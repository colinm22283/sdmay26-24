// This is the unpowered netlist.
module vga_m (clk_i,
    enable_i,
    fb_i,
    hsync_o,
    nrst_i,
    vsync_o,
    base_h_active_i,
    base_h_bporch_i,
    base_h_fporch_i,
    base_h_sync_i,
    base_v_active_i,
    base_v_bporch_i,
    base_v_fporch_i,
    base_v_sync_i,
    mport_i,
    mport_o,
    pixel_o,
    prescaler_i,
    resolution_i);
 input clk_i;
 input enable_i;
 input fb_i;
 output hsync_o;
 input nrst_i;
 output vsync_o;
 input [9:0] base_h_active_i;
 input [6:0] base_h_bporch_i;
 input [4:0] base_h_fporch_i;
 input [6:0] base_h_sync_i;
 input [8:0] base_v_active_i;
 input [3:0] base_v_bporch_i;
 input [2:0] base_v_fporch_i;
 input [2:0] base_v_sync_i;
 input [33:0] mport_i;
 output [68:0] mport_o;
 output [7:0] pixel_o;
 input [3:0] prescaler_i;
 input [3:0] resolution_i;

 wire net371;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net372;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net373;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net374;
 wire net375;
 wire net376;
 wire net405;
 wire net406;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire \base_h_active[0] ;
 wire \base_h_active[1] ;
 wire \base_h_active[2] ;
 wire \base_h_active[3] ;
 wire \base_h_active[4] ;
 wire \base_h_active[5] ;
 wire \base_h_active[6] ;
 wire \base_h_active[7] ;
 wire \base_h_active[8] ;
 wire \base_h_active[9] ;
 wire \base_h_bporch[0] ;
 wire \base_h_bporch[1] ;
 wire \base_h_bporch[2] ;
 wire \base_h_bporch[3] ;
 wire \base_h_bporch[4] ;
 wire \base_h_bporch[5] ;
 wire \base_h_bporch[6] ;
 wire \base_h_counter[0] ;
 wire \base_h_counter[1] ;
 wire \base_h_counter[2] ;
 wire \base_h_counter[3] ;
 wire \base_h_counter[4] ;
 wire \base_h_counter[5] ;
 wire \base_h_counter[6] ;
 wire \base_h_counter[7] ;
 wire \base_h_counter[8] ;
 wire \base_h_counter[9] ;
 wire \base_h_fporch[0] ;
 wire \base_h_fporch[1] ;
 wire \base_h_fporch[2] ;
 wire \base_h_fporch[3] ;
 wire \base_h_fporch[4] ;
 wire \base_h_sync[0] ;
 wire \base_h_sync[1] ;
 wire \base_h_sync[2] ;
 wire \base_h_sync[3] ;
 wire \base_h_sync[4] ;
 wire \base_h_sync[5] ;
 wire \base_h_sync[6] ;
 wire \base_v_active[0] ;
 wire \base_v_active[1] ;
 wire \base_v_active[2] ;
 wire \base_v_active[3] ;
 wire \base_v_active[4] ;
 wire \base_v_active[5] ;
 wire \base_v_active[6] ;
 wire \base_v_active[7] ;
 wire \base_v_active[8] ;
 wire \base_v_bporch[0] ;
 wire \base_v_bporch[1] ;
 wire \base_v_bporch[2] ;
 wire \base_v_bporch[3] ;
 wire \base_v_counter[0] ;
 wire \base_v_counter[1] ;
 wire \base_v_counter[2] ;
 wire \base_v_counter[3] ;
 wire \base_v_counter[4] ;
 wire \base_v_counter[5] ;
 wire \base_v_counter[6] ;
 wire \base_v_counter[7] ;
 wire \base_v_counter[8] ;
 wire \base_v_counter[9] ;
 wire \base_v_fporch[0] ;
 wire \base_v_fporch[1] ;
 wire \base_v_fporch[2] ;
 wire \base_v_sync[0] ;
 wire \base_v_sync[1] ;
 wire \base_v_sync[2] ;
 wire clknet_0_clk_i;
 wire clknet_2_0_0_clk_i;
 wire clknet_2_1_0_clk_i;
 wire clknet_2_2_0_clk_i;
 wire clknet_2_3_0_clk_i;
 wire clknet_5_0__leaf_clk_i;
 wire clknet_5_10__leaf_clk_i;
 wire clknet_5_11__leaf_clk_i;
 wire clknet_5_12__leaf_clk_i;
 wire clknet_5_13__leaf_clk_i;
 wire clknet_5_14__leaf_clk_i;
 wire clknet_5_15__leaf_clk_i;
 wire clknet_5_16__leaf_clk_i;
 wire clknet_5_17__leaf_clk_i;
 wire clknet_5_18__leaf_clk_i;
 wire clknet_5_19__leaf_clk_i;
 wire clknet_5_1__leaf_clk_i;
 wire clknet_5_20__leaf_clk_i;
 wire clknet_5_21__leaf_clk_i;
 wire clknet_5_22__leaf_clk_i;
 wire clknet_5_23__leaf_clk_i;
 wire clknet_5_24__leaf_clk_i;
 wire clknet_5_25__leaf_clk_i;
 wire clknet_5_26__leaf_clk_i;
 wire clknet_5_27__leaf_clk_i;
 wire clknet_5_28__leaf_clk_i;
 wire clknet_5_29__leaf_clk_i;
 wire clknet_5_2__leaf_clk_i;
 wire clknet_5_30__leaf_clk_i;
 wire clknet_5_31__leaf_clk_i;
 wire clknet_5_3__leaf_clk_i;
 wire clknet_5_4__leaf_clk_i;
 wire clknet_5_5__leaf_clk_i;
 wire clknet_5_6__leaf_clk_i;
 wire clknet_5_7__leaf_clk_i;
 wire clknet_5_8__leaf_clk_i;
 wire clknet_5_9__leaf_clk_i;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_100_clk_i;
 wire clknet_leaf_101_clk_i;
 wire clknet_leaf_102_clk_i;
 wire clknet_leaf_103_clk_i;
 wire clknet_leaf_104_clk_i;
 wire clknet_leaf_105_clk_i;
 wire clknet_leaf_106_clk_i;
 wire clknet_leaf_107_clk_i;
 wire clknet_leaf_108_clk_i;
 wire clknet_leaf_109_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_110_clk_i;
 wire clknet_leaf_111_clk_i;
 wire clknet_leaf_112_clk_i;
 wire clknet_leaf_113_clk_i;
 wire clknet_leaf_114_clk_i;
 wire clknet_leaf_115_clk_i;
 wire clknet_leaf_116_clk_i;
 wire clknet_leaf_117_clk_i;
 wire clknet_leaf_118_clk_i;
 wire clknet_leaf_119_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_120_clk_i;
 wire clknet_leaf_121_clk_i;
 wire clknet_leaf_122_clk_i;
 wire clknet_leaf_123_clk_i;
 wire clknet_leaf_124_clk_i;
 wire clknet_leaf_125_clk_i;
 wire clknet_leaf_126_clk_i;
 wire clknet_leaf_127_clk_i;
 wire clknet_leaf_128_clk_i;
 wire clknet_leaf_129_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_130_clk_i;
 wire clknet_leaf_131_clk_i;
 wire clknet_leaf_132_clk_i;
 wire clknet_leaf_133_clk_i;
 wire clknet_leaf_134_clk_i;
 wire clknet_leaf_135_clk_i;
 wire clknet_leaf_136_clk_i;
 wire clknet_leaf_137_clk_i;
 wire clknet_leaf_138_clk_i;
 wire clknet_leaf_139_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_140_clk_i;
 wire clknet_leaf_141_clk_i;
 wire clknet_leaf_142_clk_i;
 wire clknet_leaf_143_clk_i;
 wire clknet_leaf_144_clk_i;
 wire clknet_leaf_145_clk_i;
 wire clknet_leaf_146_clk_i;
 wire clknet_leaf_147_clk_i;
 wire clknet_leaf_148_clk_i;
 wire clknet_leaf_149_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_150_clk_i;
 wire clknet_leaf_151_clk_i;
 wire clknet_leaf_152_clk_i;
 wire clknet_leaf_153_clk_i;
 wire clknet_leaf_154_clk_i;
 wire clknet_leaf_155_clk_i;
 wire clknet_leaf_156_clk_i;
 wire clknet_leaf_157_clk_i;
 wire clknet_leaf_158_clk_i;
 wire clknet_leaf_159_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_160_clk_i;
 wire clknet_leaf_161_clk_i;
 wire clknet_leaf_162_clk_i;
 wire clknet_leaf_163_clk_i;
 wire clknet_leaf_164_clk_i;
 wire clknet_leaf_165_clk_i;
 wire clknet_leaf_166_clk_i;
 wire clknet_leaf_167_clk_i;
 wire clknet_leaf_168_clk_i;
 wire clknet_leaf_169_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_170_clk_i;
 wire clknet_leaf_171_clk_i;
 wire clknet_leaf_172_clk_i;
 wire clknet_leaf_173_clk_i;
 wire clknet_leaf_174_clk_i;
 wire clknet_leaf_175_clk_i;
 wire clknet_leaf_176_clk_i;
 wire clknet_leaf_177_clk_i;
 wire clknet_leaf_178_clk_i;
 wire clknet_leaf_179_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_180_clk_i;
 wire clknet_leaf_181_clk_i;
 wire clknet_leaf_182_clk_i;
 wire clknet_leaf_183_clk_i;
 wire clknet_leaf_184_clk_i;
 wire clknet_leaf_185_clk_i;
 wire clknet_leaf_186_clk_i;
 wire clknet_leaf_187_clk_i;
 wire clknet_leaf_188_clk_i;
 wire clknet_leaf_189_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_190_clk_i;
 wire clknet_leaf_191_clk_i;
 wire clknet_leaf_192_clk_i;
 wire clknet_leaf_193_clk_i;
 wire clknet_leaf_194_clk_i;
 wire clknet_leaf_195_clk_i;
 wire clknet_leaf_196_clk_i;
 wire clknet_leaf_197_clk_i;
 wire clknet_leaf_198_clk_i;
 wire clknet_leaf_199_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_200_clk_i;
 wire clknet_leaf_201_clk_i;
 wire clknet_leaf_202_clk_i;
 wire clknet_leaf_203_clk_i;
 wire clknet_leaf_204_clk_i;
 wire clknet_leaf_205_clk_i;
 wire clknet_leaf_206_clk_i;
 wire clknet_leaf_207_clk_i;
 wire clknet_leaf_208_clk_i;
 wire clknet_leaf_209_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_210_clk_i;
 wire clknet_leaf_211_clk_i;
 wire clknet_leaf_212_clk_i;
 wire clknet_leaf_213_clk_i;
 wire clknet_leaf_214_clk_i;
 wire clknet_leaf_215_clk_i;
 wire clknet_leaf_216_clk_i;
 wire clknet_leaf_217_clk_i;
 wire clknet_leaf_218_clk_i;
 wire clknet_leaf_219_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_220_clk_i;
 wire clknet_leaf_221_clk_i;
 wire clknet_leaf_222_clk_i;
 wire clknet_leaf_223_clk_i;
 wire clknet_leaf_224_clk_i;
 wire clknet_leaf_225_clk_i;
 wire clknet_leaf_226_clk_i;
 wire clknet_leaf_227_clk_i;
 wire clknet_leaf_228_clk_i;
 wire clknet_leaf_229_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_230_clk_i;
 wire clknet_leaf_231_clk_i;
 wire clknet_leaf_232_clk_i;
 wire clknet_leaf_233_clk_i;
 wire clknet_leaf_234_clk_i;
 wire clknet_leaf_235_clk_i;
 wire clknet_leaf_236_clk_i;
 wire clknet_leaf_237_clk_i;
 wire clknet_leaf_238_clk_i;
 wire clknet_leaf_239_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_240_clk_i;
 wire clknet_leaf_241_clk_i;
 wire clknet_leaf_242_clk_i;
 wire clknet_leaf_243_clk_i;
 wire clknet_leaf_244_clk_i;
 wire clknet_leaf_245_clk_i;
 wire clknet_leaf_246_clk_i;
 wire clknet_leaf_247_clk_i;
 wire clknet_leaf_248_clk_i;
 wire clknet_leaf_249_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_250_clk_i;
 wire clknet_leaf_251_clk_i;
 wire clknet_leaf_252_clk_i;
 wire clknet_leaf_253_clk_i;
 wire clknet_leaf_254_clk_i;
 wire clknet_leaf_255_clk_i;
 wire clknet_leaf_256_clk_i;
 wire clknet_leaf_257_clk_i;
 wire clknet_leaf_258_clk_i;
 wire clknet_leaf_259_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_260_clk_i;
 wire clknet_leaf_261_clk_i;
 wire clknet_leaf_262_clk_i;
 wire clknet_leaf_263_clk_i;
 wire clknet_leaf_264_clk_i;
 wire clknet_leaf_265_clk_i;
 wire clknet_leaf_266_clk_i;
 wire clknet_leaf_267_clk_i;
 wire clknet_leaf_268_clk_i;
 wire clknet_leaf_269_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_270_clk_i;
 wire clknet_leaf_271_clk_i;
 wire clknet_leaf_272_clk_i;
 wire clknet_leaf_273_clk_i;
 wire clknet_leaf_274_clk_i;
 wire clknet_leaf_275_clk_i;
 wire clknet_leaf_276_clk_i;
 wire clknet_leaf_277_clk_i;
 wire clknet_leaf_278_clk_i;
 wire clknet_leaf_279_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_280_clk_i;
 wire clknet_leaf_281_clk_i;
 wire clknet_leaf_282_clk_i;
 wire clknet_leaf_283_clk_i;
 wire clknet_leaf_284_clk_i;
 wire clknet_leaf_285_clk_i;
 wire clknet_leaf_286_clk_i;
 wire clknet_leaf_287_clk_i;
 wire clknet_leaf_288_clk_i;
 wire clknet_leaf_289_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_290_clk_i;
 wire clknet_leaf_291_clk_i;
 wire clknet_leaf_292_clk_i;
 wire clknet_leaf_293_clk_i;
 wire clknet_leaf_294_clk_i;
 wire clknet_leaf_295_clk_i;
 wire clknet_leaf_296_clk_i;
 wire clknet_leaf_297_clk_i;
 wire clknet_leaf_298_clk_i;
 wire clknet_leaf_299_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_300_clk_i;
 wire clknet_leaf_301_clk_i;
 wire clknet_leaf_302_clk_i;
 wire clknet_leaf_303_clk_i;
 wire clknet_leaf_304_clk_i;
 wire clknet_leaf_305_clk_i;
 wire clknet_leaf_306_clk_i;
 wire clknet_leaf_307_clk_i;
 wire clknet_leaf_308_clk_i;
 wire clknet_leaf_309_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_310_clk_i;
 wire clknet_leaf_311_clk_i;
 wire clknet_leaf_312_clk_i;
 wire clknet_leaf_313_clk_i;
 wire clknet_leaf_314_clk_i;
 wire clknet_leaf_315_clk_i;
 wire clknet_leaf_316_clk_i;
 wire clknet_leaf_317_clk_i;
 wire clknet_leaf_318_clk_i;
 wire clknet_leaf_319_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_320_clk_i;
 wire clknet_leaf_321_clk_i;
 wire clknet_leaf_322_clk_i;
 wire clknet_leaf_323_clk_i;
 wire clknet_leaf_324_clk_i;
 wire clknet_leaf_325_clk_i;
 wire clknet_leaf_326_clk_i;
 wire clknet_leaf_327_clk_i;
 wire clknet_leaf_328_clk_i;
 wire clknet_leaf_329_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_330_clk_i;
 wire clknet_leaf_331_clk_i;
 wire clknet_leaf_332_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_leaf_39_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_40_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_42_clk_i;
 wire clknet_leaf_43_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_45_clk_i;
 wire clknet_leaf_46_clk_i;
 wire clknet_leaf_47_clk_i;
 wire clknet_leaf_48_clk_i;
 wire clknet_leaf_49_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_50_clk_i;
 wire clknet_leaf_51_clk_i;
 wire clknet_leaf_52_clk_i;
 wire clknet_leaf_53_clk_i;
 wire clknet_leaf_54_clk_i;
 wire clknet_leaf_55_clk_i;
 wire clknet_leaf_56_clk_i;
 wire clknet_leaf_57_clk_i;
 wire clknet_leaf_58_clk_i;
 wire clknet_leaf_59_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_60_clk_i;
 wire clknet_leaf_61_clk_i;
 wire clknet_leaf_62_clk_i;
 wire clknet_leaf_63_clk_i;
 wire clknet_leaf_64_clk_i;
 wire clknet_leaf_65_clk_i;
 wire clknet_leaf_66_clk_i;
 wire clknet_leaf_67_clk_i;
 wire clknet_leaf_68_clk_i;
 wire clknet_leaf_69_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_70_clk_i;
 wire clknet_leaf_71_clk_i;
 wire clknet_leaf_72_clk_i;
 wire clknet_leaf_73_clk_i;
 wire clknet_leaf_74_clk_i;
 wire clknet_leaf_75_clk_i;
 wire clknet_leaf_76_clk_i;
 wire clknet_leaf_77_clk_i;
 wire clknet_leaf_78_clk_i;
 wire clknet_leaf_79_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_80_clk_i;
 wire clknet_leaf_81_clk_i;
 wire clknet_leaf_83_clk_i;
 wire clknet_leaf_84_clk_i;
 wire clknet_leaf_85_clk_i;
 wire clknet_leaf_86_clk_i;
 wire clknet_leaf_87_clk_i;
 wire clknet_leaf_88_clk_i;
 wire clknet_leaf_89_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_90_clk_i;
 wire clknet_leaf_91_clk_i;
 wire clknet_leaf_92_clk_i;
 wire clknet_leaf_93_clk_i;
 wire clknet_leaf_94_clk_i;
 wire clknet_leaf_95_clk_i;
 wire clknet_leaf_96_clk_i;
 wire clknet_leaf_97_clk_i;
 wire clknet_leaf_98_clk_i;
 wire clknet_leaf_99_clk_i;
 wire clknet_leaf_9_clk_i;
 wire \fb_read_state[0] ;
 wire \fb_read_state[1] ;
 wire \fb_read_state[2] ;
 wire \line_cache[0][0] ;
 wire \line_cache[0][1] ;
 wire \line_cache[0][2] ;
 wire \line_cache[0][3] ;
 wire \line_cache[0][4] ;
 wire \line_cache[0][5] ;
 wire \line_cache[0][6] ;
 wire \line_cache[0][7] ;
 wire \line_cache[100][0] ;
 wire \line_cache[100][1] ;
 wire \line_cache[100][2] ;
 wire \line_cache[100][3] ;
 wire \line_cache[100][4] ;
 wire \line_cache[100][5] ;
 wire \line_cache[100][6] ;
 wire \line_cache[100][7] ;
 wire \line_cache[101][0] ;
 wire \line_cache[101][1] ;
 wire \line_cache[101][2] ;
 wire \line_cache[101][3] ;
 wire \line_cache[101][4] ;
 wire \line_cache[101][5] ;
 wire \line_cache[101][6] ;
 wire \line_cache[101][7] ;
 wire \line_cache[102][0] ;
 wire \line_cache[102][1] ;
 wire \line_cache[102][2] ;
 wire \line_cache[102][3] ;
 wire \line_cache[102][4] ;
 wire \line_cache[102][5] ;
 wire \line_cache[102][6] ;
 wire \line_cache[102][7] ;
 wire \line_cache[103][0] ;
 wire \line_cache[103][1] ;
 wire \line_cache[103][2] ;
 wire \line_cache[103][3] ;
 wire \line_cache[103][4] ;
 wire \line_cache[103][5] ;
 wire \line_cache[103][6] ;
 wire \line_cache[103][7] ;
 wire \line_cache[104][0] ;
 wire \line_cache[104][1] ;
 wire \line_cache[104][2] ;
 wire \line_cache[104][3] ;
 wire \line_cache[104][4] ;
 wire \line_cache[104][5] ;
 wire \line_cache[104][6] ;
 wire \line_cache[104][7] ;
 wire \line_cache[105][0] ;
 wire \line_cache[105][1] ;
 wire \line_cache[105][2] ;
 wire \line_cache[105][3] ;
 wire \line_cache[105][4] ;
 wire \line_cache[105][5] ;
 wire \line_cache[105][6] ;
 wire \line_cache[105][7] ;
 wire \line_cache[106][0] ;
 wire \line_cache[106][1] ;
 wire \line_cache[106][2] ;
 wire \line_cache[106][3] ;
 wire \line_cache[106][4] ;
 wire \line_cache[106][5] ;
 wire \line_cache[106][6] ;
 wire \line_cache[106][7] ;
 wire \line_cache[107][0] ;
 wire \line_cache[107][1] ;
 wire \line_cache[107][2] ;
 wire \line_cache[107][3] ;
 wire \line_cache[107][4] ;
 wire \line_cache[107][5] ;
 wire \line_cache[107][6] ;
 wire \line_cache[107][7] ;
 wire \line_cache[108][0] ;
 wire \line_cache[108][1] ;
 wire \line_cache[108][2] ;
 wire \line_cache[108][3] ;
 wire \line_cache[108][4] ;
 wire \line_cache[108][5] ;
 wire \line_cache[108][6] ;
 wire \line_cache[108][7] ;
 wire \line_cache[109][0] ;
 wire \line_cache[109][1] ;
 wire \line_cache[109][2] ;
 wire \line_cache[109][3] ;
 wire \line_cache[109][4] ;
 wire \line_cache[109][5] ;
 wire \line_cache[109][6] ;
 wire \line_cache[109][7] ;
 wire \line_cache[10][0] ;
 wire \line_cache[10][1] ;
 wire \line_cache[10][2] ;
 wire \line_cache[10][3] ;
 wire \line_cache[10][4] ;
 wire \line_cache[10][5] ;
 wire \line_cache[10][6] ;
 wire \line_cache[10][7] ;
 wire \line_cache[110][0] ;
 wire \line_cache[110][1] ;
 wire \line_cache[110][2] ;
 wire \line_cache[110][3] ;
 wire \line_cache[110][4] ;
 wire \line_cache[110][5] ;
 wire \line_cache[110][6] ;
 wire \line_cache[110][7] ;
 wire \line_cache[111][0] ;
 wire \line_cache[111][1] ;
 wire \line_cache[111][2] ;
 wire \line_cache[111][3] ;
 wire \line_cache[111][4] ;
 wire \line_cache[111][5] ;
 wire \line_cache[111][6] ;
 wire \line_cache[111][7] ;
 wire \line_cache[112][0] ;
 wire \line_cache[112][1] ;
 wire \line_cache[112][2] ;
 wire \line_cache[112][3] ;
 wire \line_cache[112][4] ;
 wire \line_cache[112][5] ;
 wire \line_cache[112][6] ;
 wire \line_cache[112][7] ;
 wire \line_cache[113][0] ;
 wire \line_cache[113][1] ;
 wire \line_cache[113][2] ;
 wire \line_cache[113][3] ;
 wire \line_cache[113][4] ;
 wire \line_cache[113][5] ;
 wire \line_cache[113][6] ;
 wire \line_cache[113][7] ;
 wire \line_cache[114][0] ;
 wire \line_cache[114][1] ;
 wire \line_cache[114][2] ;
 wire \line_cache[114][3] ;
 wire \line_cache[114][4] ;
 wire \line_cache[114][5] ;
 wire \line_cache[114][6] ;
 wire \line_cache[114][7] ;
 wire \line_cache[115][0] ;
 wire \line_cache[115][1] ;
 wire \line_cache[115][2] ;
 wire \line_cache[115][3] ;
 wire \line_cache[115][4] ;
 wire \line_cache[115][5] ;
 wire \line_cache[115][6] ;
 wire \line_cache[115][7] ;
 wire \line_cache[116][0] ;
 wire \line_cache[116][1] ;
 wire \line_cache[116][2] ;
 wire \line_cache[116][3] ;
 wire \line_cache[116][4] ;
 wire \line_cache[116][5] ;
 wire \line_cache[116][6] ;
 wire \line_cache[116][7] ;
 wire \line_cache[117][0] ;
 wire \line_cache[117][1] ;
 wire \line_cache[117][2] ;
 wire \line_cache[117][3] ;
 wire \line_cache[117][4] ;
 wire \line_cache[117][5] ;
 wire \line_cache[117][6] ;
 wire \line_cache[117][7] ;
 wire \line_cache[118][0] ;
 wire \line_cache[118][1] ;
 wire \line_cache[118][2] ;
 wire \line_cache[118][3] ;
 wire \line_cache[118][4] ;
 wire \line_cache[118][5] ;
 wire \line_cache[118][6] ;
 wire \line_cache[118][7] ;
 wire \line_cache[119][0] ;
 wire \line_cache[119][1] ;
 wire \line_cache[119][2] ;
 wire \line_cache[119][3] ;
 wire \line_cache[119][4] ;
 wire \line_cache[119][5] ;
 wire \line_cache[119][6] ;
 wire \line_cache[119][7] ;
 wire \line_cache[11][0] ;
 wire \line_cache[11][1] ;
 wire \line_cache[11][2] ;
 wire \line_cache[11][3] ;
 wire \line_cache[11][4] ;
 wire \line_cache[11][5] ;
 wire \line_cache[11][6] ;
 wire \line_cache[11][7] ;
 wire \line_cache[120][0] ;
 wire \line_cache[120][1] ;
 wire \line_cache[120][2] ;
 wire \line_cache[120][3] ;
 wire \line_cache[120][4] ;
 wire \line_cache[120][5] ;
 wire \line_cache[120][6] ;
 wire \line_cache[120][7] ;
 wire \line_cache[121][0] ;
 wire \line_cache[121][1] ;
 wire \line_cache[121][2] ;
 wire \line_cache[121][3] ;
 wire \line_cache[121][4] ;
 wire \line_cache[121][5] ;
 wire \line_cache[121][6] ;
 wire \line_cache[121][7] ;
 wire \line_cache[122][0] ;
 wire \line_cache[122][1] ;
 wire \line_cache[122][2] ;
 wire \line_cache[122][3] ;
 wire \line_cache[122][4] ;
 wire \line_cache[122][5] ;
 wire \line_cache[122][6] ;
 wire \line_cache[122][7] ;
 wire \line_cache[123][0] ;
 wire \line_cache[123][1] ;
 wire \line_cache[123][2] ;
 wire \line_cache[123][3] ;
 wire \line_cache[123][4] ;
 wire \line_cache[123][5] ;
 wire \line_cache[123][6] ;
 wire \line_cache[123][7] ;
 wire \line_cache[124][0] ;
 wire \line_cache[124][1] ;
 wire \line_cache[124][2] ;
 wire \line_cache[124][3] ;
 wire \line_cache[124][4] ;
 wire \line_cache[124][5] ;
 wire \line_cache[124][6] ;
 wire \line_cache[124][7] ;
 wire \line_cache[125][0] ;
 wire \line_cache[125][1] ;
 wire \line_cache[125][2] ;
 wire \line_cache[125][3] ;
 wire \line_cache[125][4] ;
 wire \line_cache[125][5] ;
 wire \line_cache[125][6] ;
 wire \line_cache[125][7] ;
 wire \line_cache[126][0] ;
 wire \line_cache[126][1] ;
 wire \line_cache[126][2] ;
 wire \line_cache[126][3] ;
 wire \line_cache[126][4] ;
 wire \line_cache[126][5] ;
 wire \line_cache[126][6] ;
 wire \line_cache[126][7] ;
 wire \line_cache[127][0] ;
 wire \line_cache[127][1] ;
 wire \line_cache[127][2] ;
 wire \line_cache[127][3] ;
 wire \line_cache[127][4] ;
 wire \line_cache[127][5] ;
 wire \line_cache[127][6] ;
 wire \line_cache[127][7] ;
 wire \line_cache[128][0] ;
 wire \line_cache[128][1] ;
 wire \line_cache[128][2] ;
 wire \line_cache[128][3] ;
 wire \line_cache[128][4] ;
 wire \line_cache[128][5] ;
 wire \line_cache[128][6] ;
 wire \line_cache[128][7] ;
 wire \line_cache[129][0] ;
 wire \line_cache[129][1] ;
 wire \line_cache[129][2] ;
 wire \line_cache[129][3] ;
 wire \line_cache[129][4] ;
 wire \line_cache[129][5] ;
 wire \line_cache[129][6] ;
 wire \line_cache[129][7] ;
 wire \line_cache[12][0] ;
 wire \line_cache[12][1] ;
 wire \line_cache[12][2] ;
 wire \line_cache[12][3] ;
 wire \line_cache[12][4] ;
 wire \line_cache[12][5] ;
 wire \line_cache[12][6] ;
 wire \line_cache[12][7] ;
 wire \line_cache[130][0] ;
 wire \line_cache[130][1] ;
 wire \line_cache[130][2] ;
 wire \line_cache[130][3] ;
 wire \line_cache[130][4] ;
 wire \line_cache[130][5] ;
 wire \line_cache[130][6] ;
 wire \line_cache[130][7] ;
 wire \line_cache[131][0] ;
 wire \line_cache[131][1] ;
 wire \line_cache[131][2] ;
 wire \line_cache[131][3] ;
 wire \line_cache[131][4] ;
 wire \line_cache[131][5] ;
 wire \line_cache[131][6] ;
 wire \line_cache[131][7] ;
 wire \line_cache[132][0] ;
 wire \line_cache[132][1] ;
 wire \line_cache[132][2] ;
 wire \line_cache[132][3] ;
 wire \line_cache[132][4] ;
 wire \line_cache[132][5] ;
 wire \line_cache[132][6] ;
 wire \line_cache[132][7] ;
 wire \line_cache[133][0] ;
 wire \line_cache[133][1] ;
 wire \line_cache[133][2] ;
 wire \line_cache[133][3] ;
 wire \line_cache[133][4] ;
 wire \line_cache[133][5] ;
 wire \line_cache[133][6] ;
 wire \line_cache[133][7] ;
 wire \line_cache[134][0] ;
 wire \line_cache[134][1] ;
 wire \line_cache[134][2] ;
 wire \line_cache[134][3] ;
 wire \line_cache[134][4] ;
 wire \line_cache[134][5] ;
 wire \line_cache[134][6] ;
 wire \line_cache[134][7] ;
 wire \line_cache[135][0] ;
 wire \line_cache[135][1] ;
 wire \line_cache[135][2] ;
 wire \line_cache[135][3] ;
 wire \line_cache[135][4] ;
 wire \line_cache[135][5] ;
 wire \line_cache[135][6] ;
 wire \line_cache[135][7] ;
 wire \line_cache[136][0] ;
 wire \line_cache[136][1] ;
 wire \line_cache[136][2] ;
 wire \line_cache[136][3] ;
 wire \line_cache[136][4] ;
 wire \line_cache[136][5] ;
 wire \line_cache[136][6] ;
 wire \line_cache[136][7] ;
 wire \line_cache[137][0] ;
 wire \line_cache[137][1] ;
 wire \line_cache[137][2] ;
 wire \line_cache[137][3] ;
 wire \line_cache[137][4] ;
 wire \line_cache[137][5] ;
 wire \line_cache[137][6] ;
 wire \line_cache[137][7] ;
 wire \line_cache[138][0] ;
 wire \line_cache[138][1] ;
 wire \line_cache[138][2] ;
 wire \line_cache[138][3] ;
 wire \line_cache[138][4] ;
 wire \line_cache[138][5] ;
 wire \line_cache[138][6] ;
 wire \line_cache[138][7] ;
 wire \line_cache[139][0] ;
 wire \line_cache[139][1] ;
 wire \line_cache[139][2] ;
 wire \line_cache[139][3] ;
 wire \line_cache[139][4] ;
 wire \line_cache[139][5] ;
 wire \line_cache[139][6] ;
 wire \line_cache[139][7] ;
 wire \line_cache[13][0] ;
 wire \line_cache[13][1] ;
 wire \line_cache[13][2] ;
 wire \line_cache[13][3] ;
 wire \line_cache[13][4] ;
 wire \line_cache[13][5] ;
 wire \line_cache[13][6] ;
 wire \line_cache[13][7] ;
 wire \line_cache[140][0] ;
 wire \line_cache[140][1] ;
 wire \line_cache[140][2] ;
 wire \line_cache[140][3] ;
 wire \line_cache[140][4] ;
 wire \line_cache[140][5] ;
 wire \line_cache[140][6] ;
 wire \line_cache[140][7] ;
 wire \line_cache[141][0] ;
 wire \line_cache[141][1] ;
 wire \line_cache[141][2] ;
 wire \line_cache[141][3] ;
 wire \line_cache[141][4] ;
 wire \line_cache[141][5] ;
 wire \line_cache[141][6] ;
 wire \line_cache[141][7] ;
 wire \line_cache[142][0] ;
 wire \line_cache[142][1] ;
 wire \line_cache[142][2] ;
 wire \line_cache[142][3] ;
 wire \line_cache[142][4] ;
 wire \line_cache[142][5] ;
 wire \line_cache[142][6] ;
 wire \line_cache[142][7] ;
 wire \line_cache[143][0] ;
 wire \line_cache[143][1] ;
 wire \line_cache[143][2] ;
 wire \line_cache[143][3] ;
 wire \line_cache[143][4] ;
 wire \line_cache[143][5] ;
 wire \line_cache[143][6] ;
 wire \line_cache[143][7] ;
 wire \line_cache[144][0] ;
 wire \line_cache[144][1] ;
 wire \line_cache[144][2] ;
 wire \line_cache[144][3] ;
 wire \line_cache[144][4] ;
 wire \line_cache[144][5] ;
 wire \line_cache[144][6] ;
 wire \line_cache[144][7] ;
 wire \line_cache[145][0] ;
 wire \line_cache[145][1] ;
 wire \line_cache[145][2] ;
 wire \line_cache[145][3] ;
 wire \line_cache[145][4] ;
 wire \line_cache[145][5] ;
 wire \line_cache[145][6] ;
 wire \line_cache[145][7] ;
 wire \line_cache[146][0] ;
 wire \line_cache[146][1] ;
 wire \line_cache[146][2] ;
 wire \line_cache[146][3] ;
 wire \line_cache[146][4] ;
 wire \line_cache[146][5] ;
 wire \line_cache[146][6] ;
 wire \line_cache[146][7] ;
 wire \line_cache[147][0] ;
 wire \line_cache[147][1] ;
 wire \line_cache[147][2] ;
 wire \line_cache[147][3] ;
 wire \line_cache[147][4] ;
 wire \line_cache[147][5] ;
 wire \line_cache[147][6] ;
 wire \line_cache[147][7] ;
 wire \line_cache[148][0] ;
 wire \line_cache[148][1] ;
 wire \line_cache[148][2] ;
 wire \line_cache[148][3] ;
 wire \line_cache[148][4] ;
 wire \line_cache[148][5] ;
 wire \line_cache[148][6] ;
 wire \line_cache[148][7] ;
 wire \line_cache[149][0] ;
 wire \line_cache[149][1] ;
 wire \line_cache[149][2] ;
 wire \line_cache[149][3] ;
 wire \line_cache[149][4] ;
 wire \line_cache[149][5] ;
 wire \line_cache[149][6] ;
 wire \line_cache[149][7] ;
 wire \line_cache[14][0] ;
 wire \line_cache[14][1] ;
 wire \line_cache[14][2] ;
 wire \line_cache[14][3] ;
 wire \line_cache[14][4] ;
 wire \line_cache[14][5] ;
 wire \line_cache[14][6] ;
 wire \line_cache[14][7] ;
 wire \line_cache[150][0] ;
 wire \line_cache[150][1] ;
 wire \line_cache[150][2] ;
 wire \line_cache[150][3] ;
 wire \line_cache[150][4] ;
 wire \line_cache[150][5] ;
 wire \line_cache[150][6] ;
 wire \line_cache[150][7] ;
 wire \line_cache[151][0] ;
 wire \line_cache[151][1] ;
 wire \line_cache[151][2] ;
 wire \line_cache[151][3] ;
 wire \line_cache[151][4] ;
 wire \line_cache[151][5] ;
 wire \line_cache[151][6] ;
 wire \line_cache[151][7] ;
 wire \line_cache[152][0] ;
 wire \line_cache[152][1] ;
 wire \line_cache[152][2] ;
 wire \line_cache[152][3] ;
 wire \line_cache[152][4] ;
 wire \line_cache[152][5] ;
 wire \line_cache[152][6] ;
 wire \line_cache[152][7] ;
 wire \line_cache[153][0] ;
 wire \line_cache[153][1] ;
 wire \line_cache[153][2] ;
 wire \line_cache[153][3] ;
 wire \line_cache[153][4] ;
 wire \line_cache[153][5] ;
 wire \line_cache[153][6] ;
 wire \line_cache[153][7] ;
 wire \line_cache[154][0] ;
 wire \line_cache[154][1] ;
 wire \line_cache[154][2] ;
 wire \line_cache[154][3] ;
 wire \line_cache[154][4] ;
 wire \line_cache[154][5] ;
 wire \line_cache[154][6] ;
 wire \line_cache[154][7] ;
 wire \line_cache[155][0] ;
 wire \line_cache[155][1] ;
 wire \line_cache[155][2] ;
 wire \line_cache[155][3] ;
 wire \line_cache[155][4] ;
 wire \line_cache[155][5] ;
 wire \line_cache[155][6] ;
 wire \line_cache[155][7] ;
 wire \line_cache[156][0] ;
 wire \line_cache[156][1] ;
 wire \line_cache[156][2] ;
 wire \line_cache[156][3] ;
 wire \line_cache[156][4] ;
 wire \line_cache[156][5] ;
 wire \line_cache[156][6] ;
 wire \line_cache[156][7] ;
 wire \line_cache[157][0] ;
 wire \line_cache[157][1] ;
 wire \line_cache[157][2] ;
 wire \line_cache[157][3] ;
 wire \line_cache[157][4] ;
 wire \line_cache[157][5] ;
 wire \line_cache[157][6] ;
 wire \line_cache[157][7] ;
 wire \line_cache[158][0] ;
 wire \line_cache[158][1] ;
 wire \line_cache[158][2] ;
 wire \line_cache[158][3] ;
 wire \line_cache[158][4] ;
 wire \line_cache[158][5] ;
 wire \line_cache[158][6] ;
 wire \line_cache[158][7] ;
 wire \line_cache[159][0] ;
 wire \line_cache[159][1] ;
 wire \line_cache[159][2] ;
 wire \line_cache[159][3] ;
 wire \line_cache[159][4] ;
 wire \line_cache[159][5] ;
 wire \line_cache[159][6] ;
 wire \line_cache[159][7] ;
 wire \line_cache[15][0] ;
 wire \line_cache[15][1] ;
 wire \line_cache[15][2] ;
 wire \line_cache[15][3] ;
 wire \line_cache[15][4] ;
 wire \line_cache[15][5] ;
 wire \line_cache[15][6] ;
 wire \line_cache[15][7] ;
 wire \line_cache[160][0] ;
 wire \line_cache[160][1] ;
 wire \line_cache[160][2] ;
 wire \line_cache[160][3] ;
 wire \line_cache[160][4] ;
 wire \line_cache[160][5] ;
 wire \line_cache[160][6] ;
 wire \line_cache[160][7] ;
 wire \line_cache[161][0] ;
 wire \line_cache[161][1] ;
 wire \line_cache[161][2] ;
 wire \line_cache[161][3] ;
 wire \line_cache[161][4] ;
 wire \line_cache[161][5] ;
 wire \line_cache[161][6] ;
 wire \line_cache[161][7] ;
 wire \line_cache[162][0] ;
 wire \line_cache[162][1] ;
 wire \line_cache[162][2] ;
 wire \line_cache[162][3] ;
 wire \line_cache[162][4] ;
 wire \line_cache[162][5] ;
 wire \line_cache[162][6] ;
 wire \line_cache[162][7] ;
 wire \line_cache[163][0] ;
 wire \line_cache[163][1] ;
 wire \line_cache[163][2] ;
 wire \line_cache[163][3] ;
 wire \line_cache[163][4] ;
 wire \line_cache[163][5] ;
 wire \line_cache[163][6] ;
 wire \line_cache[163][7] ;
 wire \line_cache[164][0] ;
 wire \line_cache[164][1] ;
 wire \line_cache[164][2] ;
 wire \line_cache[164][3] ;
 wire \line_cache[164][4] ;
 wire \line_cache[164][5] ;
 wire \line_cache[164][6] ;
 wire \line_cache[164][7] ;
 wire \line_cache[165][0] ;
 wire \line_cache[165][1] ;
 wire \line_cache[165][2] ;
 wire \line_cache[165][3] ;
 wire \line_cache[165][4] ;
 wire \line_cache[165][5] ;
 wire \line_cache[165][6] ;
 wire \line_cache[165][7] ;
 wire \line_cache[166][0] ;
 wire \line_cache[166][1] ;
 wire \line_cache[166][2] ;
 wire \line_cache[166][3] ;
 wire \line_cache[166][4] ;
 wire \line_cache[166][5] ;
 wire \line_cache[166][6] ;
 wire \line_cache[166][7] ;
 wire \line_cache[167][0] ;
 wire \line_cache[167][1] ;
 wire \line_cache[167][2] ;
 wire \line_cache[167][3] ;
 wire \line_cache[167][4] ;
 wire \line_cache[167][5] ;
 wire \line_cache[167][6] ;
 wire \line_cache[167][7] ;
 wire \line_cache[168][0] ;
 wire \line_cache[168][1] ;
 wire \line_cache[168][2] ;
 wire \line_cache[168][3] ;
 wire \line_cache[168][4] ;
 wire \line_cache[168][5] ;
 wire \line_cache[168][6] ;
 wire \line_cache[168][7] ;
 wire \line_cache[169][0] ;
 wire \line_cache[169][1] ;
 wire \line_cache[169][2] ;
 wire \line_cache[169][3] ;
 wire \line_cache[169][4] ;
 wire \line_cache[169][5] ;
 wire \line_cache[169][6] ;
 wire \line_cache[169][7] ;
 wire \line_cache[16][0] ;
 wire \line_cache[16][1] ;
 wire \line_cache[16][2] ;
 wire \line_cache[16][3] ;
 wire \line_cache[16][4] ;
 wire \line_cache[16][5] ;
 wire \line_cache[16][6] ;
 wire \line_cache[16][7] ;
 wire \line_cache[170][0] ;
 wire \line_cache[170][1] ;
 wire \line_cache[170][2] ;
 wire \line_cache[170][3] ;
 wire \line_cache[170][4] ;
 wire \line_cache[170][5] ;
 wire \line_cache[170][6] ;
 wire \line_cache[170][7] ;
 wire \line_cache[171][0] ;
 wire \line_cache[171][1] ;
 wire \line_cache[171][2] ;
 wire \line_cache[171][3] ;
 wire \line_cache[171][4] ;
 wire \line_cache[171][5] ;
 wire \line_cache[171][6] ;
 wire \line_cache[171][7] ;
 wire \line_cache[172][0] ;
 wire \line_cache[172][1] ;
 wire \line_cache[172][2] ;
 wire \line_cache[172][3] ;
 wire \line_cache[172][4] ;
 wire \line_cache[172][5] ;
 wire \line_cache[172][6] ;
 wire \line_cache[172][7] ;
 wire \line_cache[173][0] ;
 wire \line_cache[173][1] ;
 wire \line_cache[173][2] ;
 wire \line_cache[173][3] ;
 wire \line_cache[173][4] ;
 wire \line_cache[173][5] ;
 wire \line_cache[173][6] ;
 wire \line_cache[173][7] ;
 wire \line_cache[174][0] ;
 wire \line_cache[174][1] ;
 wire \line_cache[174][2] ;
 wire \line_cache[174][3] ;
 wire \line_cache[174][4] ;
 wire \line_cache[174][5] ;
 wire \line_cache[174][6] ;
 wire \line_cache[174][7] ;
 wire \line_cache[175][0] ;
 wire \line_cache[175][1] ;
 wire \line_cache[175][2] ;
 wire \line_cache[175][3] ;
 wire \line_cache[175][4] ;
 wire \line_cache[175][5] ;
 wire \line_cache[175][6] ;
 wire \line_cache[175][7] ;
 wire \line_cache[176][0] ;
 wire \line_cache[176][1] ;
 wire \line_cache[176][2] ;
 wire \line_cache[176][3] ;
 wire \line_cache[176][4] ;
 wire \line_cache[176][5] ;
 wire \line_cache[176][6] ;
 wire \line_cache[176][7] ;
 wire \line_cache[177][0] ;
 wire \line_cache[177][1] ;
 wire \line_cache[177][2] ;
 wire \line_cache[177][3] ;
 wire \line_cache[177][4] ;
 wire \line_cache[177][5] ;
 wire \line_cache[177][6] ;
 wire \line_cache[177][7] ;
 wire \line_cache[178][0] ;
 wire \line_cache[178][1] ;
 wire \line_cache[178][2] ;
 wire \line_cache[178][3] ;
 wire \line_cache[178][4] ;
 wire \line_cache[178][5] ;
 wire \line_cache[178][6] ;
 wire \line_cache[178][7] ;
 wire \line_cache[179][0] ;
 wire \line_cache[179][1] ;
 wire \line_cache[179][2] ;
 wire \line_cache[179][3] ;
 wire \line_cache[179][4] ;
 wire \line_cache[179][5] ;
 wire \line_cache[179][6] ;
 wire \line_cache[179][7] ;
 wire \line_cache[17][0] ;
 wire \line_cache[17][1] ;
 wire \line_cache[17][2] ;
 wire \line_cache[17][3] ;
 wire \line_cache[17][4] ;
 wire \line_cache[17][5] ;
 wire \line_cache[17][6] ;
 wire \line_cache[17][7] ;
 wire \line_cache[180][0] ;
 wire \line_cache[180][1] ;
 wire \line_cache[180][2] ;
 wire \line_cache[180][3] ;
 wire \line_cache[180][4] ;
 wire \line_cache[180][5] ;
 wire \line_cache[180][6] ;
 wire \line_cache[180][7] ;
 wire \line_cache[181][0] ;
 wire \line_cache[181][1] ;
 wire \line_cache[181][2] ;
 wire \line_cache[181][3] ;
 wire \line_cache[181][4] ;
 wire \line_cache[181][5] ;
 wire \line_cache[181][6] ;
 wire \line_cache[181][7] ;
 wire \line_cache[182][0] ;
 wire \line_cache[182][1] ;
 wire \line_cache[182][2] ;
 wire \line_cache[182][3] ;
 wire \line_cache[182][4] ;
 wire \line_cache[182][5] ;
 wire \line_cache[182][6] ;
 wire \line_cache[182][7] ;
 wire \line_cache[183][0] ;
 wire \line_cache[183][1] ;
 wire \line_cache[183][2] ;
 wire \line_cache[183][3] ;
 wire \line_cache[183][4] ;
 wire \line_cache[183][5] ;
 wire \line_cache[183][6] ;
 wire \line_cache[183][7] ;
 wire \line_cache[184][0] ;
 wire \line_cache[184][1] ;
 wire \line_cache[184][2] ;
 wire \line_cache[184][3] ;
 wire \line_cache[184][4] ;
 wire \line_cache[184][5] ;
 wire \line_cache[184][6] ;
 wire \line_cache[184][7] ;
 wire \line_cache[185][0] ;
 wire \line_cache[185][1] ;
 wire \line_cache[185][2] ;
 wire \line_cache[185][3] ;
 wire \line_cache[185][4] ;
 wire \line_cache[185][5] ;
 wire \line_cache[185][6] ;
 wire \line_cache[185][7] ;
 wire \line_cache[186][0] ;
 wire \line_cache[186][1] ;
 wire \line_cache[186][2] ;
 wire \line_cache[186][3] ;
 wire \line_cache[186][4] ;
 wire \line_cache[186][5] ;
 wire \line_cache[186][6] ;
 wire \line_cache[186][7] ;
 wire \line_cache[187][0] ;
 wire \line_cache[187][1] ;
 wire \line_cache[187][2] ;
 wire \line_cache[187][3] ;
 wire \line_cache[187][4] ;
 wire \line_cache[187][5] ;
 wire \line_cache[187][6] ;
 wire \line_cache[187][7] ;
 wire \line_cache[188][0] ;
 wire \line_cache[188][1] ;
 wire \line_cache[188][2] ;
 wire \line_cache[188][3] ;
 wire \line_cache[188][4] ;
 wire \line_cache[188][5] ;
 wire \line_cache[188][6] ;
 wire \line_cache[188][7] ;
 wire \line_cache[189][0] ;
 wire \line_cache[189][1] ;
 wire \line_cache[189][2] ;
 wire \line_cache[189][3] ;
 wire \line_cache[189][4] ;
 wire \line_cache[189][5] ;
 wire \line_cache[189][6] ;
 wire \line_cache[189][7] ;
 wire \line_cache[18][0] ;
 wire \line_cache[18][1] ;
 wire \line_cache[18][2] ;
 wire \line_cache[18][3] ;
 wire \line_cache[18][4] ;
 wire \line_cache[18][5] ;
 wire \line_cache[18][6] ;
 wire \line_cache[18][7] ;
 wire \line_cache[190][0] ;
 wire \line_cache[190][1] ;
 wire \line_cache[190][2] ;
 wire \line_cache[190][3] ;
 wire \line_cache[190][4] ;
 wire \line_cache[190][5] ;
 wire \line_cache[190][6] ;
 wire \line_cache[190][7] ;
 wire \line_cache[191][0] ;
 wire \line_cache[191][1] ;
 wire \line_cache[191][2] ;
 wire \line_cache[191][3] ;
 wire \line_cache[191][4] ;
 wire \line_cache[191][5] ;
 wire \line_cache[191][6] ;
 wire \line_cache[191][7] ;
 wire \line_cache[192][0] ;
 wire \line_cache[192][1] ;
 wire \line_cache[192][2] ;
 wire \line_cache[192][3] ;
 wire \line_cache[192][4] ;
 wire \line_cache[192][5] ;
 wire \line_cache[192][6] ;
 wire \line_cache[192][7] ;
 wire \line_cache[193][0] ;
 wire \line_cache[193][1] ;
 wire \line_cache[193][2] ;
 wire \line_cache[193][3] ;
 wire \line_cache[193][4] ;
 wire \line_cache[193][5] ;
 wire \line_cache[193][6] ;
 wire \line_cache[193][7] ;
 wire \line_cache[194][0] ;
 wire \line_cache[194][1] ;
 wire \line_cache[194][2] ;
 wire \line_cache[194][3] ;
 wire \line_cache[194][4] ;
 wire \line_cache[194][5] ;
 wire \line_cache[194][6] ;
 wire \line_cache[194][7] ;
 wire \line_cache[195][0] ;
 wire \line_cache[195][1] ;
 wire \line_cache[195][2] ;
 wire \line_cache[195][3] ;
 wire \line_cache[195][4] ;
 wire \line_cache[195][5] ;
 wire \line_cache[195][6] ;
 wire \line_cache[195][7] ;
 wire \line_cache[196][0] ;
 wire \line_cache[196][1] ;
 wire \line_cache[196][2] ;
 wire \line_cache[196][3] ;
 wire \line_cache[196][4] ;
 wire \line_cache[196][5] ;
 wire \line_cache[196][6] ;
 wire \line_cache[196][7] ;
 wire \line_cache[197][0] ;
 wire \line_cache[197][1] ;
 wire \line_cache[197][2] ;
 wire \line_cache[197][3] ;
 wire \line_cache[197][4] ;
 wire \line_cache[197][5] ;
 wire \line_cache[197][6] ;
 wire \line_cache[197][7] ;
 wire \line_cache[198][0] ;
 wire \line_cache[198][1] ;
 wire \line_cache[198][2] ;
 wire \line_cache[198][3] ;
 wire \line_cache[198][4] ;
 wire \line_cache[198][5] ;
 wire \line_cache[198][6] ;
 wire \line_cache[198][7] ;
 wire \line_cache[199][0] ;
 wire \line_cache[199][1] ;
 wire \line_cache[199][2] ;
 wire \line_cache[199][3] ;
 wire \line_cache[199][4] ;
 wire \line_cache[199][5] ;
 wire \line_cache[199][6] ;
 wire \line_cache[199][7] ;
 wire \line_cache[19][0] ;
 wire \line_cache[19][1] ;
 wire \line_cache[19][2] ;
 wire \line_cache[19][3] ;
 wire \line_cache[19][4] ;
 wire \line_cache[19][5] ;
 wire \line_cache[19][6] ;
 wire \line_cache[19][7] ;
 wire \line_cache[1][0] ;
 wire \line_cache[1][1] ;
 wire \line_cache[1][2] ;
 wire \line_cache[1][3] ;
 wire \line_cache[1][4] ;
 wire \line_cache[1][5] ;
 wire \line_cache[1][6] ;
 wire \line_cache[1][7] ;
 wire \line_cache[200][0] ;
 wire \line_cache[200][1] ;
 wire \line_cache[200][2] ;
 wire \line_cache[200][3] ;
 wire \line_cache[200][4] ;
 wire \line_cache[200][5] ;
 wire \line_cache[200][6] ;
 wire \line_cache[200][7] ;
 wire \line_cache[201][0] ;
 wire \line_cache[201][1] ;
 wire \line_cache[201][2] ;
 wire \line_cache[201][3] ;
 wire \line_cache[201][4] ;
 wire \line_cache[201][5] ;
 wire \line_cache[201][6] ;
 wire \line_cache[201][7] ;
 wire \line_cache[202][0] ;
 wire \line_cache[202][1] ;
 wire \line_cache[202][2] ;
 wire \line_cache[202][3] ;
 wire \line_cache[202][4] ;
 wire \line_cache[202][5] ;
 wire \line_cache[202][6] ;
 wire \line_cache[202][7] ;
 wire \line_cache[203][0] ;
 wire \line_cache[203][1] ;
 wire \line_cache[203][2] ;
 wire \line_cache[203][3] ;
 wire \line_cache[203][4] ;
 wire \line_cache[203][5] ;
 wire \line_cache[203][6] ;
 wire \line_cache[203][7] ;
 wire \line_cache[204][0] ;
 wire \line_cache[204][1] ;
 wire \line_cache[204][2] ;
 wire \line_cache[204][3] ;
 wire \line_cache[204][4] ;
 wire \line_cache[204][5] ;
 wire \line_cache[204][6] ;
 wire \line_cache[204][7] ;
 wire \line_cache[205][0] ;
 wire \line_cache[205][1] ;
 wire \line_cache[205][2] ;
 wire \line_cache[205][3] ;
 wire \line_cache[205][4] ;
 wire \line_cache[205][5] ;
 wire \line_cache[205][6] ;
 wire \line_cache[205][7] ;
 wire \line_cache[206][0] ;
 wire \line_cache[206][1] ;
 wire \line_cache[206][2] ;
 wire \line_cache[206][3] ;
 wire \line_cache[206][4] ;
 wire \line_cache[206][5] ;
 wire \line_cache[206][6] ;
 wire \line_cache[206][7] ;
 wire \line_cache[207][0] ;
 wire \line_cache[207][1] ;
 wire \line_cache[207][2] ;
 wire \line_cache[207][3] ;
 wire \line_cache[207][4] ;
 wire \line_cache[207][5] ;
 wire \line_cache[207][6] ;
 wire \line_cache[207][7] ;
 wire \line_cache[208][0] ;
 wire \line_cache[208][1] ;
 wire \line_cache[208][2] ;
 wire \line_cache[208][3] ;
 wire \line_cache[208][4] ;
 wire \line_cache[208][5] ;
 wire \line_cache[208][6] ;
 wire \line_cache[208][7] ;
 wire \line_cache[209][0] ;
 wire \line_cache[209][1] ;
 wire \line_cache[209][2] ;
 wire \line_cache[209][3] ;
 wire \line_cache[209][4] ;
 wire \line_cache[209][5] ;
 wire \line_cache[209][6] ;
 wire \line_cache[209][7] ;
 wire \line_cache[20][0] ;
 wire \line_cache[20][1] ;
 wire \line_cache[20][2] ;
 wire \line_cache[20][3] ;
 wire \line_cache[20][4] ;
 wire \line_cache[20][5] ;
 wire \line_cache[20][6] ;
 wire \line_cache[20][7] ;
 wire \line_cache[210][0] ;
 wire \line_cache[210][1] ;
 wire \line_cache[210][2] ;
 wire \line_cache[210][3] ;
 wire \line_cache[210][4] ;
 wire \line_cache[210][5] ;
 wire \line_cache[210][6] ;
 wire \line_cache[210][7] ;
 wire \line_cache[211][0] ;
 wire \line_cache[211][1] ;
 wire \line_cache[211][2] ;
 wire \line_cache[211][3] ;
 wire \line_cache[211][4] ;
 wire \line_cache[211][5] ;
 wire \line_cache[211][6] ;
 wire \line_cache[211][7] ;
 wire \line_cache[212][0] ;
 wire \line_cache[212][1] ;
 wire \line_cache[212][2] ;
 wire \line_cache[212][3] ;
 wire \line_cache[212][4] ;
 wire \line_cache[212][5] ;
 wire \line_cache[212][6] ;
 wire \line_cache[212][7] ;
 wire \line_cache[213][0] ;
 wire \line_cache[213][1] ;
 wire \line_cache[213][2] ;
 wire \line_cache[213][3] ;
 wire \line_cache[213][4] ;
 wire \line_cache[213][5] ;
 wire \line_cache[213][6] ;
 wire \line_cache[213][7] ;
 wire \line_cache[214][0] ;
 wire \line_cache[214][1] ;
 wire \line_cache[214][2] ;
 wire \line_cache[214][3] ;
 wire \line_cache[214][4] ;
 wire \line_cache[214][5] ;
 wire \line_cache[214][6] ;
 wire \line_cache[214][7] ;
 wire \line_cache[215][0] ;
 wire \line_cache[215][1] ;
 wire \line_cache[215][2] ;
 wire \line_cache[215][3] ;
 wire \line_cache[215][4] ;
 wire \line_cache[215][5] ;
 wire \line_cache[215][6] ;
 wire \line_cache[215][7] ;
 wire \line_cache[216][0] ;
 wire \line_cache[216][1] ;
 wire \line_cache[216][2] ;
 wire \line_cache[216][3] ;
 wire \line_cache[216][4] ;
 wire \line_cache[216][5] ;
 wire \line_cache[216][6] ;
 wire \line_cache[216][7] ;
 wire \line_cache[217][0] ;
 wire \line_cache[217][1] ;
 wire \line_cache[217][2] ;
 wire \line_cache[217][3] ;
 wire \line_cache[217][4] ;
 wire \line_cache[217][5] ;
 wire \line_cache[217][6] ;
 wire \line_cache[217][7] ;
 wire \line_cache[218][0] ;
 wire \line_cache[218][1] ;
 wire \line_cache[218][2] ;
 wire \line_cache[218][3] ;
 wire \line_cache[218][4] ;
 wire \line_cache[218][5] ;
 wire \line_cache[218][6] ;
 wire \line_cache[218][7] ;
 wire \line_cache[219][0] ;
 wire \line_cache[219][1] ;
 wire \line_cache[219][2] ;
 wire \line_cache[219][3] ;
 wire \line_cache[219][4] ;
 wire \line_cache[219][5] ;
 wire \line_cache[219][6] ;
 wire \line_cache[219][7] ;
 wire \line_cache[21][0] ;
 wire \line_cache[21][1] ;
 wire \line_cache[21][2] ;
 wire \line_cache[21][3] ;
 wire \line_cache[21][4] ;
 wire \line_cache[21][5] ;
 wire \line_cache[21][6] ;
 wire \line_cache[21][7] ;
 wire \line_cache[220][0] ;
 wire \line_cache[220][1] ;
 wire \line_cache[220][2] ;
 wire \line_cache[220][3] ;
 wire \line_cache[220][4] ;
 wire \line_cache[220][5] ;
 wire \line_cache[220][6] ;
 wire \line_cache[220][7] ;
 wire \line_cache[221][0] ;
 wire \line_cache[221][1] ;
 wire \line_cache[221][2] ;
 wire \line_cache[221][3] ;
 wire \line_cache[221][4] ;
 wire \line_cache[221][5] ;
 wire \line_cache[221][6] ;
 wire \line_cache[221][7] ;
 wire \line_cache[222][0] ;
 wire \line_cache[222][1] ;
 wire \line_cache[222][2] ;
 wire \line_cache[222][3] ;
 wire \line_cache[222][4] ;
 wire \line_cache[222][5] ;
 wire \line_cache[222][6] ;
 wire \line_cache[222][7] ;
 wire \line_cache[223][0] ;
 wire \line_cache[223][1] ;
 wire \line_cache[223][2] ;
 wire \line_cache[223][3] ;
 wire \line_cache[223][4] ;
 wire \line_cache[223][5] ;
 wire \line_cache[223][6] ;
 wire \line_cache[223][7] ;
 wire \line_cache[224][0] ;
 wire \line_cache[224][1] ;
 wire \line_cache[224][2] ;
 wire \line_cache[224][3] ;
 wire \line_cache[224][4] ;
 wire \line_cache[224][5] ;
 wire \line_cache[224][6] ;
 wire \line_cache[224][7] ;
 wire \line_cache[225][0] ;
 wire \line_cache[225][1] ;
 wire \line_cache[225][2] ;
 wire \line_cache[225][3] ;
 wire \line_cache[225][4] ;
 wire \line_cache[225][5] ;
 wire \line_cache[225][6] ;
 wire \line_cache[225][7] ;
 wire \line_cache[226][0] ;
 wire \line_cache[226][1] ;
 wire \line_cache[226][2] ;
 wire \line_cache[226][3] ;
 wire \line_cache[226][4] ;
 wire \line_cache[226][5] ;
 wire \line_cache[226][6] ;
 wire \line_cache[226][7] ;
 wire \line_cache[227][0] ;
 wire \line_cache[227][1] ;
 wire \line_cache[227][2] ;
 wire \line_cache[227][3] ;
 wire \line_cache[227][4] ;
 wire \line_cache[227][5] ;
 wire \line_cache[227][6] ;
 wire \line_cache[227][7] ;
 wire \line_cache[228][0] ;
 wire \line_cache[228][1] ;
 wire \line_cache[228][2] ;
 wire \line_cache[228][3] ;
 wire \line_cache[228][4] ;
 wire \line_cache[228][5] ;
 wire \line_cache[228][6] ;
 wire \line_cache[228][7] ;
 wire \line_cache[229][0] ;
 wire \line_cache[229][1] ;
 wire \line_cache[229][2] ;
 wire \line_cache[229][3] ;
 wire \line_cache[229][4] ;
 wire \line_cache[229][5] ;
 wire \line_cache[229][6] ;
 wire \line_cache[229][7] ;
 wire \line_cache[22][0] ;
 wire \line_cache[22][1] ;
 wire \line_cache[22][2] ;
 wire \line_cache[22][3] ;
 wire \line_cache[22][4] ;
 wire \line_cache[22][5] ;
 wire \line_cache[22][6] ;
 wire \line_cache[22][7] ;
 wire \line_cache[230][0] ;
 wire \line_cache[230][1] ;
 wire \line_cache[230][2] ;
 wire \line_cache[230][3] ;
 wire \line_cache[230][4] ;
 wire \line_cache[230][5] ;
 wire \line_cache[230][6] ;
 wire \line_cache[230][7] ;
 wire \line_cache[231][0] ;
 wire \line_cache[231][1] ;
 wire \line_cache[231][2] ;
 wire \line_cache[231][3] ;
 wire \line_cache[231][4] ;
 wire \line_cache[231][5] ;
 wire \line_cache[231][6] ;
 wire \line_cache[231][7] ;
 wire \line_cache[232][0] ;
 wire \line_cache[232][1] ;
 wire \line_cache[232][2] ;
 wire \line_cache[232][3] ;
 wire \line_cache[232][4] ;
 wire \line_cache[232][5] ;
 wire \line_cache[232][6] ;
 wire \line_cache[232][7] ;
 wire \line_cache[233][0] ;
 wire \line_cache[233][1] ;
 wire \line_cache[233][2] ;
 wire \line_cache[233][3] ;
 wire \line_cache[233][4] ;
 wire \line_cache[233][5] ;
 wire \line_cache[233][6] ;
 wire \line_cache[233][7] ;
 wire \line_cache[234][0] ;
 wire \line_cache[234][1] ;
 wire \line_cache[234][2] ;
 wire \line_cache[234][3] ;
 wire \line_cache[234][4] ;
 wire \line_cache[234][5] ;
 wire \line_cache[234][6] ;
 wire \line_cache[234][7] ;
 wire \line_cache[235][0] ;
 wire \line_cache[235][1] ;
 wire \line_cache[235][2] ;
 wire \line_cache[235][3] ;
 wire \line_cache[235][4] ;
 wire \line_cache[235][5] ;
 wire \line_cache[235][6] ;
 wire \line_cache[235][7] ;
 wire \line_cache[236][0] ;
 wire \line_cache[236][1] ;
 wire \line_cache[236][2] ;
 wire \line_cache[236][3] ;
 wire \line_cache[236][4] ;
 wire \line_cache[236][5] ;
 wire \line_cache[236][6] ;
 wire \line_cache[236][7] ;
 wire \line_cache[237][0] ;
 wire \line_cache[237][1] ;
 wire \line_cache[237][2] ;
 wire \line_cache[237][3] ;
 wire \line_cache[237][4] ;
 wire \line_cache[237][5] ;
 wire \line_cache[237][6] ;
 wire \line_cache[237][7] ;
 wire \line_cache[238][0] ;
 wire \line_cache[238][1] ;
 wire \line_cache[238][2] ;
 wire \line_cache[238][3] ;
 wire \line_cache[238][4] ;
 wire \line_cache[238][5] ;
 wire \line_cache[238][6] ;
 wire \line_cache[238][7] ;
 wire \line_cache[239][0] ;
 wire \line_cache[239][1] ;
 wire \line_cache[239][2] ;
 wire \line_cache[239][3] ;
 wire \line_cache[239][4] ;
 wire \line_cache[239][5] ;
 wire \line_cache[239][6] ;
 wire \line_cache[239][7] ;
 wire \line_cache[23][0] ;
 wire \line_cache[23][1] ;
 wire \line_cache[23][2] ;
 wire \line_cache[23][3] ;
 wire \line_cache[23][4] ;
 wire \line_cache[23][5] ;
 wire \line_cache[23][6] ;
 wire \line_cache[23][7] ;
 wire \line_cache[240][0] ;
 wire \line_cache[240][1] ;
 wire \line_cache[240][2] ;
 wire \line_cache[240][3] ;
 wire \line_cache[240][4] ;
 wire \line_cache[240][5] ;
 wire \line_cache[240][6] ;
 wire \line_cache[240][7] ;
 wire \line_cache[241][0] ;
 wire \line_cache[241][1] ;
 wire \line_cache[241][2] ;
 wire \line_cache[241][3] ;
 wire \line_cache[241][4] ;
 wire \line_cache[241][5] ;
 wire \line_cache[241][6] ;
 wire \line_cache[241][7] ;
 wire \line_cache[242][0] ;
 wire \line_cache[242][1] ;
 wire \line_cache[242][2] ;
 wire \line_cache[242][3] ;
 wire \line_cache[242][4] ;
 wire \line_cache[242][5] ;
 wire \line_cache[242][6] ;
 wire \line_cache[242][7] ;
 wire \line_cache[243][0] ;
 wire \line_cache[243][1] ;
 wire \line_cache[243][2] ;
 wire \line_cache[243][3] ;
 wire \line_cache[243][4] ;
 wire \line_cache[243][5] ;
 wire \line_cache[243][6] ;
 wire \line_cache[243][7] ;
 wire \line_cache[244][0] ;
 wire \line_cache[244][1] ;
 wire \line_cache[244][2] ;
 wire \line_cache[244][3] ;
 wire \line_cache[244][4] ;
 wire \line_cache[244][5] ;
 wire \line_cache[244][6] ;
 wire \line_cache[244][7] ;
 wire \line_cache[245][0] ;
 wire \line_cache[245][1] ;
 wire \line_cache[245][2] ;
 wire \line_cache[245][3] ;
 wire \line_cache[245][4] ;
 wire \line_cache[245][5] ;
 wire \line_cache[245][6] ;
 wire \line_cache[245][7] ;
 wire \line_cache[246][0] ;
 wire \line_cache[246][1] ;
 wire \line_cache[246][2] ;
 wire \line_cache[246][3] ;
 wire \line_cache[246][4] ;
 wire \line_cache[246][5] ;
 wire \line_cache[246][6] ;
 wire \line_cache[246][7] ;
 wire \line_cache[247][0] ;
 wire \line_cache[247][1] ;
 wire \line_cache[247][2] ;
 wire \line_cache[247][3] ;
 wire \line_cache[247][4] ;
 wire \line_cache[247][5] ;
 wire \line_cache[247][6] ;
 wire \line_cache[247][7] ;
 wire \line_cache[248][0] ;
 wire \line_cache[248][1] ;
 wire \line_cache[248][2] ;
 wire \line_cache[248][3] ;
 wire \line_cache[248][4] ;
 wire \line_cache[248][5] ;
 wire \line_cache[248][6] ;
 wire \line_cache[248][7] ;
 wire \line_cache[249][0] ;
 wire \line_cache[249][1] ;
 wire \line_cache[249][2] ;
 wire \line_cache[249][3] ;
 wire \line_cache[249][4] ;
 wire \line_cache[249][5] ;
 wire \line_cache[249][6] ;
 wire \line_cache[249][7] ;
 wire \line_cache[24][0] ;
 wire \line_cache[24][1] ;
 wire \line_cache[24][2] ;
 wire \line_cache[24][3] ;
 wire \line_cache[24][4] ;
 wire \line_cache[24][5] ;
 wire \line_cache[24][6] ;
 wire \line_cache[24][7] ;
 wire \line_cache[250][0] ;
 wire \line_cache[250][1] ;
 wire \line_cache[250][2] ;
 wire \line_cache[250][3] ;
 wire \line_cache[250][4] ;
 wire \line_cache[250][5] ;
 wire \line_cache[250][6] ;
 wire \line_cache[250][7] ;
 wire \line_cache[251][0] ;
 wire \line_cache[251][1] ;
 wire \line_cache[251][2] ;
 wire \line_cache[251][3] ;
 wire \line_cache[251][4] ;
 wire \line_cache[251][5] ;
 wire \line_cache[251][6] ;
 wire \line_cache[251][7] ;
 wire \line_cache[252][0] ;
 wire \line_cache[252][1] ;
 wire \line_cache[252][2] ;
 wire \line_cache[252][3] ;
 wire \line_cache[252][4] ;
 wire \line_cache[252][5] ;
 wire \line_cache[252][6] ;
 wire \line_cache[252][7] ;
 wire \line_cache[253][0] ;
 wire \line_cache[253][1] ;
 wire \line_cache[253][2] ;
 wire \line_cache[253][3] ;
 wire \line_cache[253][4] ;
 wire \line_cache[253][5] ;
 wire \line_cache[253][6] ;
 wire \line_cache[253][7] ;
 wire \line_cache[254][0] ;
 wire \line_cache[254][1] ;
 wire \line_cache[254][2] ;
 wire \line_cache[254][3] ;
 wire \line_cache[254][4] ;
 wire \line_cache[254][5] ;
 wire \line_cache[254][6] ;
 wire \line_cache[254][7] ;
 wire \line_cache[255][0] ;
 wire \line_cache[255][1] ;
 wire \line_cache[255][2] ;
 wire \line_cache[255][3] ;
 wire \line_cache[255][4] ;
 wire \line_cache[255][5] ;
 wire \line_cache[255][6] ;
 wire \line_cache[255][7] ;
 wire \line_cache[256][0] ;
 wire \line_cache[256][1] ;
 wire \line_cache[256][2] ;
 wire \line_cache[256][3] ;
 wire \line_cache[256][4] ;
 wire \line_cache[256][5] ;
 wire \line_cache[256][6] ;
 wire \line_cache[256][7] ;
 wire \line_cache[257][0] ;
 wire \line_cache[257][1] ;
 wire \line_cache[257][2] ;
 wire \line_cache[257][3] ;
 wire \line_cache[257][4] ;
 wire \line_cache[257][5] ;
 wire \line_cache[257][6] ;
 wire \line_cache[257][7] ;
 wire \line_cache[258][0] ;
 wire \line_cache[258][1] ;
 wire \line_cache[258][2] ;
 wire \line_cache[258][3] ;
 wire \line_cache[258][4] ;
 wire \line_cache[258][5] ;
 wire \line_cache[258][6] ;
 wire \line_cache[258][7] ;
 wire \line_cache[259][0] ;
 wire \line_cache[259][1] ;
 wire \line_cache[259][2] ;
 wire \line_cache[259][3] ;
 wire \line_cache[259][4] ;
 wire \line_cache[259][5] ;
 wire \line_cache[259][6] ;
 wire \line_cache[259][7] ;
 wire \line_cache[25][0] ;
 wire \line_cache[25][1] ;
 wire \line_cache[25][2] ;
 wire \line_cache[25][3] ;
 wire \line_cache[25][4] ;
 wire \line_cache[25][5] ;
 wire \line_cache[25][6] ;
 wire \line_cache[25][7] ;
 wire \line_cache[260][0] ;
 wire \line_cache[260][1] ;
 wire \line_cache[260][2] ;
 wire \line_cache[260][3] ;
 wire \line_cache[260][4] ;
 wire \line_cache[260][5] ;
 wire \line_cache[260][6] ;
 wire \line_cache[260][7] ;
 wire \line_cache[261][0] ;
 wire \line_cache[261][1] ;
 wire \line_cache[261][2] ;
 wire \line_cache[261][3] ;
 wire \line_cache[261][4] ;
 wire \line_cache[261][5] ;
 wire \line_cache[261][6] ;
 wire \line_cache[261][7] ;
 wire \line_cache[262][0] ;
 wire \line_cache[262][1] ;
 wire \line_cache[262][2] ;
 wire \line_cache[262][3] ;
 wire \line_cache[262][4] ;
 wire \line_cache[262][5] ;
 wire \line_cache[262][6] ;
 wire \line_cache[262][7] ;
 wire \line_cache[263][0] ;
 wire \line_cache[263][1] ;
 wire \line_cache[263][2] ;
 wire \line_cache[263][3] ;
 wire \line_cache[263][4] ;
 wire \line_cache[263][5] ;
 wire \line_cache[263][6] ;
 wire \line_cache[263][7] ;
 wire \line_cache[264][0] ;
 wire \line_cache[264][1] ;
 wire \line_cache[264][2] ;
 wire \line_cache[264][3] ;
 wire \line_cache[264][4] ;
 wire \line_cache[264][5] ;
 wire \line_cache[264][6] ;
 wire \line_cache[264][7] ;
 wire \line_cache[265][0] ;
 wire \line_cache[265][1] ;
 wire \line_cache[265][2] ;
 wire \line_cache[265][3] ;
 wire \line_cache[265][4] ;
 wire \line_cache[265][5] ;
 wire \line_cache[265][6] ;
 wire \line_cache[265][7] ;
 wire \line_cache[266][0] ;
 wire \line_cache[266][1] ;
 wire \line_cache[266][2] ;
 wire \line_cache[266][3] ;
 wire \line_cache[266][4] ;
 wire \line_cache[266][5] ;
 wire \line_cache[266][6] ;
 wire \line_cache[266][7] ;
 wire \line_cache[267][0] ;
 wire \line_cache[267][1] ;
 wire \line_cache[267][2] ;
 wire \line_cache[267][3] ;
 wire \line_cache[267][4] ;
 wire \line_cache[267][5] ;
 wire \line_cache[267][6] ;
 wire \line_cache[267][7] ;
 wire \line_cache[268][0] ;
 wire \line_cache[268][1] ;
 wire \line_cache[268][2] ;
 wire \line_cache[268][3] ;
 wire \line_cache[268][4] ;
 wire \line_cache[268][5] ;
 wire \line_cache[268][6] ;
 wire \line_cache[268][7] ;
 wire \line_cache[269][0] ;
 wire \line_cache[269][1] ;
 wire \line_cache[269][2] ;
 wire \line_cache[269][3] ;
 wire \line_cache[269][4] ;
 wire \line_cache[269][5] ;
 wire \line_cache[269][6] ;
 wire \line_cache[269][7] ;
 wire \line_cache[26][0] ;
 wire \line_cache[26][1] ;
 wire \line_cache[26][2] ;
 wire \line_cache[26][3] ;
 wire \line_cache[26][4] ;
 wire \line_cache[26][5] ;
 wire \line_cache[26][6] ;
 wire \line_cache[26][7] ;
 wire \line_cache[270][0] ;
 wire \line_cache[270][1] ;
 wire \line_cache[270][2] ;
 wire \line_cache[270][3] ;
 wire \line_cache[270][4] ;
 wire \line_cache[270][5] ;
 wire \line_cache[270][6] ;
 wire \line_cache[270][7] ;
 wire \line_cache[271][0] ;
 wire \line_cache[271][1] ;
 wire \line_cache[271][2] ;
 wire \line_cache[271][3] ;
 wire \line_cache[271][4] ;
 wire \line_cache[271][5] ;
 wire \line_cache[271][6] ;
 wire \line_cache[271][7] ;
 wire \line_cache[272][0] ;
 wire \line_cache[272][1] ;
 wire \line_cache[272][2] ;
 wire \line_cache[272][3] ;
 wire \line_cache[272][4] ;
 wire \line_cache[272][5] ;
 wire \line_cache[272][6] ;
 wire \line_cache[272][7] ;
 wire \line_cache[273][0] ;
 wire \line_cache[273][1] ;
 wire \line_cache[273][2] ;
 wire \line_cache[273][3] ;
 wire \line_cache[273][4] ;
 wire \line_cache[273][5] ;
 wire \line_cache[273][6] ;
 wire \line_cache[273][7] ;
 wire \line_cache[274][0] ;
 wire \line_cache[274][1] ;
 wire \line_cache[274][2] ;
 wire \line_cache[274][3] ;
 wire \line_cache[274][4] ;
 wire \line_cache[274][5] ;
 wire \line_cache[274][6] ;
 wire \line_cache[274][7] ;
 wire \line_cache[275][0] ;
 wire \line_cache[275][1] ;
 wire \line_cache[275][2] ;
 wire \line_cache[275][3] ;
 wire \line_cache[275][4] ;
 wire \line_cache[275][5] ;
 wire \line_cache[275][6] ;
 wire \line_cache[275][7] ;
 wire \line_cache[276][0] ;
 wire \line_cache[276][1] ;
 wire \line_cache[276][2] ;
 wire \line_cache[276][3] ;
 wire \line_cache[276][4] ;
 wire \line_cache[276][5] ;
 wire \line_cache[276][6] ;
 wire \line_cache[276][7] ;
 wire \line_cache[277][0] ;
 wire \line_cache[277][1] ;
 wire \line_cache[277][2] ;
 wire \line_cache[277][3] ;
 wire \line_cache[277][4] ;
 wire \line_cache[277][5] ;
 wire \line_cache[277][6] ;
 wire \line_cache[277][7] ;
 wire \line_cache[278][0] ;
 wire \line_cache[278][1] ;
 wire \line_cache[278][2] ;
 wire \line_cache[278][3] ;
 wire \line_cache[278][4] ;
 wire \line_cache[278][5] ;
 wire \line_cache[278][6] ;
 wire \line_cache[278][7] ;
 wire \line_cache[279][0] ;
 wire \line_cache[279][1] ;
 wire \line_cache[279][2] ;
 wire \line_cache[279][3] ;
 wire \line_cache[279][4] ;
 wire \line_cache[279][5] ;
 wire \line_cache[279][6] ;
 wire \line_cache[279][7] ;
 wire \line_cache[27][0] ;
 wire \line_cache[27][1] ;
 wire \line_cache[27][2] ;
 wire \line_cache[27][3] ;
 wire \line_cache[27][4] ;
 wire \line_cache[27][5] ;
 wire \line_cache[27][6] ;
 wire \line_cache[27][7] ;
 wire \line_cache[280][0] ;
 wire \line_cache[280][1] ;
 wire \line_cache[280][2] ;
 wire \line_cache[280][3] ;
 wire \line_cache[280][4] ;
 wire \line_cache[280][5] ;
 wire \line_cache[280][6] ;
 wire \line_cache[280][7] ;
 wire \line_cache[281][0] ;
 wire \line_cache[281][1] ;
 wire \line_cache[281][2] ;
 wire \line_cache[281][3] ;
 wire \line_cache[281][4] ;
 wire \line_cache[281][5] ;
 wire \line_cache[281][6] ;
 wire \line_cache[281][7] ;
 wire \line_cache[282][0] ;
 wire \line_cache[282][1] ;
 wire \line_cache[282][2] ;
 wire \line_cache[282][3] ;
 wire \line_cache[282][4] ;
 wire \line_cache[282][5] ;
 wire \line_cache[282][6] ;
 wire \line_cache[282][7] ;
 wire \line_cache[283][0] ;
 wire \line_cache[283][1] ;
 wire \line_cache[283][2] ;
 wire \line_cache[283][3] ;
 wire \line_cache[283][4] ;
 wire \line_cache[283][5] ;
 wire \line_cache[283][6] ;
 wire \line_cache[283][7] ;
 wire \line_cache[284][0] ;
 wire \line_cache[284][1] ;
 wire \line_cache[284][2] ;
 wire \line_cache[284][3] ;
 wire \line_cache[284][4] ;
 wire \line_cache[284][5] ;
 wire \line_cache[284][6] ;
 wire \line_cache[284][7] ;
 wire \line_cache[285][0] ;
 wire \line_cache[285][1] ;
 wire \line_cache[285][2] ;
 wire \line_cache[285][3] ;
 wire \line_cache[285][4] ;
 wire \line_cache[285][5] ;
 wire \line_cache[285][6] ;
 wire \line_cache[285][7] ;
 wire \line_cache[286][0] ;
 wire \line_cache[286][1] ;
 wire \line_cache[286][2] ;
 wire \line_cache[286][3] ;
 wire \line_cache[286][4] ;
 wire \line_cache[286][5] ;
 wire \line_cache[286][6] ;
 wire \line_cache[286][7] ;
 wire \line_cache[287][0] ;
 wire \line_cache[287][1] ;
 wire \line_cache[287][2] ;
 wire \line_cache[287][3] ;
 wire \line_cache[287][4] ;
 wire \line_cache[287][5] ;
 wire \line_cache[287][6] ;
 wire \line_cache[287][7] ;
 wire \line_cache[288][0] ;
 wire \line_cache[288][1] ;
 wire \line_cache[288][2] ;
 wire \line_cache[288][3] ;
 wire \line_cache[288][4] ;
 wire \line_cache[288][5] ;
 wire \line_cache[288][6] ;
 wire \line_cache[288][7] ;
 wire \line_cache[289][0] ;
 wire \line_cache[289][1] ;
 wire \line_cache[289][2] ;
 wire \line_cache[289][3] ;
 wire \line_cache[289][4] ;
 wire \line_cache[289][5] ;
 wire \line_cache[289][6] ;
 wire \line_cache[289][7] ;
 wire \line_cache[28][0] ;
 wire \line_cache[28][1] ;
 wire \line_cache[28][2] ;
 wire \line_cache[28][3] ;
 wire \line_cache[28][4] ;
 wire \line_cache[28][5] ;
 wire \line_cache[28][6] ;
 wire \line_cache[28][7] ;
 wire \line_cache[290][0] ;
 wire \line_cache[290][1] ;
 wire \line_cache[290][2] ;
 wire \line_cache[290][3] ;
 wire \line_cache[290][4] ;
 wire \line_cache[290][5] ;
 wire \line_cache[290][6] ;
 wire \line_cache[290][7] ;
 wire \line_cache[291][0] ;
 wire \line_cache[291][1] ;
 wire \line_cache[291][2] ;
 wire \line_cache[291][3] ;
 wire \line_cache[291][4] ;
 wire \line_cache[291][5] ;
 wire \line_cache[291][6] ;
 wire \line_cache[291][7] ;
 wire \line_cache[292][0] ;
 wire \line_cache[292][1] ;
 wire \line_cache[292][2] ;
 wire \line_cache[292][3] ;
 wire \line_cache[292][4] ;
 wire \line_cache[292][5] ;
 wire \line_cache[292][6] ;
 wire \line_cache[292][7] ;
 wire \line_cache[293][0] ;
 wire \line_cache[293][1] ;
 wire \line_cache[293][2] ;
 wire \line_cache[293][3] ;
 wire \line_cache[293][4] ;
 wire \line_cache[293][5] ;
 wire \line_cache[293][6] ;
 wire \line_cache[293][7] ;
 wire \line_cache[294][0] ;
 wire \line_cache[294][1] ;
 wire \line_cache[294][2] ;
 wire \line_cache[294][3] ;
 wire \line_cache[294][4] ;
 wire \line_cache[294][5] ;
 wire \line_cache[294][6] ;
 wire \line_cache[294][7] ;
 wire \line_cache[295][0] ;
 wire \line_cache[295][1] ;
 wire \line_cache[295][2] ;
 wire \line_cache[295][3] ;
 wire \line_cache[295][4] ;
 wire \line_cache[295][5] ;
 wire \line_cache[295][6] ;
 wire \line_cache[295][7] ;
 wire \line_cache[296][0] ;
 wire \line_cache[296][1] ;
 wire \line_cache[296][2] ;
 wire \line_cache[296][3] ;
 wire \line_cache[296][4] ;
 wire \line_cache[296][5] ;
 wire \line_cache[296][6] ;
 wire \line_cache[296][7] ;
 wire \line_cache[297][0] ;
 wire \line_cache[297][1] ;
 wire \line_cache[297][2] ;
 wire \line_cache[297][3] ;
 wire \line_cache[297][4] ;
 wire \line_cache[297][5] ;
 wire \line_cache[297][6] ;
 wire \line_cache[297][7] ;
 wire \line_cache[298][0] ;
 wire \line_cache[298][1] ;
 wire \line_cache[298][2] ;
 wire \line_cache[298][3] ;
 wire \line_cache[298][4] ;
 wire \line_cache[298][5] ;
 wire \line_cache[298][6] ;
 wire \line_cache[298][7] ;
 wire \line_cache[299][0] ;
 wire \line_cache[299][1] ;
 wire \line_cache[299][2] ;
 wire \line_cache[299][3] ;
 wire \line_cache[299][4] ;
 wire \line_cache[299][5] ;
 wire \line_cache[299][6] ;
 wire \line_cache[299][7] ;
 wire \line_cache[29][0] ;
 wire \line_cache[29][1] ;
 wire \line_cache[29][2] ;
 wire \line_cache[29][3] ;
 wire \line_cache[29][4] ;
 wire \line_cache[29][5] ;
 wire \line_cache[29][6] ;
 wire \line_cache[29][7] ;
 wire \line_cache[2][0] ;
 wire \line_cache[2][1] ;
 wire \line_cache[2][2] ;
 wire \line_cache[2][3] ;
 wire \line_cache[2][4] ;
 wire \line_cache[2][5] ;
 wire \line_cache[2][6] ;
 wire \line_cache[2][7] ;
 wire \line_cache[300][0] ;
 wire \line_cache[300][1] ;
 wire \line_cache[300][2] ;
 wire \line_cache[300][3] ;
 wire \line_cache[300][4] ;
 wire \line_cache[300][5] ;
 wire \line_cache[300][6] ;
 wire \line_cache[300][7] ;
 wire \line_cache[301][0] ;
 wire \line_cache[301][1] ;
 wire \line_cache[301][2] ;
 wire \line_cache[301][3] ;
 wire \line_cache[301][4] ;
 wire \line_cache[301][5] ;
 wire \line_cache[301][6] ;
 wire \line_cache[301][7] ;
 wire \line_cache[302][0] ;
 wire \line_cache[302][1] ;
 wire \line_cache[302][2] ;
 wire \line_cache[302][3] ;
 wire \line_cache[302][4] ;
 wire \line_cache[302][5] ;
 wire \line_cache[302][6] ;
 wire \line_cache[302][7] ;
 wire \line_cache[303][0] ;
 wire \line_cache[303][1] ;
 wire \line_cache[303][2] ;
 wire \line_cache[303][3] ;
 wire \line_cache[303][4] ;
 wire \line_cache[303][5] ;
 wire \line_cache[303][6] ;
 wire \line_cache[303][7] ;
 wire \line_cache[304][0] ;
 wire \line_cache[304][1] ;
 wire \line_cache[304][2] ;
 wire \line_cache[304][3] ;
 wire \line_cache[304][4] ;
 wire \line_cache[304][5] ;
 wire \line_cache[304][6] ;
 wire \line_cache[304][7] ;
 wire \line_cache[305][0] ;
 wire \line_cache[305][1] ;
 wire \line_cache[305][2] ;
 wire \line_cache[305][3] ;
 wire \line_cache[305][4] ;
 wire \line_cache[305][5] ;
 wire \line_cache[305][6] ;
 wire \line_cache[305][7] ;
 wire \line_cache[306][0] ;
 wire \line_cache[306][1] ;
 wire \line_cache[306][2] ;
 wire \line_cache[306][3] ;
 wire \line_cache[306][4] ;
 wire \line_cache[306][5] ;
 wire \line_cache[306][6] ;
 wire \line_cache[306][7] ;
 wire \line_cache[307][0] ;
 wire \line_cache[307][1] ;
 wire \line_cache[307][2] ;
 wire \line_cache[307][3] ;
 wire \line_cache[307][4] ;
 wire \line_cache[307][5] ;
 wire \line_cache[307][6] ;
 wire \line_cache[307][7] ;
 wire \line_cache[308][0] ;
 wire \line_cache[308][1] ;
 wire \line_cache[308][2] ;
 wire \line_cache[308][3] ;
 wire \line_cache[308][4] ;
 wire \line_cache[308][5] ;
 wire \line_cache[308][6] ;
 wire \line_cache[308][7] ;
 wire \line_cache[309][0] ;
 wire \line_cache[309][1] ;
 wire \line_cache[309][2] ;
 wire \line_cache[309][3] ;
 wire \line_cache[309][4] ;
 wire \line_cache[309][5] ;
 wire \line_cache[309][6] ;
 wire \line_cache[309][7] ;
 wire \line_cache[30][0] ;
 wire \line_cache[30][1] ;
 wire \line_cache[30][2] ;
 wire \line_cache[30][3] ;
 wire \line_cache[30][4] ;
 wire \line_cache[30][5] ;
 wire \line_cache[30][6] ;
 wire \line_cache[30][7] ;
 wire \line_cache[310][0] ;
 wire \line_cache[310][1] ;
 wire \line_cache[310][2] ;
 wire \line_cache[310][3] ;
 wire \line_cache[310][4] ;
 wire \line_cache[310][5] ;
 wire \line_cache[310][6] ;
 wire \line_cache[310][7] ;
 wire \line_cache[311][0] ;
 wire \line_cache[311][1] ;
 wire \line_cache[311][2] ;
 wire \line_cache[311][3] ;
 wire \line_cache[311][4] ;
 wire \line_cache[311][5] ;
 wire \line_cache[311][6] ;
 wire \line_cache[311][7] ;
 wire \line_cache[312][0] ;
 wire \line_cache[312][1] ;
 wire \line_cache[312][2] ;
 wire \line_cache[312][3] ;
 wire \line_cache[312][4] ;
 wire \line_cache[312][5] ;
 wire \line_cache[312][6] ;
 wire \line_cache[312][7] ;
 wire \line_cache[313][0] ;
 wire \line_cache[313][1] ;
 wire \line_cache[313][2] ;
 wire \line_cache[313][3] ;
 wire \line_cache[313][4] ;
 wire \line_cache[313][5] ;
 wire \line_cache[313][6] ;
 wire \line_cache[313][7] ;
 wire \line_cache[314][0] ;
 wire \line_cache[314][1] ;
 wire \line_cache[314][2] ;
 wire \line_cache[314][3] ;
 wire \line_cache[314][4] ;
 wire \line_cache[314][5] ;
 wire \line_cache[314][6] ;
 wire \line_cache[314][7] ;
 wire \line_cache[315][0] ;
 wire \line_cache[315][1] ;
 wire \line_cache[315][2] ;
 wire \line_cache[315][3] ;
 wire \line_cache[315][4] ;
 wire \line_cache[315][5] ;
 wire \line_cache[315][6] ;
 wire \line_cache[315][7] ;
 wire \line_cache[316][0] ;
 wire \line_cache[316][1] ;
 wire \line_cache[316][2] ;
 wire \line_cache[316][3] ;
 wire \line_cache[316][4] ;
 wire \line_cache[316][5] ;
 wire \line_cache[316][6] ;
 wire \line_cache[316][7] ;
 wire \line_cache[317][0] ;
 wire \line_cache[317][1] ;
 wire \line_cache[317][2] ;
 wire \line_cache[317][3] ;
 wire \line_cache[317][4] ;
 wire \line_cache[317][5] ;
 wire \line_cache[317][6] ;
 wire \line_cache[317][7] ;
 wire \line_cache[318][0] ;
 wire \line_cache[318][1] ;
 wire \line_cache[318][2] ;
 wire \line_cache[318][3] ;
 wire \line_cache[318][4] ;
 wire \line_cache[318][5] ;
 wire \line_cache[318][6] ;
 wire \line_cache[318][7] ;
 wire \line_cache[319][0] ;
 wire \line_cache[319][1] ;
 wire \line_cache[319][2] ;
 wire \line_cache[319][3] ;
 wire \line_cache[319][4] ;
 wire \line_cache[319][5] ;
 wire \line_cache[319][6] ;
 wire \line_cache[319][7] ;
 wire \line_cache[31][0] ;
 wire \line_cache[31][1] ;
 wire \line_cache[31][2] ;
 wire \line_cache[31][3] ;
 wire \line_cache[31][4] ;
 wire \line_cache[31][5] ;
 wire \line_cache[31][6] ;
 wire \line_cache[31][7] ;
 wire \line_cache[32][0] ;
 wire \line_cache[32][1] ;
 wire \line_cache[32][2] ;
 wire \line_cache[32][3] ;
 wire \line_cache[32][4] ;
 wire \line_cache[32][5] ;
 wire \line_cache[32][6] ;
 wire \line_cache[32][7] ;
 wire \line_cache[33][0] ;
 wire \line_cache[33][1] ;
 wire \line_cache[33][2] ;
 wire \line_cache[33][3] ;
 wire \line_cache[33][4] ;
 wire \line_cache[33][5] ;
 wire \line_cache[33][6] ;
 wire \line_cache[33][7] ;
 wire \line_cache[34][0] ;
 wire \line_cache[34][1] ;
 wire \line_cache[34][2] ;
 wire \line_cache[34][3] ;
 wire \line_cache[34][4] ;
 wire \line_cache[34][5] ;
 wire \line_cache[34][6] ;
 wire \line_cache[34][7] ;
 wire \line_cache[35][0] ;
 wire \line_cache[35][1] ;
 wire \line_cache[35][2] ;
 wire \line_cache[35][3] ;
 wire \line_cache[35][4] ;
 wire \line_cache[35][5] ;
 wire \line_cache[35][6] ;
 wire \line_cache[35][7] ;
 wire \line_cache[36][0] ;
 wire \line_cache[36][1] ;
 wire \line_cache[36][2] ;
 wire \line_cache[36][3] ;
 wire \line_cache[36][4] ;
 wire \line_cache[36][5] ;
 wire \line_cache[36][6] ;
 wire \line_cache[36][7] ;
 wire \line_cache[37][0] ;
 wire \line_cache[37][1] ;
 wire \line_cache[37][2] ;
 wire \line_cache[37][3] ;
 wire \line_cache[37][4] ;
 wire \line_cache[37][5] ;
 wire \line_cache[37][6] ;
 wire \line_cache[37][7] ;
 wire \line_cache[38][0] ;
 wire \line_cache[38][1] ;
 wire \line_cache[38][2] ;
 wire \line_cache[38][3] ;
 wire \line_cache[38][4] ;
 wire \line_cache[38][5] ;
 wire \line_cache[38][6] ;
 wire \line_cache[38][7] ;
 wire \line_cache[39][0] ;
 wire \line_cache[39][1] ;
 wire \line_cache[39][2] ;
 wire \line_cache[39][3] ;
 wire \line_cache[39][4] ;
 wire \line_cache[39][5] ;
 wire \line_cache[39][6] ;
 wire \line_cache[39][7] ;
 wire \line_cache[3][0] ;
 wire \line_cache[3][1] ;
 wire \line_cache[3][2] ;
 wire \line_cache[3][3] ;
 wire \line_cache[3][4] ;
 wire \line_cache[3][5] ;
 wire \line_cache[3][6] ;
 wire \line_cache[3][7] ;
 wire \line_cache[40][0] ;
 wire \line_cache[40][1] ;
 wire \line_cache[40][2] ;
 wire \line_cache[40][3] ;
 wire \line_cache[40][4] ;
 wire \line_cache[40][5] ;
 wire \line_cache[40][6] ;
 wire \line_cache[40][7] ;
 wire \line_cache[41][0] ;
 wire \line_cache[41][1] ;
 wire \line_cache[41][2] ;
 wire \line_cache[41][3] ;
 wire \line_cache[41][4] ;
 wire \line_cache[41][5] ;
 wire \line_cache[41][6] ;
 wire \line_cache[41][7] ;
 wire \line_cache[42][0] ;
 wire \line_cache[42][1] ;
 wire \line_cache[42][2] ;
 wire \line_cache[42][3] ;
 wire \line_cache[42][4] ;
 wire \line_cache[42][5] ;
 wire \line_cache[42][6] ;
 wire \line_cache[42][7] ;
 wire \line_cache[43][0] ;
 wire \line_cache[43][1] ;
 wire \line_cache[43][2] ;
 wire \line_cache[43][3] ;
 wire \line_cache[43][4] ;
 wire \line_cache[43][5] ;
 wire \line_cache[43][6] ;
 wire \line_cache[43][7] ;
 wire \line_cache[44][0] ;
 wire \line_cache[44][1] ;
 wire \line_cache[44][2] ;
 wire \line_cache[44][3] ;
 wire \line_cache[44][4] ;
 wire \line_cache[44][5] ;
 wire \line_cache[44][6] ;
 wire \line_cache[44][7] ;
 wire \line_cache[45][0] ;
 wire \line_cache[45][1] ;
 wire \line_cache[45][2] ;
 wire \line_cache[45][3] ;
 wire \line_cache[45][4] ;
 wire \line_cache[45][5] ;
 wire \line_cache[45][6] ;
 wire \line_cache[45][7] ;
 wire \line_cache[46][0] ;
 wire \line_cache[46][1] ;
 wire \line_cache[46][2] ;
 wire \line_cache[46][3] ;
 wire \line_cache[46][4] ;
 wire \line_cache[46][5] ;
 wire \line_cache[46][6] ;
 wire \line_cache[46][7] ;
 wire \line_cache[47][0] ;
 wire \line_cache[47][1] ;
 wire \line_cache[47][2] ;
 wire \line_cache[47][3] ;
 wire \line_cache[47][4] ;
 wire \line_cache[47][5] ;
 wire \line_cache[47][6] ;
 wire \line_cache[47][7] ;
 wire \line_cache[48][0] ;
 wire \line_cache[48][1] ;
 wire \line_cache[48][2] ;
 wire \line_cache[48][3] ;
 wire \line_cache[48][4] ;
 wire \line_cache[48][5] ;
 wire \line_cache[48][6] ;
 wire \line_cache[48][7] ;
 wire \line_cache[49][0] ;
 wire \line_cache[49][1] ;
 wire \line_cache[49][2] ;
 wire \line_cache[49][3] ;
 wire \line_cache[49][4] ;
 wire \line_cache[49][5] ;
 wire \line_cache[49][6] ;
 wire \line_cache[49][7] ;
 wire \line_cache[4][0] ;
 wire \line_cache[4][1] ;
 wire \line_cache[4][2] ;
 wire \line_cache[4][3] ;
 wire \line_cache[4][4] ;
 wire \line_cache[4][5] ;
 wire \line_cache[4][6] ;
 wire \line_cache[4][7] ;
 wire \line_cache[50][0] ;
 wire \line_cache[50][1] ;
 wire \line_cache[50][2] ;
 wire \line_cache[50][3] ;
 wire \line_cache[50][4] ;
 wire \line_cache[50][5] ;
 wire \line_cache[50][6] ;
 wire \line_cache[50][7] ;
 wire \line_cache[51][0] ;
 wire \line_cache[51][1] ;
 wire \line_cache[51][2] ;
 wire \line_cache[51][3] ;
 wire \line_cache[51][4] ;
 wire \line_cache[51][5] ;
 wire \line_cache[51][6] ;
 wire \line_cache[51][7] ;
 wire \line_cache[52][0] ;
 wire \line_cache[52][1] ;
 wire \line_cache[52][2] ;
 wire \line_cache[52][3] ;
 wire \line_cache[52][4] ;
 wire \line_cache[52][5] ;
 wire \line_cache[52][6] ;
 wire \line_cache[52][7] ;
 wire \line_cache[53][0] ;
 wire \line_cache[53][1] ;
 wire \line_cache[53][2] ;
 wire \line_cache[53][3] ;
 wire \line_cache[53][4] ;
 wire \line_cache[53][5] ;
 wire \line_cache[53][6] ;
 wire \line_cache[53][7] ;
 wire \line_cache[54][0] ;
 wire \line_cache[54][1] ;
 wire \line_cache[54][2] ;
 wire \line_cache[54][3] ;
 wire \line_cache[54][4] ;
 wire \line_cache[54][5] ;
 wire \line_cache[54][6] ;
 wire \line_cache[54][7] ;
 wire \line_cache[55][0] ;
 wire \line_cache[55][1] ;
 wire \line_cache[55][2] ;
 wire \line_cache[55][3] ;
 wire \line_cache[55][4] ;
 wire \line_cache[55][5] ;
 wire \line_cache[55][6] ;
 wire \line_cache[55][7] ;
 wire \line_cache[56][0] ;
 wire \line_cache[56][1] ;
 wire \line_cache[56][2] ;
 wire \line_cache[56][3] ;
 wire \line_cache[56][4] ;
 wire \line_cache[56][5] ;
 wire \line_cache[56][6] ;
 wire \line_cache[56][7] ;
 wire \line_cache[57][0] ;
 wire \line_cache[57][1] ;
 wire \line_cache[57][2] ;
 wire \line_cache[57][3] ;
 wire \line_cache[57][4] ;
 wire \line_cache[57][5] ;
 wire \line_cache[57][6] ;
 wire \line_cache[57][7] ;
 wire \line_cache[58][0] ;
 wire \line_cache[58][1] ;
 wire \line_cache[58][2] ;
 wire \line_cache[58][3] ;
 wire \line_cache[58][4] ;
 wire \line_cache[58][5] ;
 wire \line_cache[58][6] ;
 wire \line_cache[58][7] ;
 wire \line_cache[59][0] ;
 wire \line_cache[59][1] ;
 wire \line_cache[59][2] ;
 wire \line_cache[59][3] ;
 wire \line_cache[59][4] ;
 wire \line_cache[59][5] ;
 wire \line_cache[59][6] ;
 wire \line_cache[59][7] ;
 wire \line_cache[5][0] ;
 wire \line_cache[5][1] ;
 wire \line_cache[5][2] ;
 wire \line_cache[5][3] ;
 wire \line_cache[5][4] ;
 wire \line_cache[5][5] ;
 wire \line_cache[5][6] ;
 wire \line_cache[5][7] ;
 wire \line_cache[60][0] ;
 wire \line_cache[60][1] ;
 wire \line_cache[60][2] ;
 wire \line_cache[60][3] ;
 wire \line_cache[60][4] ;
 wire \line_cache[60][5] ;
 wire \line_cache[60][6] ;
 wire \line_cache[60][7] ;
 wire \line_cache[61][0] ;
 wire \line_cache[61][1] ;
 wire \line_cache[61][2] ;
 wire \line_cache[61][3] ;
 wire \line_cache[61][4] ;
 wire \line_cache[61][5] ;
 wire \line_cache[61][6] ;
 wire \line_cache[61][7] ;
 wire \line_cache[62][0] ;
 wire \line_cache[62][1] ;
 wire \line_cache[62][2] ;
 wire \line_cache[62][3] ;
 wire \line_cache[62][4] ;
 wire \line_cache[62][5] ;
 wire \line_cache[62][6] ;
 wire \line_cache[62][7] ;
 wire \line_cache[63][0] ;
 wire \line_cache[63][1] ;
 wire \line_cache[63][2] ;
 wire \line_cache[63][3] ;
 wire \line_cache[63][4] ;
 wire \line_cache[63][5] ;
 wire \line_cache[63][6] ;
 wire \line_cache[63][7] ;
 wire \line_cache[64][0] ;
 wire \line_cache[64][1] ;
 wire \line_cache[64][2] ;
 wire \line_cache[64][3] ;
 wire \line_cache[64][4] ;
 wire \line_cache[64][5] ;
 wire \line_cache[64][6] ;
 wire \line_cache[64][7] ;
 wire \line_cache[65][0] ;
 wire \line_cache[65][1] ;
 wire \line_cache[65][2] ;
 wire \line_cache[65][3] ;
 wire \line_cache[65][4] ;
 wire \line_cache[65][5] ;
 wire \line_cache[65][6] ;
 wire \line_cache[65][7] ;
 wire \line_cache[66][0] ;
 wire \line_cache[66][1] ;
 wire \line_cache[66][2] ;
 wire \line_cache[66][3] ;
 wire \line_cache[66][4] ;
 wire \line_cache[66][5] ;
 wire \line_cache[66][6] ;
 wire \line_cache[66][7] ;
 wire \line_cache[67][0] ;
 wire \line_cache[67][1] ;
 wire \line_cache[67][2] ;
 wire \line_cache[67][3] ;
 wire \line_cache[67][4] ;
 wire \line_cache[67][5] ;
 wire \line_cache[67][6] ;
 wire \line_cache[67][7] ;
 wire \line_cache[68][0] ;
 wire \line_cache[68][1] ;
 wire \line_cache[68][2] ;
 wire \line_cache[68][3] ;
 wire \line_cache[68][4] ;
 wire \line_cache[68][5] ;
 wire \line_cache[68][6] ;
 wire \line_cache[68][7] ;
 wire \line_cache[69][0] ;
 wire \line_cache[69][1] ;
 wire \line_cache[69][2] ;
 wire \line_cache[69][3] ;
 wire \line_cache[69][4] ;
 wire \line_cache[69][5] ;
 wire \line_cache[69][6] ;
 wire \line_cache[69][7] ;
 wire \line_cache[6][0] ;
 wire \line_cache[6][1] ;
 wire \line_cache[6][2] ;
 wire \line_cache[6][3] ;
 wire \line_cache[6][4] ;
 wire \line_cache[6][5] ;
 wire \line_cache[6][6] ;
 wire \line_cache[6][7] ;
 wire \line_cache[70][0] ;
 wire \line_cache[70][1] ;
 wire \line_cache[70][2] ;
 wire \line_cache[70][3] ;
 wire \line_cache[70][4] ;
 wire \line_cache[70][5] ;
 wire \line_cache[70][6] ;
 wire \line_cache[70][7] ;
 wire \line_cache[71][0] ;
 wire \line_cache[71][1] ;
 wire \line_cache[71][2] ;
 wire \line_cache[71][3] ;
 wire \line_cache[71][4] ;
 wire \line_cache[71][5] ;
 wire \line_cache[71][6] ;
 wire \line_cache[71][7] ;
 wire \line_cache[72][0] ;
 wire \line_cache[72][1] ;
 wire \line_cache[72][2] ;
 wire \line_cache[72][3] ;
 wire \line_cache[72][4] ;
 wire \line_cache[72][5] ;
 wire \line_cache[72][6] ;
 wire \line_cache[72][7] ;
 wire \line_cache[73][0] ;
 wire \line_cache[73][1] ;
 wire \line_cache[73][2] ;
 wire \line_cache[73][3] ;
 wire \line_cache[73][4] ;
 wire \line_cache[73][5] ;
 wire \line_cache[73][6] ;
 wire \line_cache[73][7] ;
 wire \line_cache[74][0] ;
 wire \line_cache[74][1] ;
 wire \line_cache[74][2] ;
 wire \line_cache[74][3] ;
 wire \line_cache[74][4] ;
 wire \line_cache[74][5] ;
 wire \line_cache[74][6] ;
 wire \line_cache[74][7] ;
 wire \line_cache[75][0] ;
 wire \line_cache[75][1] ;
 wire \line_cache[75][2] ;
 wire \line_cache[75][3] ;
 wire \line_cache[75][4] ;
 wire \line_cache[75][5] ;
 wire \line_cache[75][6] ;
 wire \line_cache[75][7] ;
 wire \line_cache[76][0] ;
 wire \line_cache[76][1] ;
 wire \line_cache[76][2] ;
 wire \line_cache[76][3] ;
 wire \line_cache[76][4] ;
 wire \line_cache[76][5] ;
 wire \line_cache[76][6] ;
 wire \line_cache[76][7] ;
 wire \line_cache[77][0] ;
 wire \line_cache[77][1] ;
 wire \line_cache[77][2] ;
 wire \line_cache[77][3] ;
 wire \line_cache[77][4] ;
 wire \line_cache[77][5] ;
 wire \line_cache[77][6] ;
 wire \line_cache[77][7] ;
 wire \line_cache[78][0] ;
 wire \line_cache[78][1] ;
 wire \line_cache[78][2] ;
 wire \line_cache[78][3] ;
 wire \line_cache[78][4] ;
 wire \line_cache[78][5] ;
 wire \line_cache[78][6] ;
 wire \line_cache[78][7] ;
 wire \line_cache[79][0] ;
 wire \line_cache[79][1] ;
 wire \line_cache[79][2] ;
 wire \line_cache[79][3] ;
 wire \line_cache[79][4] ;
 wire \line_cache[79][5] ;
 wire \line_cache[79][6] ;
 wire \line_cache[79][7] ;
 wire \line_cache[7][0] ;
 wire \line_cache[7][1] ;
 wire \line_cache[7][2] ;
 wire \line_cache[7][3] ;
 wire \line_cache[7][4] ;
 wire \line_cache[7][5] ;
 wire \line_cache[7][6] ;
 wire \line_cache[7][7] ;
 wire \line_cache[80][0] ;
 wire \line_cache[80][1] ;
 wire \line_cache[80][2] ;
 wire \line_cache[80][3] ;
 wire \line_cache[80][4] ;
 wire \line_cache[80][5] ;
 wire \line_cache[80][6] ;
 wire \line_cache[80][7] ;
 wire \line_cache[81][0] ;
 wire \line_cache[81][1] ;
 wire \line_cache[81][2] ;
 wire \line_cache[81][3] ;
 wire \line_cache[81][4] ;
 wire \line_cache[81][5] ;
 wire \line_cache[81][6] ;
 wire \line_cache[81][7] ;
 wire \line_cache[82][0] ;
 wire \line_cache[82][1] ;
 wire \line_cache[82][2] ;
 wire \line_cache[82][3] ;
 wire \line_cache[82][4] ;
 wire \line_cache[82][5] ;
 wire \line_cache[82][6] ;
 wire \line_cache[82][7] ;
 wire \line_cache[83][0] ;
 wire \line_cache[83][1] ;
 wire \line_cache[83][2] ;
 wire \line_cache[83][3] ;
 wire \line_cache[83][4] ;
 wire \line_cache[83][5] ;
 wire \line_cache[83][6] ;
 wire \line_cache[83][7] ;
 wire \line_cache[84][0] ;
 wire \line_cache[84][1] ;
 wire \line_cache[84][2] ;
 wire \line_cache[84][3] ;
 wire \line_cache[84][4] ;
 wire \line_cache[84][5] ;
 wire \line_cache[84][6] ;
 wire \line_cache[84][7] ;
 wire \line_cache[85][0] ;
 wire \line_cache[85][1] ;
 wire \line_cache[85][2] ;
 wire \line_cache[85][3] ;
 wire \line_cache[85][4] ;
 wire \line_cache[85][5] ;
 wire \line_cache[85][6] ;
 wire \line_cache[85][7] ;
 wire \line_cache[86][0] ;
 wire \line_cache[86][1] ;
 wire \line_cache[86][2] ;
 wire \line_cache[86][3] ;
 wire \line_cache[86][4] ;
 wire \line_cache[86][5] ;
 wire \line_cache[86][6] ;
 wire \line_cache[86][7] ;
 wire \line_cache[87][0] ;
 wire \line_cache[87][1] ;
 wire \line_cache[87][2] ;
 wire \line_cache[87][3] ;
 wire \line_cache[87][4] ;
 wire \line_cache[87][5] ;
 wire \line_cache[87][6] ;
 wire \line_cache[87][7] ;
 wire \line_cache[88][0] ;
 wire \line_cache[88][1] ;
 wire \line_cache[88][2] ;
 wire \line_cache[88][3] ;
 wire \line_cache[88][4] ;
 wire \line_cache[88][5] ;
 wire \line_cache[88][6] ;
 wire \line_cache[88][7] ;
 wire \line_cache[89][0] ;
 wire \line_cache[89][1] ;
 wire \line_cache[89][2] ;
 wire \line_cache[89][3] ;
 wire \line_cache[89][4] ;
 wire \line_cache[89][5] ;
 wire \line_cache[89][6] ;
 wire \line_cache[89][7] ;
 wire \line_cache[8][0] ;
 wire \line_cache[8][1] ;
 wire \line_cache[8][2] ;
 wire \line_cache[8][3] ;
 wire \line_cache[8][4] ;
 wire \line_cache[8][5] ;
 wire \line_cache[8][6] ;
 wire \line_cache[8][7] ;
 wire \line_cache[90][0] ;
 wire \line_cache[90][1] ;
 wire \line_cache[90][2] ;
 wire \line_cache[90][3] ;
 wire \line_cache[90][4] ;
 wire \line_cache[90][5] ;
 wire \line_cache[90][6] ;
 wire \line_cache[90][7] ;
 wire \line_cache[91][0] ;
 wire \line_cache[91][1] ;
 wire \line_cache[91][2] ;
 wire \line_cache[91][3] ;
 wire \line_cache[91][4] ;
 wire \line_cache[91][5] ;
 wire \line_cache[91][6] ;
 wire \line_cache[91][7] ;
 wire \line_cache[92][0] ;
 wire \line_cache[92][1] ;
 wire \line_cache[92][2] ;
 wire \line_cache[92][3] ;
 wire \line_cache[92][4] ;
 wire \line_cache[92][5] ;
 wire \line_cache[92][6] ;
 wire \line_cache[92][7] ;
 wire \line_cache[93][0] ;
 wire \line_cache[93][1] ;
 wire \line_cache[93][2] ;
 wire \line_cache[93][3] ;
 wire \line_cache[93][4] ;
 wire \line_cache[93][5] ;
 wire \line_cache[93][6] ;
 wire \line_cache[93][7] ;
 wire \line_cache[94][0] ;
 wire \line_cache[94][1] ;
 wire \line_cache[94][2] ;
 wire \line_cache[94][3] ;
 wire \line_cache[94][4] ;
 wire \line_cache[94][5] ;
 wire \line_cache[94][6] ;
 wire \line_cache[94][7] ;
 wire \line_cache[95][0] ;
 wire \line_cache[95][1] ;
 wire \line_cache[95][2] ;
 wire \line_cache[95][3] ;
 wire \line_cache[95][4] ;
 wire \line_cache[95][5] ;
 wire \line_cache[95][6] ;
 wire \line_cache[95][7] ;
 wire \line_cache[96][0] ;
 wire \line_cache[96][1] ;
 wire \line_cache[96][2] ;
 wire \line_cache[96][3] ;
 wire \line_cache[96][4] ;
 wire \line_cache[96][5] ;
 wire \line_cache[96][6] ;
 wire \line_cache[96][7] ;
 wire \line_cache[97][0] ;
 wire \line_cache[97][1] ;
 wire \line_cache[97][2] ;
 wire \line_cache[97][3] ;
 wire \line_cache[97][4] ;
 wire \line_cache[97][5] ;
 wire \line_cache[97][6] ;
 wire \line_cache[97][7] ;
 wire \line_cache[98][0] ;
 wire \line_cache[98][1] ;
 wire \line_cache[98][2] ;
 wire \line_cache[98][3] ;
 wire \line_cache[98][4] ;
 wire \line_cache[98][5] ;
 wire \line_cache[98][6] ;
 wire \line_cache[98][7] ;
 wire \line_cache[99][0] ;
 wire \line_cache[99][1] ;
 wire \line_cache[99][2] ;
 wire \line_cache[99][3] ;
 wire \line_cache[99][4] ;
 wire \line_cache[99][5] ;
 wire \line_cache[99][6] ;
 wire \line_cache[99][7] ;
 wire \line_cache[9][0] ;
 wire \line_cache[9][1] ;
 wire \line_cache[9][2] ;
 wire \line_cache[9][3] ;
 wire \line_cache[9][4] ;
 wire \line_cache[9][5] ;
 wire \line_cache[9][6] ;
 wire \line_cache[9][7] ;
 wire \line_cache_idx[2] ;
 wire \line_cache_idx[3] ;
 wire \line_cache_idx[4] ;
 wire \line_cache_idx[5] ;
 wire \line_cache_idx[6] ;
 wire \line_cache_idx[7] ;
 wire \line_cache_idx[8] ;
 wire \line_cache_idx[9] ;
 wire \line_double_counter[0] ;
 wire \line_double_counter[1] ;
 wire \line_double_counter[2] ;
 wire \line_double_counter[3] ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net247;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net249;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net254;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net256;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net259;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net26;
 wire net260;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net263;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net264;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net268;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net269;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net274;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net297;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net298;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net303;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net304;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net305;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net306;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net31;
 wire net310;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net311;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net315;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net317;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net324;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net325;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net329;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net33;
 wire net330;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net332;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net336;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net339;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net342;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net344;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net345;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net346;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net354;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net355;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net356;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net357;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net358;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net359;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net360;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net361;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net362;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net363;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net364;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net365;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net366;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net367;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net368;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net369;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net37;
 wire net370;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net38;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net39;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4;
 wire net40;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net407;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net408;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net409;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net41;
 wire net410;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net411;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net412;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net413;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net414;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net415;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net416;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net417;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net418;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net419;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net42;
 wire net420;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net421;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net422;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net423;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net424;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net425;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net426;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net427;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net428;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net429;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net43;
 wire net430;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net431;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net432;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net433;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \pixel_double_counter[0] ;
 wire \pixel_double_counter[1] ;
 wire \pixel_double_counter[2] ;
 wire \pixel_double_counter[3] ;
 wire \prescaler[0] ;
 wire \prescaler[1] ;
 wire \prescaler[2] ;
 wire \prescaler[3] ;
 wire \prescaler_counter[0] ;
 wire \prescaler_counter[1] ;
 wire \prescaler_counter[2] ;
 wire \prescaler_counter[3] ;
 wire \prescaler_counter[4] ;
 wire \prescaler_counter[5] ;
 wire \prescaler_counter[6] ;
 wire \prescaler_counter[7] ;
 wire \prescaler_counter[8] ;
 wire \res_h_active[0] ;
 wire \res_h_active[1] ;
 wire \res_h_active[2] ;
 wire \res_h_active[3] ;
 wire \res_h_active[4] ;
 wire \res_h_active[5] ;
 wire \res_h_active[6] ;
 wire \res_h_active[7] ;
 wire \res_h_active[8] ;
 wire \res_h_counter[0] ;
 wire \res_h_counter[1] ;
 wire \res_h_counter[2] ;
 wire \res_h_counter[3] ;
 wire \res_h_counter[4] ;
 wire \res_h_counter[5] ;
 wire \res_h_counter[6] ;
 wire \res_h_counter[7] ;
 wire \res_h_counter[8] ;
 wire \res_h_counter[9] ;
 wire \res_v_active[0] ;
 wire \res_v_active[1] ;
 wire \res_v_active[2] ;
 wire \res_v_active[3] ;
 wire \res_v_active[4] ;
 wire \res_v_active[5] ;
 wire \res_v_active[6] ;
 wire \res_v_active[7] ;
 wire \res_v_counter[0] ;
 wire \res_v_counter[1] ;
 wire \res_v_counter[2] ;
 wire \res_v_counter[3] ;
 wire \res_v_counter[4] ;
 wire \res_v_counter[5] ;
 wire \res_v_counter[6] ;
 wire \res_v_counter[7] ;
 wire \res_v_counter[8] ;
 wire \res_v_counter[9] ;
 wire \resolution[0] ;
 wire \resolution[1] ;
 wire \resolution[2] ;
 wire \resolution[3] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_10503_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_10503_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_10503_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_06249_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_06618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_06909_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_06935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_07105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_07231_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_07525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__A (.DIODE(\base_h_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__A (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__B (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__B2 (.DIODE(_08547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__A (.DIODE(\base_v_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__B (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B1 (.DIODE(_08547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B2 (.DIODE(_08604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__B (.DIODE(_08613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A (.DIODE(_08632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__A (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__A (.DIODE(_08661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__A (.DIODE(_08722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__B1 (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__11862__A (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11862__B (.DIODE(_08726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__B (.DIODE(net2713));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__B1_N (.DIODE(_08771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A1 (.DIODE(net4316));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A2 (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__B1 (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__C1 (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__D1 (.DIODE(net2713));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__A (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__B (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__A1 (.DIODE(_08661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11927__A (.DIODE(_08726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__A (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A1 (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A2 (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A3 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__B1 (.DIODE(net4215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__A1 (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__A2 (.DIODE(net2713));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__B1 (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__C1 (.DIODE(_08726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__A (.DIODE(_08632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__B (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__A1 (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__A2 (.DIODE(net2713));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__B1 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__B (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A1 (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__B1 (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__B (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__A1 (.DIODE(\base_h_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__B (.DIODE(\base_h_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12113__A1_N (.DIODE(\base_h_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__B (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__A (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__B (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12124__B (.DIODE(\base_h_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__B (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__B (.DIODE(\base_v_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A (.DIODE(\base_v_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__B (.DIODE(\base_v_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A (.DIODE(_09163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__A (.DIODE(_09168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A (.DIODE(_09179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A (.DIODE(_09184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__A (.DIODE(_09187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__A (.DIODE(_08726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__B (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12350__A (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12367__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__A (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__A (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__A2 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12381__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12383__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__A (.DIODE(_09238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12410__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__A (.DIODE(_09252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12415__A (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A2 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__12433__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__A (.DIODE(_09276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__B (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__A2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A (.DIODE(_09283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__A (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__B (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A (.DIODE(_09293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__B2 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__A (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__B (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__A (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__A (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__B2 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__A1 (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A3 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A3 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A3 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A3 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__A (.DIODE(_09331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12516__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A3 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__A (.DIODE(_09337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12530__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__C (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__A (.DIODE(_09353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12554__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12571__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__A1 (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__A2_N (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A2_N (.DIODE(_09310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A1 (.DIODE(_09303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12640__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12651__A (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__A2 (.DIODE(_09273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A (.DIODE(_09381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__B (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__A (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__B2 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12692__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__A (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12700__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12702__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12727__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__C (.DIODE(_09360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A (.DIODE(_09391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12766__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12769__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__12769__B (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__A2 (.DIODE(_09504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12775__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A (.DIODE(_09509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A1 (.DIODE(_09412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__A (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A2 (.DIODE(_09432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A (.DIODE(_09484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A (.DIODE(_09513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12862__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12865__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12870__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12877__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12879__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12887__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__C (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12889__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__A (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__B (.DIODE(_09199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__A (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12907__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12909__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12915__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__A1 (.DIODE(_09527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12932__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12947__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12949__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__A2 (.DIODE(_09552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__A (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13001__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__A (.DIODE(_09622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13052__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__C (.DIODE(_09602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13076__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13086__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13088__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__A1 (.DIODE(_09613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13092__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13101__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13112__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__A (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__A (.DIODE(_09376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__A (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A3 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__A3 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__A2 (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A3 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__A3 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A3 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A3 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13179__A (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A3 (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__A3 (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__A3 (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__A3 (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13210__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__A (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__C (.DIODE(_09696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__A1 (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13216__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__A2_N (.DIODE(_09743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__B (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__A3 (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__A (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__A (.DIODE(_09717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13228__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13247__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13250__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13263__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__A1 (.DIODE(_09712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13276__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13277__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13278__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__A (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13280__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13282__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__A (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13284__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13286__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13291__A (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13291__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13291__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13292__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__A (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13297__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13298__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13299__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13300__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__A2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13307__A (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13307__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13307__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13309__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13313__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13314__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__A (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13317__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__B1 (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13373__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13385__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13411__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__A2_N (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13414__A2_N (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13414__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13416__A2_N (.DIODE(_09861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13416__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13426__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13427__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13429__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13443__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13446__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13449__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13451__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13455__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13474__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13478__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13479__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13482__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13484__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__A2 (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13488__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__A2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13495__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__A (.DIODE(_09926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13503__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13505__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13507__B (.DIODE(_09982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__B1 (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13519__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13519__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__A3 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__A3 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13527__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13527__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13527__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__A (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__B1 (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__B1 (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13536__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13536__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__A3 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__B1 (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13544__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13544__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__A1 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__A3 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13546__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13548__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13548__A3 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13550__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__C (.DIODE(_09833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__A3 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13569__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13569__A3 (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13574__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13579__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13579__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13579__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__A3 (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A (.DIODE(_09985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__A1 (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__A2_N (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__A2_N (.DIODE(_09993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__B (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__A3 (.DIODE(_09990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13604__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13605__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13606__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13608__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13614__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13618__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__A2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13629__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13631__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13632__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13633__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13634__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13635__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13638__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13639__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13640__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13641__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13642__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13643__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13643__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13643__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13644__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13646__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13648__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13648__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13648__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__A2 (.DIODE(_09977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13650__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13655__A2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13661__A2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13663__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13667__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13669__A (.DIODE(_10042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13669__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13669__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13672__A2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13678__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13682__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__A (.DIODE(_10097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13693__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13696__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13702__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13717__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13719__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13725__A2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13728__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13731__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13738__A2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13744__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13750__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13756__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13758__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__13760__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13765__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__A (.DIODE(_09716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13777__A2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13779__A (.DIODE(_09283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13781__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13784__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13787__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13788__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13789__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13790__A (.DIODE(_09733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13791__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13795__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13796__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13801__A1 (.DIODE(_10010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__A (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13805__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13812__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13814__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13815__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13816__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__A2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13823__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13825__A (.DIODE(_09331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13827__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13829__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13830__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13832__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13834__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13835__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__A (.DIODE(_09238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13838__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13841__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13843__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13844__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13845__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13845__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13845__C (.DIODE(_10019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13846__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13848__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13849__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13850__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13850__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13850__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13851__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13853__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13856__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13866__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13868__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13868__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13868__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13869__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13871__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__A (.DIODE(_10174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13874__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13877__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13878__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13879__B1 (.DIODE(_09298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13880__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13881__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13882__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13886__B (.DIODE(_10233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13888__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13888__B (.DIODE(_10235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__A (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__B (.DIODE(_10235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__B2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13900__A (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__A3 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__B (.DIODE(_10235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13903__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13904__A1 (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13904__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13905__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13906__A1 (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13906__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13907__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13908__A (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13909__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13909__B1 (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13909__B2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13910__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13911__A (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__A3 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13913__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13916__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13917__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__13919__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13919__B1 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13919__B2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__A (.DIODE(_09331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__B1 (.DIODE(_10259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__B2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13929__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13930__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13932__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13935__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13936__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__A (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__A3 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13940__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13941__A (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13942__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13942__A2 (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13942__A3 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13943__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13944__A1 (.DIODE(_10181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13946__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__B1 (.DIODE(_10273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__B2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13949__A2 (.DIODE(_10083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13950__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13951__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__13952__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13952__B1 (.DIODE(_10276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13952__B2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13953__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13954__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13955__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13956__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13957__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13959__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13960__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13961__A (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__A2 (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__A3 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13963__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__A (.DIODE(_09283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__B1 (.DIODE(_10285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__B2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13966__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13967__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13971__A (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13972__A2_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13972__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13972__B2 (.DIODE(_10235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13973__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__A (.DIODE(_10291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__A (.DIODE(_10233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13978__B (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13979__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__B2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13986__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13986__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13987__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13987__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13989__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13989__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13998__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13998__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14000__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14004__A (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14006__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14010__A (.DIODE(_09331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14011__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14014__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14014__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14015__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14015__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14020__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14028__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14028__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__A1 (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14030__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__A3 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14036__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14040__A3 (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14042__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14046__B2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14048__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14048__B (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14049__A3 (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14050__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14050__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14051__A3 (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__A (.DIODE(_09283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14057__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__A (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14063__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14065__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__B1 (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__B1 (.DIODE(_10300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__A (.DIODE(_10355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__A (.DIODE(_10233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__B (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14079__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14090__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14092__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14095__B2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14097__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14100__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14103__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14106__B2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14110__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14112__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14112__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14114__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__B2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14119__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14120__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14120__C (.DIODE(_10210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14122__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14124__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14125__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14127__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14130__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14132__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__A (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14136__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14138__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14141__B2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14143__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14145__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14146__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14148__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14152__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14153__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14155__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14156__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__14160__A (.DIODE(_10233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14160__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14161__A (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14162__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14164__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14165__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14167__B2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14170__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14172__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14174__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14175__B2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14177__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14179__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14181__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14183__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14185__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14187__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14188__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14190__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14191__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14193__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14194__B2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14196__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14197__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14199__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14201__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14202__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14204__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14206__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14208__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14210__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__B2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14213__B (.DIODE(_09351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14215__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14216__B2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14218__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14219__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14221__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14223__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14224__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14226__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14228__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14230__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14233__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14237__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14239__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14240__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14243__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__14245__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14247__A (.DIODE(_09509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14247__B (.DIODE(_10466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14250__A (.DIODE(_10467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14250__B (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14251__B (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14253__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14255__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14256__A (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14257__B1 (.DIODE(_10475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14259__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14261__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14263__B1 (.DIODE(_10479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14264__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14265__B (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14265__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14268__B1 (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14271__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14271__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14273__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14274__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__A (.DIODE(_10226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14277__B1 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14278__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14279__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__B1 (.DIODE(_10259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14281__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14283__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14285__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14286__A (.DIODE(_09337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__B1 (.DIODE(_10493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14288__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14288__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14290__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14292__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14294__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14295__A (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14296__B1 (.DIODE(_10498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14299__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__14300__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14300__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14302__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14303__A (.DIODE(_09353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14304__B1 (.DIODE(_10503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14306__B1 (.DIODE(_10273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14309__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__B1 (.DIODE(_10276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14311__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14311__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14313__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14315__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14315__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14317__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__B1 (.DIODE(_10285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14321__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14321__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14324__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14326__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14327__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__14329__A (.DIODE(_10467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14329__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14331__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14335__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14338__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14339__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14339__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14341__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14343__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14343__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14344__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14345__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14346__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14346__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14351__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14352__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14352__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14354__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14354__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14355__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14356__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14359__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14360__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14360__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14362__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14363__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14363__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14365__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14366__A (.DIODE(_09230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14367__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14368__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14369__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14370__A (.DIODE(_09236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14371__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14372__A (.DIODE(_10350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14373__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14373__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14375__A (.DIODE(_09243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14376__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14377__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14378__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14379__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14379__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14380__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14381__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14382__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14385__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14386__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14387__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14389__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14389__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__B (.DIODE(_09266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14392__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14394__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14394__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14403__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14403__A2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14406__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14406__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14409__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14409__A2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14412__A1 (.DIODE(_10524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14412__A2 (.DIODE(_09504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14414__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14415__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14416__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14417__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14418__A (.DIODE(_10467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14418__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14420__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14424__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14424__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14425__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14426__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14426__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14427__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14428__A (.DIODE(_09188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14428__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14429__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14430__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14432__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14434__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__14435__A (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14437__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14438__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14438__C (.DIODE(_10480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14439__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14440__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14440__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14441__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14442__A (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14444__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14446__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14446__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14449__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14452__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14455__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14458__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14459__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14460__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14460__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14461__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14461__A3 (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14466__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14468__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14468__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14469__A1 (.DIODE(_10542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14469__A3 (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14470__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14471__B (.DIODE(_09345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14472__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14473__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14474__A (.DIODE(_09253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14474__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__A3 (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14477__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14478__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14478__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14479__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14479__A3 (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14481__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14483__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14485__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14486__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14487__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14488__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14490__B (.DIODE(_09274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14491__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__A (.DIODE(_09277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__B (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__A3 (.DIODE(_10579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14495__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14496__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14498__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14501__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14502__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14504__A2 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14505__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14506__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14507__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14509__A (.DIODE(_10467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14509__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14511__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14515__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14515__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__B1 (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14521__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14522__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14525__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14526__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14527__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14528__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14529__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14531__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14533__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__A (.DIODE(_09216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14537__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14538__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14539__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14541__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14542__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14544__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A3 (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__A (.DIODE(_09233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14548__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14548__A3 (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14549__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14549__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__A3 (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14554__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14555__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14555__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__A3 (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14560__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14563__A (.DIODE(_09252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__A3 (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14567__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14568__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14569__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14571__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14574__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14575__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14576__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14577__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14581__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14582__A (.DIODE(_09276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14583__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14583__B (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14584__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14584__A3 (.DIODE(_10638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14585__B (.DIODE(_09369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14586__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14587__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14588__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14590__B (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14591__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14593__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14593__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14594__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14595__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14598__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14599__A (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14599__B (.DIODE(_10466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14600__A (.DIODE(_10691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14600__B (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14601__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14604__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14606__A (.DIODE(_09185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__A (.DIODE(_09187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14609__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14610__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14610__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14611__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14612__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14613__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14613__B1 (.DIODE(_10479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__A1 (.DIODE(_10611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14616__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14617__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14617__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14618__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14619__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14620__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14621__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14621__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14624__A1 (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14624__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14625__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14625__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__14626__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14627__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14627__B1 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14628__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14629__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14629__B1 (.DIODE(_10259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14630__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14631__A3 (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__A1 (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14633__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14633__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14636__A1 (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14636__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__A2 (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14638__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14640__A1 (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14640__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14641__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14641__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__14642__A (.DIODE(_10488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14643__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14643__B1 (.DIODE(_10498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14644__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14646__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14646__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14648__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14650__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14651__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__B1 (.DIODE(_10273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14655__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__B1 (.DIODE(_10276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14657__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14657__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14659__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14660__A (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__B1 (.DIODE(_10727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__14663__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14663__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14665__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14666__A2_N (.DIODE(_10694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14666__B1 (.DIODE(_10285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14667__A1 (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14667__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__A2 (.DIODE(_09373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14669__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14669__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14671__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A (.DIODE(_10691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14678__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14680__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14683__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14687__A (.DIODE(_09184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14688__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14688__B (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14689__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14690__A (.DIODE(_10619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14691__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14695__A2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14701__A2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14703__A (.DIODE(_09209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14704__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14705__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14705__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14706__A1 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14706__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14707__A (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14709__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14710__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14710__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14715__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14717__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14718__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14718__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14719__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14720__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14721__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14721__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14722__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14723__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14723__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14725__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14730__A2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14732__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14732__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14733__A1 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14733__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14735__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14738__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14740__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14741__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14741__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14743__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14745__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14745__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14746__A1 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14746__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14751__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14754__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14757__A1 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14757__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14759__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14762__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__14764__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14764__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__A1 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__A2 (.DIODE(_10646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14766__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__A2_N (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14768__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14769__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14769__A3 (.DIODE(_10745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14770__A (.DIODE(_10691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14770__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14773__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14777__A2 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14780__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__A3 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14782__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14783__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14783__A3 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14784__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14785__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14785__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14786__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14786__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14787__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14787__C (.DIODE(_10687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14789__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14790__B (.DIODE(_09395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14791__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14791__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14792__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14793__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14794__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14796__B (.DIODE(_09326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14797__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14797__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14798__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14799__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14799__A3 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14800__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14801__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14804__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14806__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14807__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14807__A3 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14808__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14809__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14809__A3 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14810__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14811__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14812__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14814__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14815__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14816__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__14819__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14820__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14820__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14821__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14822__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14824__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14825__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14827__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14830__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14831__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14833__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14834__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14836__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14837__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14839__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14840__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14840__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14841__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14842__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14843__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14844__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14844__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14845__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14846__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14848__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__14849__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14850__A1 (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14850__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14852__A2 (.DIODE(_09504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14854__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__A2_N (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14856__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__A2_N (.DIODE(_10806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14858__A (.DIODE(_10691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14858__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14860__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14861__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14864__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14865__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14868__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__A1 (.DIODE(_10759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__A3 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14870__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14871__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14872__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14873__A3 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14874__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14875__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14875__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14876__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14877__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14877__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14878__A (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14879__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14880__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14882__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14883__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14884__A3 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14885__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__14886__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14887__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14887__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14888__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14889__A3 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14890__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14891__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14893__A (.DIODE(_10814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14894__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14896__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14898__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14900__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14902__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14903__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14904__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14906__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14908__A (.DIODE(_09246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14910__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14911__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14911__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14912__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14913__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14915__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14916__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14916__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14917__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14918__A2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14920__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14921__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14923__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14924__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14924__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14925__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14926__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14929__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14929__A2 (.DIODE(_10809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14931__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14933__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14934__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14935__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14935__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14936__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14937__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14939__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14941__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14942__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14942__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14943__A1 (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14943__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14944__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14945__A2_N (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14945__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14946__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14947__A2_N (.DIODE(_10862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14947__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14948__A (.DIODE(_10466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14948__B (.DIODE(_09982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14949__A (.DIODE(_10912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14949__B (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14952__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14955__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14957__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14959__B (.DIODE(_09463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14959__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14961__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14961__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14963__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14964__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14966__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14968__A (.DIODE(_10395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14969__B2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14971__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14971__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14973__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14975__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14976__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14977__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14980__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14981__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14983__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14985__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14986__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14988__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14990__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14991__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14993__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14996__B2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14998__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14998__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15000__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15002__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15002__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15004__A (.DIODE(_09260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15006__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15007__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15009__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15010__B2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15012__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15013__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15015__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15016__B2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15018__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15019__B2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15024__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15025__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15027__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15028__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15031__B2 (.DIODE(_09504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15033__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15034__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15036__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15037__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__15039__A (.DIODE(_10912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15039__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15041__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15042__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15045__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15046__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15049__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15051__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15052__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15055__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15056__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15058__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15058__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15059__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15061__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15063__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15065__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15066__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15068__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15070__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15071__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15073__A (.DIODE(_10884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15078__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15080__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15082__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15082__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15084__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15087__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15089__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15089__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15090__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15091__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15093__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15095__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15097__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15098__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15099__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15100__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15102__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15105__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15108__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15110__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15110__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15111__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15113__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15115__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15115__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15116__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15118__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15121__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__15123__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15123__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15124__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15125__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15126__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15127__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__A (.DIODE(_10912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15131__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15132__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15136__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15139__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15140__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15141__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15142__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15143__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__15144__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15144__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15145__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15147__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15150__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15153__A2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15156__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15159__A2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15162__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15165__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15167__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15168__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15169__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15170__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15171__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15172__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15173__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15173__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15174__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15175__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15176__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15177__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15178__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15179__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15179__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15180__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15182__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15184__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15184__C (.DIODE(_10908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15185__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15186__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15188__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15190__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15196__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15198__A (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15199__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15199__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15200__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15202__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15204__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15204__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15205__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15207__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15209__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15209__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15210__A2 (.DIODE(_10903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15212__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15212__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15213__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15214__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15215__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15216__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15217__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15218__A (.DIODE(_10912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15218__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15220__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15222__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15226__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15232__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15235__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15238__A2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15241__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15245__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15248__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15251__A2 (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15254__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15259__A (.DIODE(_10349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15261__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15264__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15267__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15271__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15274__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15277__A2 (.DIODE(_09414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15283__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15286__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15288__A (.DIODE(_09353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15290__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15293__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15296__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15302__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15305__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15310__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15311__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15312__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15313__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15316__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__15318__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15319__A2 (.DIODE(_09504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15321__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15322__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15323__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15324__B1 (.DIODE(_09442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15326__A (.DIODE(_11161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15326__B (.DIODE(_09168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__A (.DIODE(_11162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__B (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15328__B (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15331__A (.DIODE(_09181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15332__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15333__A (.DIODE(_10721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15335__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15336__B1 (.DIODE(_10475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15337__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15338__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15339__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15339__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15340__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15342__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15343__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15344__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15345__B1 (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15346__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15347__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15348__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15348__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15349__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15350__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15351__A1 (.DIODE(_11009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15352__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15353__B1 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15354__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15355__B1 (.DIODE(_10259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15356__A1 (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15356__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15357__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15357__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__15358__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15359__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15360__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15361__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15362__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15363__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15363__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15364__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15365__A1 (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15365__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15366__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15366__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__15367__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15368__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15369__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15369__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15370__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15371__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15372__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15373__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15373__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15374__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15375__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15376__B1 (.DIODE(_10503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15377__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15378__B1 (.DIODE(_10273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15379__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15379__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15380__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15381__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15382__B1 (.DIODE(_10276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15383__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15383__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15384__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15385__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15386__B1 (.DIODE(_10727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15387__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15387__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15388__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15389__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15390__B1 (.DIODE(_10285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15391__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15391__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15392__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15393__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15393__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15394__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15395__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15396__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15398__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15399__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__15401__A (.DIODE(_11162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15401__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15403__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15406__A (.DIODE(_09179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15409__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15410__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15411__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15412__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15414__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15415__A2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15417__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15417__C (.DIODE(_11074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15418__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15419__A (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15420__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15421__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15422__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15423__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15424__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15426__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15429__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15430__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15432__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15433__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15434__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15435__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15437__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15438__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15440__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15441__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15442__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15443__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15445__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15446__A1 (.DIODE(_11182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15447__B (.DIODE(_09341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15448__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15449__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15450__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15451__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15452__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15453__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15454__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15455__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15456__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15457__A2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15459__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15460__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15461__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15462__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15463__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15464__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15466__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15467__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15468__A (.DIODE(_11152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15469__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15471__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15472__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15473__A2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15475__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15476__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15477__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15478__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15479__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15480__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15482__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15483__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15484__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15485__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__15487__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15488__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15489__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15490__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15491__A (.DIODE(_11162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15491__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15493__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15494__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15497__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15498__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15500__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15501__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15504__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15505__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15506__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15507__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15510__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15511__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15512__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15515__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15516__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15517__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15518__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15519__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15521__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15523__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15524__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15526__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15527__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15528__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15529__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15530__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15533__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__15534__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15535__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15536__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15537__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15538__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15539__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15540__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15541__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15543__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15544__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15545__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15546__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15547__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15548__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15550__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15551__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15553__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15554__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15555__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15556__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15558__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15559__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15560__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15561__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15562__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15563__A2 (.DIODE(_11082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15564__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15565__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15567__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15568__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15569__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15570__B (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15571__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15573__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15574__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15575__A (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15576__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15577__A (.DIODE(_11162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15577__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15583__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15584__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15585__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15586__A (.DIODE(_11251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15587__A2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15589__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15590__A1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15591__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15592__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15592__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15595__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15596__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15597__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15600__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15602__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15603__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15606__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15607__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15608__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__15610__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15613__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15614__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15616__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15617__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15618__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15619__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15620__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15621__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15622__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15623__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15624__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15626__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15628__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15629__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15630__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15630__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15631__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15632__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15633__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15634__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15634__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15635__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15636__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15637__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15638__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15639__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15641__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15641__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15642__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15644__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15646__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15647__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__15649__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15650__A2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15652__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15653__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15655__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15656__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15658__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15659__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15662__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__15664__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15665__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15666__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15667__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15668__A (.DIODE(_09509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15668__B (.DIODE(_11161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15669__A (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15669__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15670__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15673__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15674__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15675__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15676__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15678__B2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15680__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15681__B2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15683__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15683__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15684__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15685__A (.DIODE(_10931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15686__B2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15688__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__15689__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15689__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15690__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15691__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15692__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15693__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15693__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15694__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15695__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15697__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15700__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15703__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15705__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15706__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15707__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15708__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15709__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15710__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15711__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15711__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15712__A1 (.DIODE(_11345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15714__B2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15716__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15717__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15718__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15719__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15719__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15720__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15721__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15722__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15723__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15723__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15724__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15725__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15726__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15728__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15730__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15730__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15731__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15733__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15735__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15735__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15736__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15737__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15738__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15740__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15743__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15745__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15745__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15746__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15747__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__15748__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15748__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15749__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15750__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15751__A2 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15752__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15753__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15754__A (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15754__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15755__B (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15758__A (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15759__A (.DIODE(_10291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15759__C (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15761__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15761__B1 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15761__B2 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15764__A (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__B2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15768__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15768__B2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15771__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15771__B2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15774__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15774__B2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15777__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15777__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__B2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__B2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15785__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15787__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15787__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15790__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15790__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15793__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15793__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15796__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15796__B2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15799__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15799__B2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15802__A1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15802__B2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15806__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15809__B2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15812__B2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15815__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15815__B2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15818__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15818__B2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15821__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15821__B2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15824__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15824__B2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15830__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15830__B2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15833__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15833__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15835__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15836__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15837__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15837__B2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15840__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15840__B2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15842__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15843__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15843__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15845__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15846__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15846__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15848__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15849__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15849__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15851__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15852__B1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15852__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__15854__A (.DIODE(_11331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15855__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15855__B1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15857__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__A1 (.DIODE(_11436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__A3 (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__B1 (.DIODE(_11432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15860__A (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15860__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15861__B (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15864__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15865__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15866__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15867__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15868__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15869__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15870__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15871__A (.DIODE(_10355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15871__C (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15873__B2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15875__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15875__C (.DIODE(_11328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15876__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15877__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15878__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15878__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15879__A1 (.DIODE(_11408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15880__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15881__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15883__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15883__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15885__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15886__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15888__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15889__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15891__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15892__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15894__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15896__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15897__B2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15899__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15901__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15902__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15904__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15906__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15907__B2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15909__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15910__B2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15912__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15914__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15914__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15916__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15918__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15919__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15921__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15921__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15923__A (.DIODE(_11487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15924__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15926__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15926__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15928__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15930__B2 (.DIODE(_09366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15935__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15938__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15940__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15940__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15942__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15944__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15947__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15949__A (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15949__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15951__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15953__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15957__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15960__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15963__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15966__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15969__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15972__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15974__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15977__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15978__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15981__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15984__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15986__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15988__A (.DIODE(_10864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15989__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15990__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15991__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15992__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15994__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15996__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15997__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15999__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__16001__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16001__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16002__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16004__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16007__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16009__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16010__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16014__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16014__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16015__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16017__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16020__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16022__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16023__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16024__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16026__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16026__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16027__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16028__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16029__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16031__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16032__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16035__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16036__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16037__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16038__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16039__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16040__A (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16040__B (.DIODE(_11161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16041__A (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16041__B (.DIODE(_11620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16043__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16047__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16048__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16049__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16050__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16051__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16052__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16053__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16053__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16054__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16055__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16055__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16056__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16057__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16058__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16059__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16061__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16062__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16063__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16064__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16066__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16067__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16068__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16069__A2 (.DIODE(_10122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16071__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16072__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16074__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16075__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16076__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16077__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16078__A (.DIODE(_10602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16079__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16080__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16080__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16081__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16082__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16083__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16085__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16086__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16087__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16089__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16090__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16092__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16093__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16095__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16096__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16098__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16099__A2 (.DIODE(_10149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16101__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16101__C (.DIODE(_11516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16102__A2 (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16103__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16104__A2 (.DIODE(_10154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16106__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16107__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16108__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16109__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16110__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16111__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16112__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16113__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16115__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16116__A2 (.DIODE(_10164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16118__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16119__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16120__A (.DIODE(_11609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16121__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16123__A (.DIODE(_11174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16124__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16125__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16126__A1 (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16127__A (.DIODE(_11620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16127__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16128__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16131__A (.DIODE(_11620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16132__A (.DIODE(_10291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16132__C (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16134__B1 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16136__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16137__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16139__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16141__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16143__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16145__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16147__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16149__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16152__B2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16154__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16157__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16160__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16163__B2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16165__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16168__B2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16170__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16173__B2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16175__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16177__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16179__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16182__B2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16184__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16187__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16189__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16192__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16195__B2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16197__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16199__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16202__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16204__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16205__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16208__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16210__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16211__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16212__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16214__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16216__A (.DIODE(_11620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16216__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16217__B (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16220__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16222__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16224__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16226__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16228__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16230__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16232__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16234__A (.DIODE(_10355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16234__C (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16236__B2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16238__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16241__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16244__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16247__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16249__A (.DIODE(_10657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16251__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16253__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16254__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16256__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16259__B2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16262__B2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16264__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16266__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16268__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16269__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16269__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16271__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16272__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16273__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16275__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16278__B2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16281__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16283__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16283__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16284__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16285__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16286__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16288__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16291__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16294__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16297__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16299__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16300__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16302__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16303__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__A (.DIODE(_11620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16307__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16308__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16311__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16312__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16312__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16315__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16316__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16317__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16318__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16318__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16320__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16321__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16321__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16323__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16323__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16324__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16328__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16329__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16330__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16331__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16331__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16333__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16334__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16335__A (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16336__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16337__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16337__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16339__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16340__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16340__A2 (.DIODE(_10195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16342__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16343__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16344__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16345__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16346__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16347__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16348__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16349__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16349__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16350__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16351__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16352__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16353__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16354__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16355__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16355__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16356__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16357__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16358__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16359__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16360__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16360__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16362__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16363__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16364__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__16365__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16366__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16366__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16368__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16369__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16369__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16371__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__16372__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16373__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16373__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16375__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16375__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16376__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16377__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16378__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16378__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16380__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16380__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16381__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16382__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__16383__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16384__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16384__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16386__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16388__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16388__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__16390__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16390__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16391__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16392__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16393__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16394__B1 (.DIODE(_10289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16395__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16396__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16397__A (.DIODE(_11161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16397__B (.DIODE(_09982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16398__A (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16398__B (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16400__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16404__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16405__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16405__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16406__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16407__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16407__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16408__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16409__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16409__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16410__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16412__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16415__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16418__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16421__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16424__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16427__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__16430__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16432__A (.DIODE(_09331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16434__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16436__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16437__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16438__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16438__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16439__A (.DIODE(_10767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16440__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16440__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16441__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16443__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16443__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16444__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16444__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16445__A (.DIODE(_10663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16447__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__A3 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16449__B (.DIODE(_10667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16449__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16450__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16450__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16452__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16454__B (.DIODE(_10500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16454__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16455__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16455__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16456__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16457__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16461__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16461__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16462__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16462__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16464__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16466__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16466__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16467__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16467__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16468__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16471__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16474__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16476__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16476__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16477__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16477__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16478__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16478__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16479__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16479__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16480__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16481__A (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16482__A2_N (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16482__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16483__A (.DIODE(_09300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16484__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16485__A (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16485__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16486__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__A (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16490__A (.DIODE(_10291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16490__C (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16492__B1 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16495__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16496__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16497__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16498__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16499__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16499__C (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16501__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16502__B (.DIODE(_10587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16503__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16504__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16505__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16506__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16507__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16509__B2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16512__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16514__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16516__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16518__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16519__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16521__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16522__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16523__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16524__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16525__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16526__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16527__B2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16530__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16532__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16533__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16535__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16537__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__16538__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16540__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16542__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__16543__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16545__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16547__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16548__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16550__B (.DIODE(_10617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16552__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16553__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16555__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16556__B2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16558__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16560__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16562__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16563__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16565__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16566__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16568__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16571__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16574__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16576__A (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16576__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16577__B (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16580__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16582__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16584__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16586__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16588__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16590__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16591__A (.DIODE(_10355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16591__C (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16592__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16594__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16595__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16597__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16599__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16602__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16604__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16605__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16608__B2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16610__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16612__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16614__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16615__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16617__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16621__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16623__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16625__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16627__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16629__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16630__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16632__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__16633__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16635__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16636__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16640__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16642__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16644__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16645__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16647__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16648__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16648__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16650__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16651__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16651__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16652__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16653__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16655__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16658__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16660__A (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16660__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16662__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16663__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16667__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16670__A (.DIODE(_10746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16671__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16673__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16676__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16679__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16682__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16685__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16690__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16691__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16693__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16696__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16699__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16701__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16702__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16703__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16704__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16706__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16708__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16709__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16710__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16711__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16712__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16712__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16713__A2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16715__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16717__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16718__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16718__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16719__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16721__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16724__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16726__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16726__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16727__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16728__A (.DIODE(_11151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16729__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16730__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16732__B (.DIODE(_10679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16732__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16733__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16734__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16735__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16736__B (.DIODE(_10728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16736__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16737__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16738__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16739__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16742__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16744__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16745__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16746__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16747__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16748__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16751__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16751__B (.DIODE(_09168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16752__A (.DIODE(_03164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16752__B (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16753__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16756__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16757__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16758__A (.DIODE(_09184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16759__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16760__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16761__A (.DIODE(_10698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16762__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16763__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16764__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16765__B1 (.DIODE(_10479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16766__A1 (.DIODE(_09302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16766__B2 (.DIODE(_09227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16767__A1 (.DIODE(_09193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16767__A2 (.DIODE(_09321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16768__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16768__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16769__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16770__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16771__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16772__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16772__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16773__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16774__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16775__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16776__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16777__B1 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16778__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16779__B1 (.DIODE(_10259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16780__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16781__A1 (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16782__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16783__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16784__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16785__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16786__B1 (.DIODE(_10493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16787__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16787__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16788__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16789__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16790__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16791__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16792__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16793__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16793__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16794__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16795__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16796__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16798__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16799__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16800__B1 (.DIODE(_10503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16801__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16802__B1 (.DIODE(_10273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16804__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16805__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16806__B1 (.DIODE(_10276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16807__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__16808__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16808__C (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16809__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16810__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16811__B1 (.DIODE(_10727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16812__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16814__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16814__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16816__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__B1 (.DIODE(_10285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16818__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16818__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16819__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16820__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16820__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16822__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16823__A1 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16825__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16826__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16827__A (.DIODE(_03164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16827__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16829__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16830__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16833__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16834__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16836__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16837__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16840__A (.DIODE(_09187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16841__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16842__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16843__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16843__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16844__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16845__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16845__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16846__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16847__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16847__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16848__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16849__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16850__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16852__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16853__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16855__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16856__A2 (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16858__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16859__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16861__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16862__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16864__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16865__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16866__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__A1 (.DIODE(_03183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16868__A (.DIODE(_02772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16869__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16870__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16871__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16872__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16874__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16875__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16876__A (.DIODE(_11002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16877__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16878__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16878__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16879__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16880__A (.DIODE(_10669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16881__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16882__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16883__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16885__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16886__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16887__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16888__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16890__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16890__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16891__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16892__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16893__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16895__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16895__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16896__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16897__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16898__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16900__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16900__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16901__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16902__A (.DIODE(_03150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16903__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16905__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16905__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16906__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16907__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16907__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16908__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16909__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16910__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16911__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16912__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16913__A (.DIODE(_03164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16913__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16915__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16919__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16919__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16920__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16921__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16921__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16922__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16923__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16925__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16926__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16927__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16927__B1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16929__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16929__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16930__A2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16931__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16932__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16932__B1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16934__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16935__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16935__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16936__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16937__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16937__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16938__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16939__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16939__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16940__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16941__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16942__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__16942__B1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16944__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16945__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16945__B1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16947__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16948__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16950__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16950__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16951__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16952__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16952__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16953__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16953__A3 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16954__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16954__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16955__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16955__A3 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16956__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16956__C (.DIODE(_03200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16957__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16958__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16959__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16962__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16962__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16963__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16963__A3 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16964__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16965__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16965__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16966__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16967__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16968__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16970__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16970__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16971__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16972__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16973__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16975__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16976__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16978__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16978__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16979__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16980__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16981__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16983__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16983__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16984__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16985__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16985__B (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16986__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16986__A3 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16987__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16988__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16990__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16991__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16993__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16993__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16994__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16995__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16995__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16996__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16997__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16998__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16999__A (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17000__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17001__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17002__A (.DIODE(_03164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17002__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17004__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17006__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17009__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17010__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17012__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17013__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17015__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17016__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17018__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17019__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17021__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17023__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17026__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17029__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17032__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17035__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__17038__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17041__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17044__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17047__A2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17050__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17054__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17060__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17063__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17066__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17069__A2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17071__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17072__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17073__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17075__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17076__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17078__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17079__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17081__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17082__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17084__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17085__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__17087__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17088__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17090__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17091__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17093__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17094__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17096__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17097__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__17099__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17100__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17102__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17103__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17104__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17105__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17106__A (.DIODE(_09509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17106__B (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17107__A (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17107__B (.DIODE(_03391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17108__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17111__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17112__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17113__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17114__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17115__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17116__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17117__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17119__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17119__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17121__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17123__B (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17125__B2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17127__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17127__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17129__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17131__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17131__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17133__A (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17136__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17139__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17141__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17143__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17146__B2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17148__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17148__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17150__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17153__B2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17156__B2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17159__B2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17161__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17161__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17164__B2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17167__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17169__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17169__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17172__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17174__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17174__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17176__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17179__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17182__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17185__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17187__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17187__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17189__A (.DIODE(_09196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17190__A2 (.DIODE(_10348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17191__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17193__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17194__A (.DIODE(_03391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17194__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17195__B (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17198__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17200__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17202__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17205__A (.DIODE(_03391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17206__A (.DIODE(_10291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17206__C (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17208__B2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17211__B2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17213__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17213__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17216__B2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17218__A (.DIODE(_10930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17220__B2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17223__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17226__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17229__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17231__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17233__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17235__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17237__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17237__C (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17240__B2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17242__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17244__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17245__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17247__A (.DIODE(_09252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17248__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17251__B2 (.DIODE(_09256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17253__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17256__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17258__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17261__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17263__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17265__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17268__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17271__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17273__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17274__B (.DIODE(_10848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17276__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17278__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17279__A1 (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17281__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17283__A (.DIODE(_03391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17283__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17284__B (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17287__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17289__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17291__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17293__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17295__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17298__A (.DIODE(_10355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17298__C (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17302__A (.DIODE(_10872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17304__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17306__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17309__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17312__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17314__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17316__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17319__B2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17321__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17323__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17325__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17328__B2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17330__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17331__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17333__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17336__B2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17339__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17341__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17343__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17344__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17345__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17347__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17349__A (.DIODE(_10681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17351__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17352__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17354__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17355__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17357__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__17358__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17360__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17361__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17363__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17364__A1 (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17366__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17367__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17369__A (.DIODE(_03391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17369__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17371__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17375__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17377__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17379__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17381__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17382__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17383__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17384__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17385__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17386__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17387__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17388__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17389__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17391__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17392__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17394__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17395__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__17397__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17399__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17402__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17405__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17407__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17410__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17412__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17413__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17414__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17416__A2 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17418__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17420__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17421__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17422__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17425__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17427__A (.DIODE(_11010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17430__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17433__A2 (.DIODE(_09425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17436__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17439__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__17441__A (.DIODE(_09276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17442__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17444__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17445__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17447__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17450__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__17453__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17455__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17456__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17457__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17458__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17459__A (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17459__B (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17460__A (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17460__B (.DIODE(_03616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17462__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17466__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17468__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17470__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17472__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17474__B (.DIODE(_11040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17475__A2 (.DIODE(_03278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17476__A (.DIODE(_10645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17477__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17479__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17481__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17482__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17483__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17484__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17486__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17487__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17489__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17494__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17495__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17496__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17497__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17498__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17499__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17500__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17502__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17503__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17504__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17506__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17507__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17509__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17511__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17512__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17513__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17515__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17516__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17518__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17519__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17521__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17522__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17524__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17525__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17527__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17529__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17530__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17531__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17533__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17534__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17536__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17538__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17540__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17541__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17542__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17543__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17543__A3 (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17545__A (.DIODE(_03616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17545__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17546__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17549__A (.DIODE(_11210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17550__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17551__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17552__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17553__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17554__A (.DIODE(_03616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17555__A (.DIODE(_10291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17555__C (.DIODE(_08778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17557__B2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17559__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__17560__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17561__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17562__B2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17564__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17565__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17566__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17567__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17568__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17569__B2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17571__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17572__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17573__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17574__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17576__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17577__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17579__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17580__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17581__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17582__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17583__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17584__A1 (.DIODE(_03632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17585__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17586__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17587__B (.DIODE(_11291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17587__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17589__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17591__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17592__B2 (.DIODE(_09415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17594__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17594__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17596__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17597__B2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17599__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17599__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17601__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17603__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17604__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17606__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17606__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17609__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17611__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17612__B2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17614__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17616__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17616__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17618__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17619__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17621__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17621__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17623__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17623__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17625__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17626__A1 (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17628__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17629__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17631__A (.DIODE(_03616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17631__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17632__B (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17634__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17635__A (.DIODE(_10355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17635__C (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17636__B1 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17638__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17641__B2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17644__B2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17647__B2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17650__B2 (.DIODE(_09201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17653__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17656__B2 (.DIODE(_09398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17659__B2 (.DIODE(_09212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17662__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17665__B2 (.DIODE(_10313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17668__B2 (.DIODE(_10316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17671__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17674__B2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17676__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17679__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17681__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17683__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17685__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17685__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17687__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17689__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17690__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17690__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17692__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17695__B2 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17697__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17697__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17700__B2 (.DIODE(_10335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17702__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17702__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17704__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17707__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17710__B2 (.DIODE(_10342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17712__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17712__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17714__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17714__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17716__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17717__A1 (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17719__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17720__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17722__A (.DIODE(_03616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17722__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17724__A (.DIODE(_08727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17728__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17730__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17732__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17734__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__17734__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17736__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17737__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17738__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17742__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17743__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17745__B (.DIODE(_10874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17745__C (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17747__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17748__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__17750__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17751__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17753__A (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17754__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17756__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17758__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17760__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17762__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17765__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17767__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17769__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17769__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17771__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17773__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17774__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17775__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17777__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17778__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17779__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17780__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17781__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17783__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17783__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17785__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17786__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17788__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17789__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__17791__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17792__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17793__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17794__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17796__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17797__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17799__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17800__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__17802__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17803__A (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17804__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__17804__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17805__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17806__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17807__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17808__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17809__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17810__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17810__B (.DIODE(_09982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17811__A (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17811__B (.DIODE(_10469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17813__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17817__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17818__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17819__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17820__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17821__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17822__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17823__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__17823__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17824__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17825__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17825__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17826__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17827__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17827__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17828__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17829__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17830__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17831__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17833__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17834__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17836__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17837__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17838__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17839__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17841__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17842__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17844__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17845__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17847__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17848__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17849__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17850__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17851__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__17851__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17852__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17853__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17854__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17856__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17857__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17859__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17859__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17860__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17861__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17862__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17863__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17863__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17864__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17865__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17866__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17868__A (.DIODE(_03815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17869__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17871__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17871__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17872__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17873__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17874__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17875__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17877__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17877__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17878__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17879__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17880__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17881__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17881__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17882__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17883__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17884__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17886__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17886__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17887__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17888__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__17888__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17889__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17890__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17891__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17892__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17893__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17894__A (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17894__B (.DIODE(_10292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__B (.DIODE(_10413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17898__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17899__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17900__A (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17902__A (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17903__A (.DIODE(_10291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17903__C (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17905__B2 (.DIODE(_09315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17908__B2 (.DIODE(_09460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17910__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__17910__C (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17911__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17912__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17913__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17913__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17914__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17918__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17919__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17920__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__17920__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17921__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17922__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17923__A1 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17925__B2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17928__B2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17930__A (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17931__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17934__B2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17936__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17939__B2 (.DIODE(_09239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17941__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17943__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17945__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17945__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17948__B2 (.DIODE(_09348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17950__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17950__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17953__B2 (.DIODE(_09354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17956__B2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17958__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17958__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17961__B2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17964__B2 (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17966__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17971__B2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17973__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17973__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17975__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__17975__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17978__A1 (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17980__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17982__A (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17982__B (.DIODE(_10356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17983__B (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17986__A (.DIODE(_10355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17986__C (.DIODE(_08725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17988__B1 (.DIODE(_09451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17993__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17996__B2 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18001__B2 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18003__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18005__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18006__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18006__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18007__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__B2 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18011__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18012__B2 (.DIODE(_09219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18014__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18015__B2 (.DIODE(_09332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18017__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18018__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18019__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18020__B2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18022__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18023__B2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18025__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__18025__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18026__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18027__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18028__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18031__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18032__B2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18035__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18036__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18036__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18037__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18038__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18039__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18040__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18041__B2 (.DIODE(_09263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18043__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18043__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18044__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18045__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18046__B2 (.DIODE(_09269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18048__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18048__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18050__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18052__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18053__B2 (.DIODE(_09280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18055__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18056__B2 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18058__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18059__B2 (.DIODE(_09288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18061__A (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18062__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__18064__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18065__A1 (.DIODE(_09296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18067__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18068__A1 (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18070__A (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18070__B (.DIODE(_10411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18072__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18076__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18077__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18078__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18079__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18080__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18082__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18083__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18085__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__18085__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18086__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18087__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18088__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18090__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18091__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18093__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18094__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18095__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18095__C (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18096__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18097__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18098__A2 (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18100__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18101__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18103__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18104__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18106__A (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18107__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18108__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18109__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18110__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18111__A1 (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18112__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18113__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18115__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18116__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18117__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18118__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18119__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__18121__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18122__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18122__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18123__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18124__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18125__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18126__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18126__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18127__A2 (.DIODE(_03835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18129__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18130__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18133__A (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18134__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18134__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18135__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18136__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18139__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18140__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18141__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__18143__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18144__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18146__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18147__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18149__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18150__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18152__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18152__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18153__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18154__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18154__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18155__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18156__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18157__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18158__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18159__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18161__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18162__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18167__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18168__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18169__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__B1 (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18173__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18174__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18174__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__18174__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18175__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18176__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18177__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18177__B1 (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18179__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18180__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18180__B1 (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18182__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18183__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18183__B1 (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18185__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18186__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18188__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18188__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18189__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18190__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18191__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18193__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18194__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18197__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18198__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18198__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18199__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18200__A (.DIODE(_02845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18200__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18201__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18203__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18204__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18204__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18205__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18206__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18206__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18207__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18208__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18209__A2 (.DIODE(_09249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18211__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18212__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18214__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18214__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18214__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18215__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18216__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18217__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18219__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18220__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18222__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18222__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18222__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18223__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18224__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18225__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18227__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18227__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18227__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18228__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18229__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18229__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18230__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18230__A3 (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18231__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18232__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18233__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18235__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18236__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18238__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18238__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18238__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18239__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18240__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18240__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18240__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18241__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18242__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18243__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18244__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18244__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18245__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18245__A3 (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18247__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18248__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18252__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18253__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18255__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18256__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18257__A1 (.DIODE(_04033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18258__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18258__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__18258__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18259__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18260__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18260__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18260__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18261__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18262__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18263__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18264__A2 (.DIODE(_10869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18266__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18267__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18268__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18269__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18270__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18272__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18273__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18274__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18275__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18277__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18278__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18280__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18281__A2 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18283__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18285__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18286__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18287__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18288__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18290__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18291__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18293__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18294__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18296__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18297__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18298__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18299__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18299__B (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18299__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18300__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18301__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18302__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18304__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18305__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18307__A (.DIODE(_11219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18308__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18308__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18308__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18309__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18310__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18311__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18314__A2 (.DIODE(_04044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18315__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18316__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18317__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18318__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18320__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18321__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18323__A (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18324__A (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18324__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18324__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18325__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18326__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18327__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18328__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18329__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18330__A (.DIODE(_03317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18331__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18333__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18334__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18338__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18339__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18340__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18341__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18342__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18343__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18344__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18346__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18346__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__18346__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18347__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18348__A (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18349__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18351__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18351__B (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18351__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18352__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18353__A (.DIODE(_08775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18354__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18356__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18358__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18358__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18358__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18359__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18361__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__18364__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18367__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18370__A2 (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18372__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18373__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18374__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18375__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18376__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18376__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__18376__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18377__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18378__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18379__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18380__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18381__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18382__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18382__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__18382__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18383__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18384__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18385__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18386__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18386__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__18386__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18387__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18388__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18389__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18391__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18393__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18393__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18393__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18394__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18396__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__18402__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18405__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18408__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18411__A2 (.DIODE(_09287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18413__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18414__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18415__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18416__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18417__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18418__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18419__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18421__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18422__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18426__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18427__A1 (.DIODE(_04129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18428__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18430__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18432__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18433__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18434__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18436__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18438__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18438__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18438__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18439__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18440__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18440__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18440__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18441__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18442__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18443__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18445__A2 (.DIODE(_10591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18448__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__18450__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18451__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18452__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18454__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18455__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18457__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18458__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18459__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18460__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18461__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18462__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18463__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18464__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__A (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18467__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18468__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18469__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18471__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18471__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__18471__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18472__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18473__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18474__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18475__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18475__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__18475__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18476__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18477__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18478__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18479__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18480__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18482__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18482__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18482__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18483__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18485__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18487__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18488__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__18490__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18491__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__C (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18493__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18494__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18495__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18497__A (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18498__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18498__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18498__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18499__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18501__A2 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18502__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18503__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18504__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18505__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18508__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18510__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18513__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18514__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18516__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18517__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18519__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18520__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18522__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18523__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18525__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18526__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18528__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18529__A2 (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18531__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18532__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18534__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18535__A2 (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18537__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18539__A2 (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18542__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18545__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18548__A2 (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18551__A2 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18555__A2 (.DIODE(_09338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18558__A2 (.DIODE(_10202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18561__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18564__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__18567__A2 (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18570__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18573__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18576__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__A2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18582__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18585__A2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18587__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18589__A2 (.DIODE(_09494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18592__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18595__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18598__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18601__A2 (.DIODE(_09287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18603__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18604__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18605__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18606__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18607__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18608__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18610__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18611__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18614__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18614__B (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__A3 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18620__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18620__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18620__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18626__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18626__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18626__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18628__A (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18629__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18629__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18629__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18630__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18630__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18631__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18631__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18631__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18632__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18632__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18633__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18633__B (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18634__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18634__A3 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18636__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18636__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18638__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18638__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__18638__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18641__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18641__A2 (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18641__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18644__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18644__A2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18644__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18647__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18647__A2 (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18647__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18650__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18650__A2 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18650__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18652__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18652__B (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18653__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18653__A3 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18654__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18654__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__18654__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18655__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18655__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18656__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18656__B (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18657__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18657__A3 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18659__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18659__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18659__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18662__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18662__A2 (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18662__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18665__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18665__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18665__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18667__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18668__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18669__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18669__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18669__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18671__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18672__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18672__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18674__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18675__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18675__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__18677__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18677__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18677__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18678__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18678__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18679__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18680__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18680__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18682__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18682__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18682__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18683__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18683__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18684__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18684__B (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18685__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18685__A3 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18686__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18686__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18686__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18687__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18687__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18688__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18689__A1 (.DIODE(_04357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18689__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18691__A (.DIODE(_04350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18691__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18691__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18692__A1 (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18692__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18693__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__A2_N (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__B1 (.DIODE(_09294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18695__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__A2_N (.DIODE(_04354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__B1 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18697__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18698__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18698__A3 (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18701__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18702__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18706__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18707__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18708__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18709__A1 (.DIODE(_04235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18710__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18711__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18712__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18714__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18715__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18716__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18717__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18719__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18719__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18719__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18720__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18721__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18722__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18723__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18723__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18723__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18724__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18725__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18726__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18727__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18728__A2 (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18730__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18731__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__18733__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18734__A2 (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18736__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18737__A2 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18739__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18740__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18742__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18743__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18744__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18745__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__A2 (.DIODE(_09414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18750__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18751__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18752__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18752__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__18752__C (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18753__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18754__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18755__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18756__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18757__A2 (.DIODE(_09262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18759__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18760__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18762__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18763__A2 (.DIODE(_09268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18765__A (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18767__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18768__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18771__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18771__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18771__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18772__A2 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18773__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18774__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18776__A (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18777__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18777__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18777__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18778__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18779__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18780__B1 (.DIODE(_09293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18781__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18782__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18783__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18784__B1 (.DIODE(_11316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18786__A (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18787__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18789__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18792__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18794__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18797__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18798__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18799__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18800__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18802__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18805__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18808__A2 (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18811__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18814__A2 (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18816__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18817__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18819__A2 (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18822__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__18824__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18825__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18827__A2 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18830__A2 (.DIODE(_09337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18832__A (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18832__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__18832__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18833__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18835__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18837__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18838__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18840__A2 (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18843__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18845__A (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18845__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__18845__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18846__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18848__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18851__A2 (.DIODE(_09262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18854__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18856__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18857__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18858__A2 (.DIODE(_09268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18860__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18861__A2 (.DIODE(_09494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18863__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18864__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18865__A (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18865__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18865__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18866__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18867__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18868__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18870__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18871__A2 (.DIODE(_09287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__A (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18874__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18875__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18876__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18877__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18878__B1 (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18880__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18881__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18885__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18886__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18886__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18887__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18888__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18889__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18891__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18892__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18892__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18893__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18894__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18896__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18900__A1 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18900__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18901__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18902__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18902__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18903__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18903__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18903__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18904__A1 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18904__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18905__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18906__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18907__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__18911__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18912__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__18914__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18915__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18916__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18917__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18918__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18919__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18920__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18921__A2 (.DIODE(_09238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18923__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18924__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18926__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18927__A3 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18928__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18929__A2 (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18931__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18933__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18934__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18936__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18938__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18939__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__18941__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18941__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18941__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18942__A1 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18942__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18943__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18944__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18946__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18946__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18946__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18947__A1 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18947__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18948__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18950__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18950__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18950__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18951__A1 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18951__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18952__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18953__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18955__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18955__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18955__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18956__A1 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18956__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18957__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18957__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18957__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18958__A1 (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18958__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18959__A (.DIODE(_04221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18960__A2_N (.DIODE(_04528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18960__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18961__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18964__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18965__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18969__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18971__A (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18973__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18975__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18976__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18977__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18978__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18980__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18980__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18980__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18981__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18982__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18982__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18982__C (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18983__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18984__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18986__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18987__A2 (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18989__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18990__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__18992__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18993__A2 (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18995__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18996__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__18998__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18999__A2 (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19001__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19005__A (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19006__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19006__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19006__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19007__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19008__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19009__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19011__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19014__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19015__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19016__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19017__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19018__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19019__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19021__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19022__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19023__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19024__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__19026__A (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19027__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19027__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__19027__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19028__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19029__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19030__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19033__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19034__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19035__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19037__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19038__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19040__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19041__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__19043__A (.DIODE(_04576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19043__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19043__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19044__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19045__A (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19046__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19047__B1 (.DIODE(_09293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19048__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19049__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19050__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19051__B1 (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19053__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19054__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19058__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19059__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19059__A3 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19060__A (.DIODE(_09184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19061__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19061__A3 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19062__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19063__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19063__A3 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19064__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19064__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__19064__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19065__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19065__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19066__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19067__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19068__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19070__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19070__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19070__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19071__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19071__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19072__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19073__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19075__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19075__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19075__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19076__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19076__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19077__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19078__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19078__A3 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19079__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19080__A2 (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19082__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19083__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19084__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19086__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19087__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19088__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19089__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19090__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19091__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19093__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19093__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19094__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19095__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19097__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19098__A2 (.DIODE(_09414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19100__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19100__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__19100__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19101__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19101__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19102__A (.DIODE(_03482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19103__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19104__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19104__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__19104__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19105__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19105__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19106__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19108__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19109__A2 (.DIODE(_09262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19112__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19114__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19115__A2 (.DIODE(_09268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19118__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19118__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19119__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19120__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19121__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19121__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19121__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19122__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19122__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19124__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__19126__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19126__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19126__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19127__A1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19127__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19128__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19129__A2_N (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19129__B1 (.DIODE(_09293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19130__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19131__A2_N (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19131__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19132__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19133__A2_N (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19133__B1 (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19135__A (.DIODE(_04683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19136__A (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19139__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19140__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19141__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19144__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19145__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19147__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19148__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19150__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19151__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19153__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19154__A2 (.DIODE(_11330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19156__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19157__A2 (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19159__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19160__A2 (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19162__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19163__A2 (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19165__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19166__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19167__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19168__A2 (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__A (.DIODE(_04653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19171__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19173__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19174__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19175__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19176__A1 (.DIODE(_04610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19177__A (.DIODE(_09164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19179__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19180__A (.DIODE(_04683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19180__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19180__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19181__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19182__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19183__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19184__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19185__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19186__A (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19188__A2 (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19190__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19191__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19193__A (.DIODE(_04683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19193__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__19193__C (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19194__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19195__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19196__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19199__A2 (.DIODE(_09262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19201__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19202__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19204__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19205__A2 (.DIODE(_09268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19207__A (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19208__A (.DIODE(_04683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19208__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__19208__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19209__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19210__A (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19211__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19212__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19213__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19215__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19216__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__19218__A (.DIODE(_04683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19218__B (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19218__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19219__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19220__A (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__A (.DIODE(_04683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19222__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19223__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19224__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19225__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19226__B1 (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19229__A (.DIODE(_09190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19230__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19233__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19234__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19234__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19234__B1 (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__A (.DIODE(_09184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19238__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19238__A3 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19239__A (.DIODE(_09187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19239__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19240__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19240__A3 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19241__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19241__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__19241__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19242__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19242__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19243__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19243__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19243__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19244__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19244__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19245__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19245__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19245__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19246__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19246__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19247__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19248__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19248__B1 (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19250__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19250__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19250__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19251__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19251__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19252__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19252__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19253__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19253__A3 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19254__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19255__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19255__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__19255__B1 (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19258__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19258__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19260__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19260__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__A3 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19262__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19263__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19263__A2 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19265__A (.DIODE(_09235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19265__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19266__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19266__A3 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19267__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19268__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19268__A2 (.DIODE(_09238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19270__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19270__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19271__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19271__A3 (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19272__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19272__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19273__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19273__A3 (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19274__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19274__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__19274__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19275__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19275__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19276__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19277__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19277__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19279__A (.DIODE(_04718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19280__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19280__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19282__A (.DIODE(_09259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19282__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19283__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19283__A3 (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19284__A (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19286__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19286__A2 (.DIODE(_09262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19288__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19288__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__19288__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19289__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19289__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19291__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19291__A2 (.DIODE(_09268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19293__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19293__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__19293__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19294__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19294__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19296__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19296__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19298__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19298__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19298__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19299__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19299__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19301__A1 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19301__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__19303__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19303__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19303__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19304__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19304__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19305__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19305__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19305__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19306__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19306__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19307__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19308__A2_N (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19308__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19309__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19309__B (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19310__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19310__A3 (.DIODE(_04749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19312__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19313__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19317__A (.DIODE(_09180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19317__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19318__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19319__A (.DIODE(_09184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19319__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19320__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19321__A (.DIODE(_09187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19321__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19322__A1 (.DIODE(_04713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19324__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19325__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19325__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19325__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19326__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19327__A (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19329__A2 (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19329__B1 (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19331__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19331__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19332__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19334__A2 (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19334__B1 (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19336__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19336__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19339__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__19339__B1 (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19342__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19342__B1 (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19345__A2 (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19345__B1 (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19347__A (.DIODE(_09232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19347__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19348__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__A2 (.DIODE(_09337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__B1 (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19352__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19352__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19352__C (.DIODE(_04732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19353__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19355__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19358__A2 (.DIODE(_09414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19360__A (.DIODE(_09226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19361__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19361__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__19361__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19362__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19363__A (.DIODE(_09252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19363__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19364__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19366__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19369__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19372__A2 (.DIODE(_09262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19374__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19374__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__19374__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19375__A2 (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19377__A2 (.DIODE(_09268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19379__A (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19380__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19381__A2 (.DIODE(_09494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19383__A (.DIODE(_09276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19383__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19384__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19385__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19385__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19385__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19386__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19387__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19388__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__19390__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19391__A2 (.DIODE(_09287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19393__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19394__B1 (.DIODE(_09293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19395__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19396__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19397__A (.DIODE(_09299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19397__B (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19398__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19398__A3 (.DIODE(_04801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19401__A (.DIODE(_08794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19403__A (.DIODE(_09166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19406__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19407__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19407__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19407__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19409__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19410__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19410__A2 (.DIODE(_09314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19410__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19412__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__A2 (.DIODE(_09459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19415__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__A2 (.DIODE(_10983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19418__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19419__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19419__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19421__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19422__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19422__A2 (.DIODE(_09204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19422__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19424__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19425__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19425__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19427__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19428__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19428__A2 (.DIODE(_09211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19428__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19430__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19431__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19431__A2 (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19431__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19433__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19436__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19439__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__A2 (.DIODE(_09588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19442__A (.DIODE(_04840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__A2 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__B1 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19446__A (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19448__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19448__A2 (.DIODE(_09337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19451__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19451__A2 (.DIODE(_09238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19454__A1 (.DIODE(_04855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19454__A2 (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19457__A2 (.DIODE(_09414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19460__A2 (.DIODE(_09248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19463__A2 (.DIODE(_09347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19466__A2 (.DIODE(_09255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19469__A2 (.DIODE(_11136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19472__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__19475__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19478__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__19481__A2 (.DIODE(_09494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19484__A2 (.DIODE(_09365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19490__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__A2 (.DIODE(_09287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19496__A2_N (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19496__B1 (.DIODE(_09293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19497__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19498__A2_N (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19498__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19499__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19500__A2_N (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19500__B1 (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19502__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19503__A (.DIODE(_08795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19504__A (.DIODE(_09625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19508__A2 (.DIODE(_10239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19511__A (.DIODE(_09184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19512__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19512__A3 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19513__A (.DIODE(_09187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__A3 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19515__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19515__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__19515__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19516__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19516__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19517__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19517__B (.DIODE(_10586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19517__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19518__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19518__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19519__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19519__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19519__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19520__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19520__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19521__A (.DIODE(_09208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19522__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19523__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19523__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19523__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19524__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19524__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19525__A (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19526__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19527__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19528__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__19530__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19531__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__A (.DIODE(_09229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19534__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19535__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__A2 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19538__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19539__A2 (.DIODE(_09337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19541__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19541__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19541__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19542__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19542__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19543__A (.DIODE(_09242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19544__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19545__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19546__A2 (.DIODE(_09414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19548__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19548__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__19548__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19549__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19549__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19550__A (.DIODE(_09252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19551__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19552__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19552__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__19552__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19553__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19553__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19554__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19555__A2 (.DIODE(_09353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19557__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19558__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__19560__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19561__A2 (.DIODE(_09424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19563__A (.DIODE(_08777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19564__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__19566__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19566__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__19566__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19567__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19567__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19568__A (.DIODE(_09276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19569__A1 (.DIODE(_09224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19571__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19571__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19572__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19572__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__19572__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19574__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19574__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19574__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19575__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19575__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19576__A (.DIODE(_04922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19576__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19576__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19577__A1 (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19577__A2 (.DIODE(_08801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19578__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19579__A2_N (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19579__B1 (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19580__A (.DIODE(_04629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19581__A2_N (.DIODE(_04930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19581__B1 (.DIODE(_09441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19583__B (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19588__C (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19592__C (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19596__B (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19600__A (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19605__B (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19611__A (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19615__B (.DIODE(_09165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19619__B1 (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19623__A (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19625__A (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19626__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19627__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19629__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19630__A (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19640__A (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19641__A (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19642__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19648__A (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19648__B (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19652__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19655__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19657__A (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19659__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__C (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__B (.DIODE(_05045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__C (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19667__A (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19667__B (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19673__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19673__B (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19673__C (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19675__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19675__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19675__C (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19678__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19680__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19682__A (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19684__A (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19684__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19689__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19689__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19689__C (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__B (.DIODE(_05071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__C (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19696__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19696__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19696__C (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19699__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19699__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19699__C (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19704__A (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19706__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19706__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19708__A (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19709__A (.DIODE(_05088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19711__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19712__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19712__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19712__C (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19714__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19716__A (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19718__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19718__B (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19718__C (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19719__A (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19720__A (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19721__A (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19722__A (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19724__B (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19724__D (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19725__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19725__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19725__C (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19727__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19727__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19727__C (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19729__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19730__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19730__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19732__A (.DIODE(_05111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19733__A (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19734__B (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19738__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19738__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19738__C (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19740__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19740__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19740__C (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19742__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19742__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19742__C (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19744__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19744__A2 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19746__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19746__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19746__C (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19748__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19748__B (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19748__C (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19751__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19751__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19751__C (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19755__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19755__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19755__C (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19762__A (.DIODE(_05141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19763__A (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19763__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19763__C (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19765__A (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19767__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19769__A (.DIODE(_05148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19769__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19771__A (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19772__A (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19772__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19773__A_N (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19773__B (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19773__C (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19777__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19781__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19782__B (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19782__C (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19782__D (.DIODE(_05161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19784__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19784__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19786__A (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19786__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19788__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19791__A (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19791__C (.DIODE(_05168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19791__D (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19792__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19794__A (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19794__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19795__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19797__A (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19797__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19799__A (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19799__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19801__A (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19801__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19802__A (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19802__B (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19805__A (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19806__A (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19807__A (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19808__A (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19810__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19811__A (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19812__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19815__A (.DIODE(_05141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19816__B (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19817__A1 (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19817__A2 (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19817__B1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19818__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19818__B (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19819__A (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19820__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19821__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19823__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19824__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19826__A (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19827__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19828__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19829__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19829__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19830__A1 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19830__A2 (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19830__A3 (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19831__A (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19831__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19832__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19832__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19833__A (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19833__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19834__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19834__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19835__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19835__B (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19837__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19837__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19838__B (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19840__A (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19841__D (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19843__A (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19843__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19844__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19844__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19845__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19845__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19846__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19846__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19847__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19848__A (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19849__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19849__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19850__A1 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19850__A2 (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19850__A3 (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19851__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__A (.DIODE(_05231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19854__A (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19854__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19855__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19855__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19856__A1 (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19856__A2 (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19856__A3 (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19857__A1 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19857__A2 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19857__A3 (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19857__B1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19859__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19859__A2 (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19861__A (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19861__B (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19862__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19863__A (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19863__B (.DIODE(_05141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__A (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__B (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__A (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__B (.DIODE(_05088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19867__A1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19867__A2 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19867__A3 (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19867__A4 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19867__B1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19869__A (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19869__B (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19870__A (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19871__A (.DIODE(_05141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19871__B (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19873__A (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19873__B (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19874__A (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19874__B (.DIODE(_05088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19876__A1 (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19876__A2 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19876__A3 (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19876__A4 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19876__B1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19877__A (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19878__A (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19879__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19879__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19879__C (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19881__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19881__B (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19881__C (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19882__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19882__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19882__C (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19883__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19883__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19883__C (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19884__B (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19884__C (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19884__D (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19885__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19885__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19885__C (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19887__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19887__B (.DIODE(_05045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19887__C (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__C (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19891__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19891__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19891__C (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19893__A (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19893__C (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__C (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19896__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19896__B (.DIODE(_05071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19896__C (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19898__A (.DIODE(_05005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19898__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19898__C (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19900__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19900__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19900__C (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19902__B (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19902__C (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19902__D (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19903__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19903__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19903__C (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19904__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19905__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19905__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__A (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__B (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__C (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19908__A (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19908__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19909__A (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19909__B (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19909__C (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19911__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19911__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19911__C (.DIODE(_05054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19913__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19913__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19913__C (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19915__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19915__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19917__A1 (.DIODE(_05111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19917__A2 (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19917__D1 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19918__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19918__B (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19918__C (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19919__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19919__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19919__C (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19921__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19921__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19921__C (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19922__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19922__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19922__C (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__A (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__B (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__C (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__D (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19924__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19924__B (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19924__C (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19925__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19925__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19925__C (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19927__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19927__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19927__C (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19928__A (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19928__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19930__A (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19930__B (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19930__C (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19930__D (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19931__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19931__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19931__C (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19933__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19933__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19933__C (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19935__A (.DIODE(_05091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19935__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19935__C (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19936__A (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19936__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19938__B (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19938__C (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19941__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19941__A2 (.DIODE(_05148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19941__A3 (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19941__A4 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19941__B1 (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19942__A (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19942__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19943__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19944__A (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19944__B (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19945__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19946__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19947__A (.DIODE(_05325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19947__B (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19948__A1 (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19948__A2 (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19948__B1 (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19949__A (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19949__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19949__C (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19950__A (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19950__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19950__C (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__A (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__B (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19953__A (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19953__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19954__A (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19954__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19955__A (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19955__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19956__A (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19956__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19959__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19959__A2 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19959__A3 (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19959__B1 (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19959__C1 (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19960__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19962__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19962__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19962__C (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19965__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19967__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19967__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19967__C (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19969__A1 (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19969__C1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19970__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19970__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19970__C (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__C (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19974__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19974__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19974__C (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19977__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19977__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19979__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19979__B (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19979__C (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19979__D (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19981__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19982__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19983__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19985__A (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19985__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19987__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19988__C (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19992__A (.DIODE(_05371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19994__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19994__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19995__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19995__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19996__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19996__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19997__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19997__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20000__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20000__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20001__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20002__A (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20002__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20002__C (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20003__A (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20003__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20004__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20004__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20005__A (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20005__B (.DIODE(_08677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20006__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20006__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20008__B2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20009__A (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20009__B (.DIODE(_05099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20010__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20010__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20011__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20011__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20012__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20012__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20013__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20013__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20014__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20016__A (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20016__B (.DIODE(_08678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20017__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20017__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20018__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20018__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20019__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20019__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20021__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20021__B (.DIODE(\line_cache[154][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20022__B1 (.DIODE(_05401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20027__A (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20029__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20030__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20031__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20032__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20032__C (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20034__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20034__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20036__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20036__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20037__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20037__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20038__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20038__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20039__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20039__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20043__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20043__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20044__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20044__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20047__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20047__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20051__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20051__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20052__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20052__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20053__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20053__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20054__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20054__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20058__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20058__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20059__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20059__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20060__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20060__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20062__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20065__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20065__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20066__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20066__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20067__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20067__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20069__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20069__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20073__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20073__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20074__A (.DIODE(_08676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20075__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20076__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20076__B (.DIODE(_05455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20077__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20077__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20078__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20078__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20080__B2 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20081__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20081__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20082__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20082__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20083__A (.DIODE(_05249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20083__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20084__A (.DIODE(_05250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20084__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20087__D (.DIODE(_05466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20088__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20088__B (.DIODE(_05455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20089__A (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20090__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20091__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20092__A (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20093__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20094__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20095__A (.DIODE(_05231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20096__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20097__A1 (.DIODE(\line_cache[191][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20097__A2 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20098__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20098__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20099__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20099__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20104__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20104__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20107__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20107__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20109__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20109__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20111__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20111__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20112__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20112__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20113__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20113__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20115__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20115__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20120__B (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20121__B (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20122__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20122__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20123__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20123__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20124__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20124__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20126__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20126__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20129__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20129__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20130__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20130__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20131__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20131__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20134__A2 (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20135__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20135__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20136__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20136__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20139__B (.DIODE(_05185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20139__C (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20140__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20140__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20141__A1 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20142__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20142__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20143__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20143__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20144__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20144__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20149__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20149__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20150__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20150__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20151__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20151__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20152__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20152__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20155__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20155__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20156__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20157__A (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20157__B (.DIODE(_05100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20157__C (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20158__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20158__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20159__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20159__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20161__B2 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20162__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20162__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20163__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20163__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20164__A (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20165__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20165__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20166__A3 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20170__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20170__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20171__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20171__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20173__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20173__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20179__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20179__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20180__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20180__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20181__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20181__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20182__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20183__A (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20183__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20186__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20186__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20187__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20187__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20188__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20188__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20189__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20189__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20193__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20193__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20194__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20194__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20195__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20195__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20196__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20196__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20199__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20199__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20200__A (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20200__B (.DIODE(_05455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20201__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20201__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20202__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20202__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20205__A (.DIODE(_05565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20207__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20207__B (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20209__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20209__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20210__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20210__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20211__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20211__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20214__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20214__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20215__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20215__B (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20217__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20217__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20218__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20218__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20222__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20222__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20223__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20223__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20224__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20224__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20225__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20225__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20228__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20228__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20229__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20229__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20230__A (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20231__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20232__A (.DIODE(_05253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20232__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20233__A1 (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20233__A3 (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20237__A (.DIODE(_05437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20237__B (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20237__C (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20240__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20240__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20243__A (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20244__A (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20250__A (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20251__A (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20255__A2 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20255__B2 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20258__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20263__A (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20263__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20272__B1 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20273__C (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20274__A (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20275__A (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20276__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20276__A2 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20277__A2 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20278__A (.DIODE(_05168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20279__A (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20280__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20282__A (.DIODE(_05161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20287__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20288__A (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20289__B (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20290__A (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20291__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20291__A2 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20293__A (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20293__B (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20293__C (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20294__A (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20295__A (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20295__B (.DIODE(_05071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20295__C (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20296__A (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20297__A (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20298__A (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20302__C (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20303__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20303__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20304__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20304__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20305__A (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20306__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20306__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20307__A (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20307__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20310__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20310__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20311__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20311__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20312__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20312__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20313__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20315__A (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20315__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20318__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20318__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__A (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__C (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20320__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20320__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20321__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20321__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20324__A (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20325__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20325__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20327__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20328__A (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20329__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20330__A (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20331__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20334__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20334__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20335__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20335__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20336__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20336__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20337__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20337__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20340__A (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20340__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20340__C (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20342__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20342__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20343__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20343__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20344__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20344__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20346__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20346__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20347__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20347__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20348__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20348__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20349__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20349__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20353__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20353__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20354__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20354__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20355__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20355__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20356__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20356__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20359__A (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20360__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20360__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20361__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20361__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20362__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20362__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20363__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20364__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20364__B (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20365__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20365__B (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20366__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20366__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20367__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20367__B (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20370__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20370__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20373__A (.DIODE(_05199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20373__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20376__D (.DIODE(_05755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20377__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20377__C (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20380__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20380__C (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20381__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20381__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20382__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20382__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20382__C (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20384__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20384__C (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20385__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20386__A2 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20387__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20387__C (.DIODE(_05042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20389__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20390__A (.DIODE(_05769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20392__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20392__B (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20392__C (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20394__A1 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20394__A2 (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20396__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20396__C (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20400__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20400__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20401__A1 (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20401__A3 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20405__A (.DIODE(_05682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20405__B (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20406__B (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20410__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20412__A (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20413__A (.DIODE(_05111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20413__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20414__A (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20414__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__A (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__A1 (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__A2 (.DIODE(\line_cache[271][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20417__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20417__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20417__C (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20419__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20419__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20421__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20421__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20422__A1 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20422__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20425__A1 (.DIODE(\line_cache[255][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20425__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20426__A (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20427__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20427__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20430__A2 (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20431__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20432__A (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20433__A (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20433__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20434__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20434__A3 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20435__A (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20435__B (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20436__A (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20436__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20438__A (.DIODE(_05148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20438__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20440__A (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20440__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20441__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20441__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20445__A (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20446__A (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20447__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20447__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20448__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20448__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20451__A (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20452__A (.DIODE(_05325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20453__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20453__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20456__A1 (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20456__B2 (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20457__A2 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20457__B2 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20460__A (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20461__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20461__A2 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20461__B1 (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20465__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20465__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20466__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20466__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20467__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20467__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20468__A2 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20468__B2 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20470__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20470__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20471__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20471__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20472__A (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20473__A2 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20474__A2 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20474__B2 (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20478__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20478__B (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20479__B1 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20480__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20480__B (.DIODE(_05383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20481__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20481__B (.DIODE(_05385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20485__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20485__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20486__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20486__B (.DIODE(_05208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20487__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20487__B (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20488__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20488__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20491__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20491__B (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20492__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20492__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20493__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20493__B (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20495__A (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20495__B (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20499__A (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20500__B (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20501__A (.DIODE(_05617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20501__B (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20502__A (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20504__A (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20507__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20507__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20508__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20508__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20515__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20516__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20517__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20518__A1 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20521__B1 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20522__A1 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20522__A2 (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20523__B2 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20531__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20534__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20534__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20535__A (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20535__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20536__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20536__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20538__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20538__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20539__A1 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20539__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20540__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20540__A3 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20547__A2 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20547__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20548__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20548__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20555__B (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20556__A (.DIODE(_05909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20557__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20557__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20558__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20558__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20559__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20559__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20560__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20574__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20574__C (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20576__A3 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20577__A2 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20578__D1 (.DIODE(_05956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20580__B (.DIODE(_05958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20583__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20583__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20584__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20584__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20585__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20585__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20587__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20587__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20588__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20588__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20589__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20589__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20590__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20590__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20599__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20600__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20601__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20602__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__A (.DIODE(_05195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20608__B (.DIODE(_05986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20612__A (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20613__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20613__B (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20615__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20615__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20616__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20616__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20618__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20620__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20620__A2 (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20621__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20623__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20625__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20625__B1 (.DIODE(\line_cache[287][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20626__D_N (.DIODE(_06004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20627__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20627__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20628__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20628__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20629__A (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20630__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20632__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20632__B2 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20637__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20637__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20638__A2 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20645__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20645__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20646__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20646__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20647__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20647__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20648__A1 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20648__B1 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20650__C (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20650__D (.DIODE(_06028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20651__A (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20652__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20655__A (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20656__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20658__A1 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20658__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20660__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20660__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20661__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20661__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20663__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20663__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20666__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20666__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20667__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20667__B2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20668__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20668__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__A3 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20671__A1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20671__A2 (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__A2 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20675__A (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20679__B (.DIODE(_06049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20680__B (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20681__C (.DIODE(_06059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20682__A (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20688__A2 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20696__A (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20703__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20703__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20706__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20706__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20709__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20709__B (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20714__B (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20715__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20715__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20719__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20723__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20723__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20728__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20728__B (.DIODE(_05201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20731__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20740__A1 (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20749__B1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20751__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20760__A2 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20763__C (.DIODE(_06141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20764__A (.DIODE(_05989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20764__B (.DIODE(_06060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20764__C (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20768__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20768__B (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20770__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20770__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20771__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20771__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20773__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20774__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20774__A2 (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20775__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20777__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20779__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20781__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20781__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20782__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20782__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20783__A (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20784__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20786__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20786__B2 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20791__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20791__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20792__A2 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20799__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20799__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20800__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20800__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20801__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20801__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20802__A1 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20802__B1 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20804__A (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20804__C (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20804__D (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20805__A (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20806__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20809__A (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20810__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20812__A1 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20812__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20814__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20814__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20815__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20815__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20817__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20817__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20820__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20820__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20821__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20821__B2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20822__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20822__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20823__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20823__A3 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20825__A1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20825__A2 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20826__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20826__A2 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20828__A (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20832__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20833__B (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20834__C (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20835__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20838__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20838__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20839__A (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20839__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20840__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20840__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20842__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20842__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20843__A1 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20843__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20844__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20844__A3 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20851__A2 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20851__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20852__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20852__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20860__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20860__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20861__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20861__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20868__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20868__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20869__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20869__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20870__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20871__A1 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20878__B1 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20880__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20881__A1 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20881__A2 (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20884__B (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20887__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20887__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20888__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20888__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20889__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20889__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20891__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20892__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20893__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20894__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20894__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20903__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20903__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20904__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20904__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20905__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20905__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20906__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20910__C (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20911__B (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20912__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20912__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20913__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20913__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20914__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20914__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20915__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20931__C (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20933__A2 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20934__D (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20936__B (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20936__D (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20938__B1 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20940__A (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20947__C (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20954__A (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20958__D (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20963__A1 (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20968__A2 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20973__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20987__B1 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20992__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20992__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20996__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21000__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21000__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21004__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21004__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21015__B (.DIODE(_06369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21016__A (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21016__B (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21016__C (.DIODE(_06393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21019__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21019__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21020__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21020__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21027__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21028__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21029__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21030__A1 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21033__B1 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21034__A1 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21034__A2 (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21035__B2 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21043__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21046__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21046__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21047__A (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21047__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21048__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21048__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21050__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21050__B (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21051__A1 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21051__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21052__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21052__A3 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21059__A2 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21059__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21060__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21060__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21068__A (.DIODE(_06419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21069__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21069__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21070__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21070__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21071__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21071__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21072__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21086__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21086__C (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21088__A3 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21089__A2 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21092__B (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21095__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21095__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21096__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21096__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21097__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21097__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21099__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21099__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21100__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21100__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21101__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21101__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21102__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21102__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21111__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21112__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21113__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21114__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21119__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21123__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21123__B (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21125__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21125__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21126__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21126__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21128__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21129__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21129__A2 (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21130__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21132__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21134__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21135__D_N (.DIODE(_06511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21136__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21136__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21137__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21137__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21138__A (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21139__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21141__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21141__B2 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21146__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21146__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21147__A2 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21154__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21154__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21156__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21156__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21157__A1 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21157__B1 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21159__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21159__D (.DIODE(_06535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21160__A (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21161__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21164__A (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21165__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21167__A1 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21167__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21169__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21169__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21170__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21170__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21172__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21172__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21175__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21175__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21176__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21176__B2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21177__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21177__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21178__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21178__A3 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21180__A1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21180__A2 (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21181__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21181__A2 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21183__A (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21187__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21188__B (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21189__C (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21195__B2 (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21203__A2 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21212__B1 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21221__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21227__B (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21230__A1 (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21239__B1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21242__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21242__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21251__A (.DIODE(_06621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21253__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21257__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21257__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21264__A (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21264__B (.DIODE(_06618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21265__A (.DIODE(_06498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21265__B (.DIODE(_06566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21265__C (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21269__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21269__B (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21271__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21271__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21272__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21272__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21274__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21275__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21275__A2 (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21276__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21278__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21280__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21281__D_N (.DIODE(_06656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21282__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21282__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21283__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21283__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21284__A (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21285__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21287__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21287__B2 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21292__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21292__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21293__A2 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21300__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21300__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21301__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21301__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21302__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21302__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21303__A1 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21303__B1 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21305__A (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21305__D (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21306__A (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21307__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21310__A (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21311__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21313__A1 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21313__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21315__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21315__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21316__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21316__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21318__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21318__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21321__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21321__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21322__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21322__B2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21323__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21323__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21324__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21324__A3 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21326__A1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21326__A2 (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21327__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21327__A2 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21329__A (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21334__B (.DIODE(_06696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21336__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21336__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21337__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21337__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21344__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21344__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21345__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21346__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21347__A1 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21350__B1 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21351__A1 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21351__A2 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21352__B2 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21362__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21362__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21363__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21363__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21364__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21364__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21366__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21367__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21368__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21369__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21369__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21378__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21378__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21379__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21379__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21380__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21380__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21381__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21386__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21387__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21387__C (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21388__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21388__C (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21389__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21398__B1 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21399__A3 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21409__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21410__B (.DIODE(_06761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21411__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21414__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21414__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21415__A (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21415__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21416__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21416__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21418__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21418__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21419__A1 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21419__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21420__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21420__A3 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21427__A2 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21427__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21428__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21428__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21439__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21442__A2 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21444__A1 (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21449__B1 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21458__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21470__A (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21476__B (.DIODE(_06845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21480__A2 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21487__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21487__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21490__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21490__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21497__B (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21499__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21503__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21503__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21510__A (.DIODE(_06841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21510__B (.DIODE(_06862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21511__A (.DIODE(_06711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21511__B (.DIODE(_06812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21511__C (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21515__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21515__B (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21517__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21517__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21518__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21518__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21520__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21521__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21521__A2 (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21522__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21524__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21526__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21527__D_N (.DIODE(_06901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21528__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21528__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21529__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21529__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21530__A (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21531__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21533__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21533__B2 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21538__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21538__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21539__A2 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21546__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21546__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21547__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21547__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21548__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21548__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21549__A1 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21549__B1 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21552__A (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21553__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21556__A (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21557__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21559__A1 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21559__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21561__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21561__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21562__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21562__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21564__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21564__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21567__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21567__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21568__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21568__B2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21569__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21569__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21570__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21570__A3 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21572__A1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21572__A2 (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21573__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21573__A2 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21575__A (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21582__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21582__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21583__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21583__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21590__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21590__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21591__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21592__A (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21593__A1 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21596__B1 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21597__A1 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21597__A2 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21598__B2 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21608__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21608__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21609__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21609__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21610__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21610__C (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21612__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21613__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21614__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21615__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21615__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21624__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21625__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21625__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21626__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21626__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21627__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21632__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21633__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21633__C (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21634__C (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21635__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21644__B1 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21645__A3 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21654__A (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21655__B (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21656__B (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21657__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21660__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21660__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21661__A (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21661__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21662__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21662__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21664__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21664__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21665__A1 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21665__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21666__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21666__A3 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21673__A2 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21673__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21674__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21674__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21680__A (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21681__B (.DIODE(_07055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21683__A (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21689__A2 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21697__A (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21704__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21704__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21708__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21712__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21712__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21716__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21716__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21729__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21743__A2 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21745__A1 (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21754__B1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21756__C (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21758__A (.DIODE(_06956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21758__B (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21758__C (.DIODE(_07132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21762__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21762__B (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21764__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21764__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21765__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21765__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21767__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21768__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21768__A2 (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21769__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21771__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21771__B (.DIODE(\line_cache[271][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21773__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21773__B1 (.DIODE(\line_cache[287][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21774__D_N (.DIODE(_07147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21775__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21775__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21776__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21776__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21777__A (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21778__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21780__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21780__B2 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21785__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21785__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21786__A2 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21793__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21793__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21794__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21794__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21795__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21795__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21796__A1 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21796__B1 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21799__A (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21800__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21803__A (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21804__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21806__A1 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21806__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21808__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21808__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21809__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21809__B (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21811__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21811__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21814__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21814__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21815__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21815__B2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21816__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21816__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21817__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21817__A3 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21819__A1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21819__A2 (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21820__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21820__A2 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21822__A (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21829__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21832__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21832__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21833__A (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21833__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21834__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21834__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21836__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21836__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21837__A1 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21837__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21838__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21838__A3 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21845__A2 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21845__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21846__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21846__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21854__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21854__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21855__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21855__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21862__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21862__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21863__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21863__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21864__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21865__A1 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21872__B1 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21874__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21875__A1 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21875__A2 (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21878__B (.DIODE(_07251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21881__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21881__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21882__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21882__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21883__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21883__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21885__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21886__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21887__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21888__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21888__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21897__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21897__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21898__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21898__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21899__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21899__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21900__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21905__B (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21906__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21906__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21907__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21907__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21908__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21908__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21909__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21925__C (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21927__A2 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21929__B (.DIODE(_07302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21930__B (.DIODE(_07252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21931__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21939__A2 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21946__B2 (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21951__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21951__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21962__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21969__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21969__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21976__A1 (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21981__A2 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21990__A2 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21995__A (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22005__A (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22005__C (.DIODE(_07378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22006__A (.DIODE(_07202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22006__B (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22006__C (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22012__A2 (.DIODE(_05519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22023__B2 (.DIODE(_05502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22028__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22028__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22031__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22031__C (.DIODE(_05562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22039__A (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22039__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22043__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22048__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22048__C (.DIODE(_05381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22059__B1 (.DIODE(_05468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22066__A1 (.DIODE(_05392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22074__B1 (.DIODE(\line_cache[168][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22075__A1 (.DIODE(_05409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22084__B1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22086__A (.DIODE(_07426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22086__D (.DIODE(_07458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22088__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22088__B (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22090__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22090__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22091__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22091__A3 (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22093__B (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22094__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22094__A2 (.DIODE(_05180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22095__A1 (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22097__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22097__B (.DIODE(\line_cache[271][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22099__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22099__B1 (.DIODE(\line_cache[287][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22100__D_N (.DIODE(_07472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22101__A1 (.DIODE(_05283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22101__B2 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22102__A1 (.DIODE(_05298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22102__B2 (.DIODE(_05300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22103__A (.DIODE(_05279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22104__A (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22106__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22106__B2 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22111__A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22111__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22112__A2 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22119__A1 (.DIODE(_05314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22119__B2 (.DIODE(_05315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22120__A1 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22120__B2 (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22121__A1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22121__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22122__A1 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22122__B1 (.DIODE(_05309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22125__A (.DIODE(_05365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22126__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22129__A (.DIODE(_05353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22130__A (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22132__A1 (.DIODE(_05355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22132__B1 (.DIODE(_05346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22134__A (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22134__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22135__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22135__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22137__A1 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22137__B2 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22140__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22140__B2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22141__A2 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22141__B2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22142__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22142__B (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22143__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22143__A3 (.DIODE(_05320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22145__A1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22145__A2 (.DIODE(_05812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22146__A1 (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22146__A2 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22148__A (.DIODE(_05270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22154__C (.DIODE(_07526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22155__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22158__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22158__B (.DIODE(_05021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22159__A (.DIODE(_05771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22159__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22160__A (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22160__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22162__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22162__B (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22163__A1 (.DIODE(_05760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22163__B2 (.DIODE(_05764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22164__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22164__A3 (.DIODE(_05364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22171__A2 (.DIODE(_05097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22171__B2 (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22172__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22172__B2 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22180__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22180__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22181__A (.DIODE(_05586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22181__C (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22188__A (.DIODE(_05470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22188__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22189__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22189__C (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22190__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22191__A1 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22198__B1 (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22200__A1 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22201__A1 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22201__A2 (.DIODE(_05151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22204__B (.DIODE(_07576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22207__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22207__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22208__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22208__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22209__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22209__C (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22211__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22212__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22213__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22214__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22214__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22223__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22224__A (.DIODE(_05610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22224__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22225__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22225__C (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22226__A (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22231__B (.DIODE(_07603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22232__A (.DIODE(_05454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22232__C (.DIODE(_05732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22233__A (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22233__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22234__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22234__C (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22235__A1 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22251__C (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22253__A2 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22255__B (.DIODE(_07627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22256__B (.DIODE(_07577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22257__A (.DIODE(_07459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22257__B (.DIODE(_07527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22259__A (.DIODE(net4215));
 sky130_fd_sc_hd__diode_2 ANTENNA__22259__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__22261__A (.DIODE(net4215));
 sky130_fd_sc_hd__diode_2 ANTENNA__22262__A (.DIODE(_08726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22262__B (.DIODE(_07632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22263__A2 (.DIODE(_07633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22263__B1 (.DIODE(_08771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22264__A (.DIODE(net2713));
 sky130_fd_sc_hd__diode_2 ANTENNA__22264__B (.DIODE(_09359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22266__A1 (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22269__A2 (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22272__B2 (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22276__B2 (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22279__B2 (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22282__B2 (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22283__A2 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22283__A3 (.DIODE(_10466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22284__A1_N (.DIODE(_10238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22284__B1 (.DIODE(_08728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22284__B2 (.DIODE(net2713));
 sky130_fd_sc_hd__diode_2 ANTENNA__22285__C (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22288__A (.DIODE(_08771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22300__B1 (.DIODE(_07632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22301__A (.DIODE(_09225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22301__B (.DIODE(_07633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22302__A (.DIODE(_07662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22302__B (.DIODE(_07663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22303__A (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22304__A (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22304__B (.DIODE(_08726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22306__A (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22307__A (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22308__A2 (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22311__A (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22312__A1 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22312__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22313__B (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22315__A (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22315__B (.DIODE(_09192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22316__A (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22318__B (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22320__B1 (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22322__A (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22323__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22325__A1 (.DIODE(_07662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22325__A2 (.DIODE(_07663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22326__A1 (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22326__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22327__A1 (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22329__B (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22330__B (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22335__A (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22337__B1 (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22340__B (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22341__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22344__A (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22348__B (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22349__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22352__A (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22356__C (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22357__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22360__A (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22361__B1 (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22363__B (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22364__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22367__A (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22371__B1 (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22371__C1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22378__A (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22379__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22379__A4 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22383__A2 (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22383__B2 (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22384__A (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22385__B1 (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22393__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22394__A3 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22394__A4 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22400__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22401__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22401__A4 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22405__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22406__A3 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22406__A4 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22412__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22413__A3 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22413__A4 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22417__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22418__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22418__A4 (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22424__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22425__A2 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22425__A4 (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22429__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22430__A3 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22430__A4 (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22434__B (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22435__A3 (.DIODE(_08791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22435__A4 (.DIODE(_07665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22439__A2 (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22439__B2 (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22441__B (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22442__A1 (.DIODE(_07664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22443__B (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22447__B1 (.DIODE(_07676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22448__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__22448__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__22449__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__22450__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__22452__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__22454__A (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22454__B (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22455__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22455__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22456__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22457__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__22458__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__22458__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__22459__A (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22460__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__22460__B1 (.DIODE(_07791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22461__B (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22463__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22465__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22465__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22466__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22467__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22470__B (.DIODE(_07791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22471__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22471__B2 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22472__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22474__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22474__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22475__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22476__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22479__B (.DIODE(_07791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22480__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22480__B2 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22481__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22483__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22483__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22484__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22485__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22487__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22487__B1 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22488__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22491__B (.DIODE(_07791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22492__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22494__A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__22494__S (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22496__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__22496__S (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22498__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__22498__S (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22500__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__22500__S (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22502__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__22502__S (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22504__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22505__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__22507__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__22509__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__22537__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22538__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22540__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22542__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22544__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22546__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22548__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22550__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22552__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22554__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22556__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22558__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22560__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22562__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22564__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22566__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22568__S (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22570__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22571__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22573__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22575__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22577__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22579__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22581__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22583__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22585__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22587__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22589__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22591__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22593__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__22593__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22593__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22593__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__22594__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__22594__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22595__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22597__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__22597__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22597__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22597__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__22598__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__22598__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22599__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22601__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__22601__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22601__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22601__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__22602__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__22602__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22603__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22605__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__22605__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22605__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22605__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__22606__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__22606__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22607__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22609__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__22609__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22609__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22609__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__22610__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__22610__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22611__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22613__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__22613__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22613__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22614__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__22614__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22615__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22617__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22617__B1 (.DIODE(_07785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22618__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__22618__A2 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22619__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22621__A2 (.DIODE(_07783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22621__B1 (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22622__S (.DIODE(_07794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22624__A (.DIODE(_07786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22736__B1 (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22738__B1 (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22739__C (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22750__C (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22759__C (.DIODE(\base_h_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22784__A (.DIODE(_08722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22784__B (.DIODE(net4316));
 sky130_fd_sc_hd__diode_2 ANTENNA__22785__B (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22787__A0 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22787__A1 (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22793__A2 (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22793__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22795__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22800__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22804__A2 (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22804__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22808__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22812__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22816__A2 (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22816__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22820__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22822__A2 (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22822__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22823__A (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22823__B (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22920__B (.DIODE(\base_v_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22921__C (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22939__B (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22940__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22947__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22953__A (.DIODE(_08722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22955__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22963__B (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22971__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22972__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22985__B (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22993__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22994__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23003__B1 (.DIODE(_03834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23009__A (.DIODE(_08722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23011__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23015__B (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23020__A (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23021__A (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23023__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23025__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23029__A1 (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23032__A (.DIODE(_08722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23034__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23038__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23044__A (.DIODE(_08722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23046__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23049__A (.DIODE(_09223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23056__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23057__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23059__B1 (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23064__B1 (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23066__A (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23067__A (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23072__B (.DIODE(_09222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23074__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23075__C (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23076__A (.DIODE(_08722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23078__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23083__C1 (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23088__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23089__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23093__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23094__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23097__B (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23100__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23104__A (.DIODE(_05061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23104__B (.DIODE(_05088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23105__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23106__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23111__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23112__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23116__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23117__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23120__B (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23121__B (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23122__B (.DIODE(_10310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23123__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23124__B (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23127__B1 (.DIODE(_08800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23128__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23132__A (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23172__B1 (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23173__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23173__B (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23174__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23181__B1 (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23182__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23184__B (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23185__A (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23186__A (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23188__A (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23193__B1 (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23194__B1 (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23195__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23200__A (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23201__B1 (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23202__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23206__B (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23208__B1 (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23209__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23213__B (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23214__A (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23216__A (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23219__B1 (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23220__A2 (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23221__C (.DIODE(_08051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23222__A2 (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23224__B (.DIODE(_08774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23227__A (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23232__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23233__C (.DIODE(_08460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23234__B (.DIODE(_08661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23237__B (.DIODE(_08464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23238__A (.DIODE(_08464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23241__A (.DIODE(_08793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23243__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23245__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23247__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23249__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23251__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__23251__S (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23253__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__23253__S (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23255__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__23255__S (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23257__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__23257__S (.DIODE(_09375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23259__B (.DIODE(_04971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23261__B (.DIODE(_08460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23267__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23273__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23276__B1 (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23278__A (.DIODE(_08318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23281__A (.DIODE(_08661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23281__B (.DIODE(_08776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23284__A1 (.DIODE(_08723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23303__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23304__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23305__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__23306__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__23307__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23308__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__23309__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23353__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23355__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23356__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23363__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23365__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23366__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23367__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23368__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23369__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23370__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23371__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23372__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23373__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23374__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23375__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23376__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23377__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23379__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23380__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23387__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23388__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23389__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23390__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23391__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23392__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23393__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23394__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23395__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23396__RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__23415__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23416__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23418__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23419__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23420__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23421__RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__23424__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23435__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23436__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23437__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23444__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23445__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23446__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23447__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23450__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23453__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23454__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__23521__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23535__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23549__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__23622__RESET_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__23627__RESET_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__23630__RESET_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__24018__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24019__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24026__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24027__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24030__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24032__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24033__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24036__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24039__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24040__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24041__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24044__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24047__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24064__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__24449__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__24455__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__24463__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__24467__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__24468__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__24475__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__24516__RESET_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__24517__RESET_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__24521__RESET_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__24522__RESET_B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__24550__RESET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__24555__RESET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__24589__RESET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__24981__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__24982__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__24998__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__25056__RESET_B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__25057__RESET_B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__25086__RESET_B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__25426__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__25434__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25436__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25438__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__25439__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25440__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25441__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__25442__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__25443__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25444__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25445__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25446__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25466__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25469__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25473__RESET_B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__25474__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__25678__CLK (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__25691__RESET_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__25692__RESET_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__25820__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__25822__RESET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__25829__RESET_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__25903__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25911__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25915__RESET_B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__25919__RESET_B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__25920__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25921__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25924__RESET_B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__25926__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25927__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25928__RESET_B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__25929__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25932__RESET_B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__25934__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25935__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25940__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__25944__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__25948__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__25951__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25956__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__25959__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__25964__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__25967__RESET_B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__26067__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_0__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_10__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_11__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_12__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_13__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_14__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_15__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_16__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_17__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_18__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_19__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_1__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_20__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_21__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_22__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_23__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_24__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_25__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_26__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_27__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_28__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_29__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_2__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_30__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_31__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_3__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_4__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_5__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_6__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_7__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_8__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_9__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_140_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_141_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_142_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_143_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_144_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_145_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_146_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_147_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_148_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_149_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_150_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_151_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_152_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_153_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_154_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_155_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_156_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_157_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_158_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_159_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_160_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_161_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_162_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_163_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_164_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_165_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_166_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_167_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_168_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_169_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_170_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_171_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_172_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_173_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_174_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_175_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_176_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_177_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_178_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_179_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_180_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_181_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_182_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_183_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_184_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_185_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_186_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_187_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_188_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_189_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_190_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_191_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_192_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_193_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_194_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_195_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_196_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_197_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_198_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_199_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_200_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_201_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_202_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_203_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_204_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_205_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_206_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_207_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_208_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_209_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_210_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_211_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_212_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_213_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_214_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_215_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_216_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_217_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_218_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_219_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_220_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_221_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_222_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_223_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_224_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_225_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_226_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_227_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_228_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_229_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_230_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_231_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_232_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_233_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_234_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_235_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_236_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_237_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_238_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_239_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_240_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_241_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_242_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_243_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_244_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_245_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_246_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_247_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_248_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_249_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_250_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_251_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_252_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_253_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_254_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_255_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_256_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_257_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_258_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_259_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_260_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_261_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_262_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_263_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_264_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_265_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_266_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_267_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_268_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_269_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_270_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_271_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_272_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_273_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_274_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_275_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_276_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_277_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_278_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_279_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_280_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_281_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_282_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_283_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_284_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_285_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_286_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_287_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_288_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_289_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_290_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_291_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_292_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_293_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_294_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_295_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_296_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_297_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_298_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_299_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_300_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_301_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_302_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_303_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_304_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_305_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_306_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_307_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_308_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_309_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_310_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_311_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_312_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_313_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_314_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_315_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_316_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_317_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_318_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_319_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_320_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_321_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_322_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_323_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_324_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_325_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_326_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_327_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_328_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_329_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_330_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_331_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_332_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout352_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout370_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2312_A (.DIODE(\line_cache[154][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2318_A (.DIODE(\line_cache[191][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3809_A (.DIODE(\fb_read_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3815_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3845_A (.DIODE(\line_cache[271][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3846_A (.DIODE(\line_cache[168][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3887_A (.DIODE(\line_cache[255][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3902_A (.DIODE(\line_cache[271][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3910_A (.DIODE(_08632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3914_A (.DIODE(\base_h_counter[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3917_A (.DIODE(\base_h_counter[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3919_A (.DIODE(\base_v_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3920_A (.DIODE(\line_cache[287][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3921_A (.DIODE(\base_h_counter[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3922_A (.DIODE(\line_cache[287][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3923_A (.DIODE(\line_cache[287][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3924_A (.DIODE(\line_cache[271][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3929_A (.DIODE(_08632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew137_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew138_A (.DIODE(_09414_));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew139_A (.DIODE(_09287_));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew141_A (.DIODE(_09494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew142_A (.DIODE(_09440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew146_A (.DIODE(_09218_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap135_A (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap136_A (.DIODE(_09504_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap140_A (.DIODE(_09283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap143_A (.DIODE(_09331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap144_A (.DIODE(_09268_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap145_A (.DIODE(_09262_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _11644_ (.A(net4266),
    .Y(_08509_));
 sky130_fd_sc_hd__inv_2 _11645_ (.A(\base_h_active[7] ),
    .Y(_08510_));
 sky130_fd_sc_hd__nor2_1 _11646_ (.A(\base_h_counter[7] ),
    .B(_08510_),
    .Y(_08511_));
 sky130_fd_sc_hd__inv_2 _11647_ (.A(net3443),
    .Y(_08512_));
 sky130_fd_sc_hd__nor2_1 _11648_ (.A(\base_h_active[7] ),
    .B(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__inv_2 _11649_ (.A(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__o21ai_1 _11650_ (.A1(_08509_),
    .A2(\base_h_active[6] ),
    .B1(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__a211oi_1 _11651_ (.A1(_08509_),
    .A2(\base_h_active[6] ),
    .B1(_08511_),
    .C1(_08515_),
    .Y(_08516_));
 sky130_fd_sc_hd__inv_2 _11652_ (.A(\base_h_active[5] ),
    .Y(_08517_));
 sky130_fd_sc_hd__nor2_1 _11653_ (.A(\base_h_counter[5] ),
    .B(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__inv_2 _11654_ (.A(net4327),
    .Y(_08519_));
 sky130_fd_sc_hd__nor2_1 _11655_ (.A(\base_h_active[5] ),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__nor2_1 _11656_ (.A(_08518_),
    .B(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__inv_2 _11657_ (.A(net3660),
    .Y(_08522_));
 sky130_fd_sc_hd__a31o_1 _11658_ (.A1(_08521_),
    .A2(\base_h_active[4] ),
    .A3(_08522_),
    .B1(_08518_),
    .X(_08523_));
 sky130_fd_sc_hd__inv_2 _11659_ (.A(net4323),
    .Y(_08524_));
 sky130_fd_sc_hd__inv_2 _11660_ (.A(\base_h_counter[0] ),
    .Y(_08525_));
 sky130_fd_sc_hd__clkbuf_4 _11661_ (.A(net4310),
    .X(_08526_));
 sky130_fd_sc_hd__inv_2 _11662_ (.A(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_08527_),
    .B(\base_h_active[1] ),
    .Y(_08528_));
 sky130_fd_sc_hd__inv_2 _11664_ (.A(\base_h_active[1] ),
    .Y(_08529_));
 sky130_fd_sc_hd__nand2_1 _11665_ (.A(_08529_),
    .B(_08526_),
    .Y(_08530_));
 sky130_fd_sc_hd__o211a_1 _11666_ (.A1(\base_h_active[0] ),
    .A2(_08525_),
    .B1(_08528_),
    .C1(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__or2b_1 _11667_ (.A(_08531_),
    .B_N(_08528_),
    .X(_08532_));
 sky130_fd_sc_hd__inv_2 _11668_ (.A(\base_h_active[2] ),
    .Y(_08533_));
 sky130_fd_sc_hd__nor2_1 _11669_ (.A(\base_h_counter[2] ),
    .B(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__inv_2 _11670_ (.A(net4320),
    .Y(_08535_));
 sky130_fd_sc_hd__nor2_1 _11671_ (.A(\base_h_active[2] ),
    .B(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__nor2_1 _11672_ (.A(_08534_),
    .B(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__nand2_1 _11673_ (.A(_08524_),
    .B(\base_h_active[3] ),
    .Y(_08538_));
 sky130_fd_sc_hd__inv_2 _11674_ (.A(\base_h_active[3] ),
    .Y(_08539_));
 sky130_fd_sc_hd__nand2_1 _11675_ (.A(_08539_),
    .B(\base_h_counter[3] ),
    .Y(_08540_));
 sky130_fd_sc_hd__and3_1 _11676_ (.A(_08537_),
    .B(_08538_),
    .C(_08540_),
    .X(_08541_));
 sky130_fd_sc_hd__and3_1 _11677_ (.A(_08534_),
    .B(_08538_),
    .C(_08540_),
    .X(_08542_));
 sky130_fd_sc_hd__a221o_1 _11678_ (.A1(_08524_),
    .A2(\base_h_active[3] ),
    .B1(_08532_),
    .B2(_08541_),
    .C1(_08542_),
    .X(_08543_));
 sky130_fd_sc_hd__nand2_1 _11679_ (.A(_08522_),
    .B(\base_h_active[4] ),
    .Y(_08544_));
 sky130_fd_sc_hd__inv_2 _11680_ (.A(\base_h_active[4] ),
    .Y(_08545_));
 sky130_fd_sc_hd__nand2_1 _11681_ (.A(_08545_),
    .B(\base_h_counter[4] ),
    .Y(_08546_));
 sky130_fd_sc_hd__and4_2 _11682_ (.A(_08516_),
    .B(_08544_),
    .C(_08546_),
    .D(_08521_),
    .X(_08547_));
 sky130_fd_sc_hd__a31o_1 _11683_ (.A1(_08514_),
    .A2(_08509_),
    .A3(\base_h_active[6] ),
    .B1(_08511_),
    .X(_08548_));
 sky130_fd_sc_hd__a221o_1 _11684_ (.A1(_08516_),
    .A2(_08523_),
    .B1(_08543_),
    .B2(_08547_),
    .C1(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__inv_2 _11685_ (.A(\base_h_active[9] ),
    .Y(_08550_));
 sky130_fd_sc_hd__nor2_1 _11686_ (.A(\base_h_counter[9] ),
    .B(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__nand2_1 _11687_ (.A(_08550_),
    .B(\base_h_counter[9] ),
    .Y(_08552_));
 sky130_fd_sc_hd__and2b_1 _11688_ (.A_N(_08551_),
    .B(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__inv_2 _11689_ (.A(net4150),
    .Y(_08554_));
 sky130_fd_sc_hd__nand2_1 _11690_ (.A(_08554_),
    .B(\base_h_active[8] ),
    .Y(_08555_));
 sky130_fd_sc_hd__or2_1 _11691_ (.A(\base_h_active[8] ),
    .B(_08554_),
    .X(_08556_));
 sky130_fd_sc_hd__and3_1 _11692_ (.A(_08553_),
    .B(_08555_),
    .C(_08556_),
    .X(_08557_));
 sky130_fd_sc_hd__a31o_1 _11693_ (.A1(_08552_),
    .A2(_08554_),
    .A3(\base_h_active[8] ),
    .B1(_08551_),
    .X(_08558_));
 sky130_fd_sc_hd__a21o_1 _11694_ (.A1(_08549_),
    .A2(_08557_),
    .B1(_08558_),
    .X(_08559_));
 sky130_fd_sc_hd__inv_2 _11695_ (.A(\base_v_active[6] ),
    .Y(_08560_));
 sky130_fd_sc_hd__nor2_1 _11696_ (.A(\base_v_counter[6] ),
    .B(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__inv_2 _11697_ (.A(net4298),
    .Y(_08562_));
 sky130_fd_sc_hd__nor2_1 _11698_ (.A(\base_v_active[6] ),
    .B(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__nor2_1 _11699_ (.A(_08561_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__inv_2 _11700_ (.A(net4321),
    .Y(_08565_));
 sky130_fd_sc_hd__nand2_1 _11701_ (.A(_08565_),
    .B(\base_v_active[7] ),
    .Y(_08566_));
 sky130_fd_sc_hd__inv_2 _11702_ (.A(\base_v_active[7] ),
    .Y(_08567_));
 sky130_fd_sc_hd__nand2_1 _11703_ (.A(_08567_),
    .B(\base_v_counter[7] ),
    .Y(_08568_));
 sky130_fd_sc_hd__and3_1 _11704_ (.A(_08564_),
    .B(_08566_),
    .C(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__inv_2 _11705_ (.A(\base_v_active[5] ),
    .Y(_08570_));
 sky130_fd_sc_hd__nor2_1 _11706_ (.A(\base_v_counter[5] ),
    .B(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__inv_2 _11707_ (.A(net4325),
    .Y(_08572_));
 sky130_fd_sc_hd__nor2_1 _11708_ (.A(\base_v_active[5] ),
    .B(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__nor2_1 _11709_ (.A(_08571_),
    .B(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__inv_2 _11710_ (.A(\base_v_active[4] ),
    .Y(_08575_));
 sky130_fd_sc_hd__nor2_1 _11711_ (.A(\base_v_counter[4] ),
    .B(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__inv_2 _11712_ (.A(net4306),
    .Y(_08577_));
 sky130_fd_sc_hd__nor2_1 _11713_ (.A(\base_v_active[4] ),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__nor2_1 _11714_ (.A(_08576_),
    .B(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__and3_1 _11715_ (.A(_08569_),
    .B(_08574_),
    .C(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__inv_2 _11716_ (.A(net4303),
    .Y(_08581_));
 sky130_fd_sc_hd__inv_2 _11717_ (.A(\base_v_active[8] ),
    .Y(_08582_));
 sky130_fd_sc_hd__nor2_1 _11718_ (.A(\base_v_counter[8] ),
    .B(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__inv_2 _11719_ (.A(net4318),
    .Y(_08584_));
 sky130_fd_sc_hd__nor2_1 _11720_ (.A(\base_v_active[8] ),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__or3_1 _11721_ (.A(\base_v_counter[9] ),
    .B(_08583_),
    .C(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__a21oi_1 _11722_ (.A1(\base_v_active[0] ),
    .A2(_08581_),
    .B1(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__inv_2 _11723_ (.A(net4300),
    .Y(_08588_));
 sky130_fd_sc_hd__nand2_1 _11724_ (.A(_08588_),
    .B(\base_v_active[3] ),
    .Y(_08589_));
 sky130_fd_sc_hd__inv_2 _11725_ (.A(\base_v_active[3] ),
    .Y(_08590_));
 sky130_fd_sc_hd__nand2_1 _11726_ (.A(_08590_),
    .B(\base_v_counter[3] ),
    .Y(_08591_));
 sky130_fd_sc_hd__nand2_1 _11727_ (.A(_08589_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__inv_2 _11728_ (.A(net4289),
    .Y(_08593_));
 sky130_fd_sc_hd__nand2_1 _11729_ (.A(_08593_),
    .B(\base_v_active[2] ),
    .Y(_08594_));
 sky130_fd_sc_hd__or2_1 _11730_ (.A(\base_v_active[2] ),
    .B(_08593_),
    .X(_08595_));
 sky130_fd_sc_hd__and3b_1 _11731_ (.A_N(_08592_),
    .B(_08594_),
    .C(_08595_),
    .X(_08596_));
 sky130_fd_sc_hd__inv_2 _11732_ (.A(\base_v_active[1] ),
    .Y(_08597_));
 sky130_fd_sc_hd__nor2_1 _11733_ (.A(\base_v_counter[1] ),
    .B(_08597_),
    .Y(_08598_));
 sky130_fd_sc_hd__inv_2 _11734_ (.A(\base_v_active[0] ),
    .Y(_08599_));
 sky130_fd_sc_hd__a22o_1 _11735_ (.A1(_08597_),
    .A2(\base_v_counter[1] ),
    .B1(_08599_),
    .B2(\base_v_counter[0] ),
    .X(_08600_));
 sky130_fd_sc_hd__nor2_1 _11736_ (.A(_08598_),
    .B(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__and2_1 _11737_ (.A(_08596_),
    .B(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__inv_2 _11738_ (.A(\base_h_active[0] ),
    .Y(_08603_));
 sky130_fd_sc_hd__o2111a_2 _11739_ (.A1(_08603_),
    .A2(\base_h_counter[0] ),
    .B1(_08531_),
    .C1(_08541_),
    .D1(_08557_),
    .X(_08604_));
 sky130_fd_sc_hd__a32o_1 _11740_ (.A1(_08580_),
    .A2(_08587_),
    .A3(_08602_),
    .B1(_08547_),
    .B2(_08604_),
    .X(_08605_));
 sky130_fd_sc_hd__inv_2 _11741_ (.A(net4229),
    .Y(_08606_));
 sky130_fd_sc_hd__a21o_1 _11742_ (.A1(_08574_),
    .A2(_08576_),
    .B1(_08571_),
    .X(_08607_));
 sky130_fd_sc_hd__o21ai_1 _11743_ (.A1(_08598_),
    .A2(_08601_),
    .B1(_08596_),
    .Y(_08608_));
 sky130_fd_sc_hd__o211ai_1 _11744_ (.A1(_08592_),
    .A2(_08594_),
    .B1(_08589_),
    .C1(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__a21bo_1 _11745_ (.A1(_08568_),
    .A2(_08561_),
    .B1_N(_08566_),
    .X(_08610_));
 sky130_fd_sc_hd__a221oi_1 _11746_ (.A1(_08569_),
    .A2(_08607_),
    .B1(_08609_),
    .B2(_08580_),
    .C1(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__o2bb2a_1 _11747_ (.A1_N(_08606_),
    .A2_N(_08583_),
    .B1(_08586_),
    .B2(_08611_),
    .X(_08612_));
 sky130_fd_sc_hd__nor2_2 _11748_ (.A(_08605_),
    .B(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__nand2_4 _11749_ (.A(_08559_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__inv_2 _11750_ (.A(_08614_),
    .Y(_08615_));
 sky130_fd_sc_hd__inv_2 _11751_ (.A(\prescaler[2] ),
    .Y(_08616_));
 sky130_fd_sc_hd__nor2_1 _11752_ (.A(\prescaler[0] ),
    .B(\prescaler[1] ),
    .Y(_08617_));
 sky130_fd_sc_hd__and2_1 _11753_ (.A(_08617_),
    .B(_08616_),
    .X(_08618_));
 sky130_fd_sc_hd__inv_2 _11754_ (.A(net2761),
    .Y(_08619_));
 sky130_fd_sc_hd__a211o_1 _11755_ (.A1(_08618_),
    .A2(\prescaler_counter[2] ),
    .B1(\prescaler_counter[3] ),
    .C1(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__or3_1 _11756_ (.A(\prescaler_counter[6] ),
    .B(net2762),
    .C(net2695),
    .X(_08621_));
 sky130_fd_sc_hd__a2111oi_1 _11757_ (.A1(net4314),
    .A2(_08619_),
    .B1(net4276),
    .C1(net2905),
    .D1(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__o311a_1 _11758_ (.A1(\prescaler_counter[2] ),
    .A2(_08616_),
    .A3(_08617_),
    .B1(_08620_),
    .C1(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__o21a_1 _11759_ (.A1(_08616_),
    .A2(_08617_),
    .B1(\prescaler_counter[2] ),
    .X(_08624_));
 sky130_fd_sc_hd__o22ai_1 _11760_ (.A1(net4314),
    .A2(_08619_),
    .B1(_08618_),
    .B2(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__or2_1 _11761_ (.A(\prescaler[1] ),
    .B(\prescaler_counter[1] ),
    .X(_08626_));
 sky130_fd_sc_hd__nand2_1 _11762_ (.A(\prescaler[1] ),
    .B(\prescaler_counter[1] ),
    .Y(_08627_));
 sky130_fd_sc_hd__a21o_1 _11763_ (.A1(_08626_),
    .A2(_08627_),
    .B1(\prescaler_counter[0] ),
    .X(_08628_));
 sky130_fd_sc_hd__a31o_1 _11764_ (.A1(_08626_),
    .A2(\prescaler_counter[0] ),
    .A3(_08627_),
    .B1(\prescaler[0] ),
    .X(_08629_));
 sky130_fd_sc_hd__a21bo_1 _11765_ (.A1(net3788),
    .A2(_08628_),
    .B1_N(_08629_),
    .X(_08630_));
 sky130_fd_sc_hd__inv_2 _11766_ (.A(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__nand3_4 _11767_ (.A(_08623_),
    .B(net4315),
    .C(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__inv_2 _11768_ (.A(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__inv_2 _11769_ (.A(net2655),
    .Y(_08634_));
 sky130_fd_sc_hd__nor2_1 _11770_ (.A(\resolution[0] ),
    .B(\resolution[1] ),
    .Y(_08635_));
 sky130_fd_sc_hd__inv_2 _11771_ (.A(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_1 _11772_ (.A(\resolution[0] ),
    .B(\resolution[1] ),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_1 _11773_ (.A(_08636_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__inv_2 _11774_ (.A(net2648),
    .Y(_08639_));
 sky130_fd_sc_hd__or2_1 _11775_ (.A(\resolution[0] ),
    .B(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__nand2_1 _11776_ (.A(_08639_),
    .B(\resolution[0] ),
    .Y(_08641_));
 sky130_fd_sc_hd__nor2_1 _11777_ (.A(\resolution[2] ),
    .B(_08636_),
    .Y(_08642_));
 sky130_fd_sc_hd__inv_2 _11778_ (.A(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__or2_1 _11779_ (.A(\resolution[3] ),
    .B(_08643_),
    .X(_08644_));
 sky130_fd_sc_hd__o21ai_1 _11780_ (.A1(_08634_),
    .A2(_08638_),
    .B1(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__a221oi_1 _11781_ (.A1(_08634_),
    .A2(_08638_),
    .B1(_08640_),
    .B2(_08641_),
    .C1(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__inv_2 _11782_ (.A(net1876),
    .Y(_08647_));
 sky130_fd_sc_hd__nand2_1 _11783_ (.A(_08643_),
    .B(\resolution[3] ),
    .Y(_08648_));
 sky130_fd_sc_hd__nand2_1 _11784_ (.A(_08644_),
    .B(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__xor2_1 _11785_ (.A(_08647_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__inv_2 _11786_ (.A(net1912),
    .Y(_08651_));
 sky130_fd_sc_hd__nand2_1 _11787_ (.A(_08636_),
    .B(\resolution[2] ),
    .Y(_08652_));
 sky130_fd_sc_hd__nand2_1 _11788_ (.A(_08643_),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__xor2_1 _11789_ (.A(_08651_),
    .B(_08653_),
    .X(_08654_));
 sky130_fd_sc_hd__and3_1 _11790_ (.A(_08646_),
    .B(_08650_),
    .C(_08654_),
    .X(_08655_));
 sky130_fd_sc_hd__xor2_1 _11791_ (.A(net2660),
    .B(_08638_),
    .X(_08656_));
 sky130_fd_sc_hd__xor2_1 _11792_ (.A(\resolution[0] ),
    .B(\line_double_counter[0] ),
    .X(_08657_));
 sky130_fd_sc_hd__nand2_1 _11793_ (.A(_08644_),
    .B(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__xor2_1 _11794_ (.A(\line_double_counter[2] ),
    .B(_08653_),
    .X(_08659_));
 sky130_fd_sc_hd__xor2_1 _11795_ (.A(net2680),
    .B(_08649_),
    .X(_08660_));
 sky130_fd_sc_hd__or4_4 _11796_ (.A(_08656_),
    .B(_08658_),
    .C(_08659_),
    .D(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__clkinv_4 _11797_ (.A(net3652),
    .Y(_08662_));
 sky130_fd_sc_hd__nor2_1 _11798_ (.A(\res_h_active[5] ),
    .B(\res_h_active[4] ),
    .Y(_08663_));
 sky130_fd_sc_hd__inv_2 _11799_ (.A(_08663_),
    .Y(_08664_));
 sky130_fd_sc_hd__nor2_1 _11800_ (.A(\res_h_active[3] ),
    .B(\res_h_active[2] ),
    .Y(_08665_));
 sky130_fd_sc_hd__nor2_1 _11801_ (.A(\res_h_active[1] ),
    .B(\res_h_active[0] ),
    .Y(_08666_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(_08665_),
    .B(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__nor2_1 _11803_ (.A(_08664_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__inv_2 _11804_ (.A(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__nor2_1 _11805_ (.A(\res_h_active[6] ),
    .B(_08669_),
    .Y(_08670_));
 sky130_fd_sc_hd__inv_2 _11806_ (.A(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__nor2_1 _11807_ (.A(\res_h_active[7] ),
    .B(_08671_),
    .Y(_08672_));
 sky130_fd_sc_hd__and2_1 _11808_ (.A(_08671_),
    .B(\res_h_active[7] ),
    .X(_08673_));
 sky130_fd_sc_hd__nor2_1 _11809_ (.A(_08672_),
    .B(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__xor2_1 _11810_ (.A(_08662_),
    .B(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__buf_12 _11811_ (.A(\res_h_counter[8] ),
    .X(_08676_));
 sky130_fd_sc_hd__clkinv_8 _11812_ (.A(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__buf_8 _11813_ (.A(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__nand2_1 _11814_ (.A(_08678_),
    .B(\res_h_active[8] ),
    .Y(_08679_));
 sky130_fd_sc_hd__or2_1 _11815_ (.A(\res_h_active[8] ),
    .B(_08677_),
    .X(_08680_));
 sky130_fd_sc_hd__a21oi_1 _11816_ (.A1(_08679_),
    .A2(_08680_),
    .B1(_08672_),
    .Y(_08681_));
 sky130_fd_sc_hd__inv_2 _11817_ (.A(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__nand2_1 _11818_ (.A(_08672_),
    .B(_08679_),
    .Y(_08683_));
 sky130_fd_sc_hd__inv_2 _11819_ (.A(net4288),
    .Y(_08684_));
 sky130_fd_sc_hd__or2_1 _11820_ (.A(\res_h_active[4] ),
    .B(_08667_),
    .X(_08685_));
 sky130_fd_sc_hd__nand2_1 _11821_ (.A(_08667_),
    .B(\res_h_active[4] ),
    .Y(_08686_));
 sky130_fd_sc_hd__nand2_1 _11822_ (.A(_08685_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__nor2_1 _11823_ (.A(_08684_),
    .B(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__inv_2 _11824_ (.A(_08688_),
    .Y(_08689_));
 sky130_fd_sc_hd__nand2_1 _11825_ (.A(_08687_),
    .B(_08684_),
    .Y(_08690_));
 sky130_fd_sc_hd__and4_1 _11826_ (.A(_08682_),
    .B(_08683_),
    .C(_08689_),
    .D(_08690_),
    .X(_08691_));
 sky130_fd_sc_hd__nor2_1 _11827_ (.A(\res_h_active[2] ),
    .B(_08666_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand2_1 _11828_ (.A(_08666_),
    .B(\res_h_active[2] ),
    .Y(_08693_));
 sky130_fd_sc_hd__or2b_1 _11829_ (.A(_08692_),
    .B_N(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__xor2_1 _11830_ (.A(\res_h_active[1] ),
    .B(\res_h_counter[1] ),
    .X(_08695_));
 sky130_fd_sc_hd__inv_2 _11831_ (.A(net2770),
    .Y(_08696_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(_08695_),
    .A1(_08696_),
    .S(\res_h_active[0] ),
    .X(_08697_));
 sky130_fd_sc_hd__nand2_1 _11833_ (.A(_08694_),
    .B(\res_h_counter[2] ),
    .Y(_08698_));
 sky130_fd_sc_hd__nand2_1 _11834_ (.A(_08695_),
    .B(_08696_),
    .Y(_08699_));
 sky130_fd_sc_hd__inv_2 _11835_ (.A(net1859),
    .Y(_08700_));
 sky130_fd_sc_hd__and3_1 _11836_ (.A(_08698_),
    .B(_08699_),
    .C(_08700_),
    .X(_08701_));
 sky130_fd_sc_hd__o211a_1 _11837_ (.A1(\res_h_counter[2] ),
    .A2(_08694_),
    .B1(_08697_),
    .C1(_08701_),
    .X(_08702_));
 sky130_fd_sc_hd__o31ai_1 _11838_ (.A1(\res_h_active[2] ),
    .A2(\res_h_active[1] ),
    .A3(\res_h_active[0] ),
    .B1(\res_h_active[3] ),
    .Y(_08703_));
 sky130_fd_sc_hd__nand2_1 _11839_ (.A(_08703_),
    .B(_08667_),
    .Y(_08704_));
 sky130_fd_sc_hd__inv_2 _11840_ (.A(net2785),
    .Y(_08705_));
 sky130_fd_sc_hd__nand2_1 _11841_ (.A(_08704_),
    .B(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__or2_1 _11842_ (.A(_08705_),
    .B(_08704_),
    .X(_08707_));
 sky130_fd_sc_hd__and4_1 _11843_ (.A(_08691_),
    .B(_08702_),
    .C(_08706_),
    .D(_08707_),
    .X(_08708_));
 sky130_fd_sc_hd__clkinv_4 _11844_ (.A(net2750),
    .Y(_08709_));
 sky130_fd_sc_hd__nand2_1 _11845_ (.A(_08669_),
    .B(\res_h_active[6] ),
    .Y(_08710_));
 sky130_fd_sc_hd__nand2_1 _11846_ (.A(_08671_),
    .B(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__or2_1 _11847_ (.A(_08709_),
    .B(_08711_),
    .X(_08712_));
 sky130_fd_sc_hd__inv_2 _11848_ (.A(\res_h_counter[5] ),
    .Y(_08713_));
 sky130_fd_sc_hd__nand2_1 _11849_ (.A(_08685_),
    .B(\res_h_active[5] ),
    .Y(_08714_));
 sky130_fd_sc_hd__nand2_1 _11850_ (.A(_08714_),
    .B(_08669_),
    .Y(_08715_));
 sky130_fd_sc_hd__or2_1 _11851_ (.A(_08713_),
    .B(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__nand2_1 _11852_ (.A(_08711_),
    .B(_08709_),
    .Y(_08717_));
 sky130_fd_sc_hd__nand2_1 _11853_ (.A(_08715_),
    .B(_08713_),
    .Y(_08718_));
 sky130_fd_sc_hd__and4_1 _11854_ (.A(_08712_),
    .B(_08716_),
    .C(_08717_),
    .D(_08718_),
    .X(_08719_));
 sky130_fd_sc_hd__nand3b_4 _11855_ (.A_N(_08675_),
    .B(_08708_),
    .C(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__nor2_2 _11856_ (.A(_08661_),
    .B(_08720_),
    .Y(_08721_));
 sky130_fd_sc_hd__clkinv_4 _11857_ (.A(net49),
    .Y(_08722_));
 sky130_fd_sc_hd__buf_6 _11858_ (.A(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__a41oi_2 _11859_ (.A1(_08615_),
    .A2(_08633_),
    .A3(_08655_),
    .A4(_08721_),
    .B1(_08723_),
    .Y(_08724_));
 sky130_fd_sc_hd__buf_12 _11860_ (.A(net75),
    .X(_08725_));
 sky130_fd_sc_hd__clkbuf_16 _11861_ (.A(\fb_read_state[1] ),
    .X(_08726_));
 sky130_fd_sc_hd__nand2_8 _11862_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__buf_12 _11863_ (.A(_08727_),
    .X(_08728_));
 sky130_fd_sc_hd__inv_2 _11864_ (.A(_08665_),
    .Y(_08729_));
 sky130_fd_sc_hd__nor2_1 _11865_ (.A(_08729_),
    .B(_08664_),
    .Y(_08730_));
 sky130_fd_sc_hd__inv_2 _11866_ (.A(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__nor2_1 _11867_ (.A(\res_h_active[6] ),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__inv_2 _11868_ (.A(_08732_),
    .Y(_08733_));
 sky130_fd_sc_hd__nor2_1 _11869_ (.A(\res_h_active[7] ),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__inv_2 _11870_ (.A(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__buf_8 _11871_ (.A(\line_cache_idx[8] ),
    .X(_08736_));
 sky130_fd_sc_hd__nand2_1 _11872_ (.A(_08735_),
    .B(\res_h_active[8] ),
    .Y(_08737_));
 sky130_fd_sc_hd__inv_2 _11873_ (.A(net2927),
    .Y(_08738_));
 sky130_fd_sc_hd__nand2_1 _11874_ (.A(_08733_),
    .B(\res_h_active[7] ),
    .Y(_08739_));
 sky130_fd_sc_hd__nand2_1 _11875_ (.A(_08735_),
    .B(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__or2_1 _11876_ (.A(_08738_),
    .B(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__inv_2 _11877_ (.A(_08741_),
    .Y(_08742_));
 sky130_fd_sc_hd__nand2_1 _11878_ (.A(_08731_),
    .B(\res_h_active[6] ),
    .Y(_08743_));
 sky130_fd_sc_hd__inv_2 _11879_ (.A(net2781),
    .Y(_08744_));
 sky130_fd_sc_hd__nand2_1 _11880_ (.A(\res_h_active[3] ),
    .B(\res_h_active[2] ),
    .Y(_08745_));
 sky130_fd_sc_hd__nand2_1 _11881_ (.A(_08729_),
    .B(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__inv_2 _11882_ (.A(\line_cache_idx[2] ),
    .Y(_08747_));
 sky130_fd_sc_hd__o21ai_1 _11883_ (.A1(_08747_),
    .A2(_08692_),
    .B1(_08693_),
    .Y(_08748_));
 sky130_fd_sc_hd__nand2_1 _11884_ (.A(_08746_),
    .B(_08744_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand2_1 _11885_ (.A(_08748_),
    .B(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__o21ai_1 _11886_ (.A1(_08744_),
    .A2(_08746_),
    .B1(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__nand2_1 _11887_ (.A(_08729_),
    .B(\res_h_active[4] ),
    .Y(_08752_));
 sky130_fd_sc_hd__inv_2 _11888_ (.A(\res_h_active[4] ),
    .Y(_08753_));
 sky130_fd_sc_hd__nand2_1 _11889_ (.A(_08665_),
    .B(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__nand2_1 _11890_ (.A(_08752_),
    .B(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__inv_2 _11891_ (.A(net3791),
    .Y(_08756_));
 sky130_fd_sc_hd__nand2_1 _11892_ (.A(_08755_),
    .B(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__inv_2 _11893_ (.A(net2787),
    .Y(_08758_));
 sky130_fd_sc_hd__nand2_1 _11894_ (.A(_08754_),
    .B(\res_h_active[5] ),
    .Y(_08759_));
 sky130_fd_sc_hd__nand2_1 _11895_ (.A(_08731_),
    .B(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__o22ai_1 _11896_ (.A1(_08756_),
    .A2(_08755_),
    .B1(_08758_),
    .B2(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__a21o_1 _11897_ (.A1(_08751_),
    .A2(_08757_),
    .B1(_08761_),
    .X(_08762_));
 sky130_fd_sc_hd__a21o_1 _11898_ (.A1(_08733_),
    .A2(_08743_),
    .B1(\line_cache_idx[6] ),
    .X(_08763_));
 sky130_fd_sc_hd__nand2_1 _11899_ (.A(_08760_),
    .B(_08758_),
    .Y(_08764_));
 sky130_fd_sc_hd__and3_1 _11900_ (.A(_08762_),
    .B(_08763_),
    .C(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__a31o_1 _11901_ (.A1(\line_cache_idx[6] ),
    .A2(_08733_),
    .A3(_08743_),
    .B1(_08765_),
    .X(_08766_));
 sky130_fd_sc_hd__nand2_1 _11902_ (.A(_08740_),
    .B(_08738_),
    .Y(_08767_));
 sky130_fd_sc_hd__o221a_1 _11903_ (.A1(_08736_),
    .A2(_08737_),
    .B1(_08742_),
    .B2(_08766_),
    .C1(_08767_),
    .X(_08768_));
 sky130_fd_sc_hd__a211o_1 _11904_ (.A1(_08736_),
    .A2(_08737_),
    .B1(\line_cache_idx[9] ),
    .C1(_08768_),
    .X(_08769_));
 sky130_fd_sc_hd__o21ai_1 _11905_ (.A1(net2712),
    .A2(_08735_),
    .B1(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__or2_4 _11906_ (.A(_08728_),
    .B(net2713),
    .X(_08771_));
 sky130_fd_sc_hd__a21bo_1 _11907_ (.A1(_08724_),
    .A2(net2702),
    .B1_N(_08771_),
    .X(_02569_));
 sky130_fd_sc_hd__inv_2 _11908_ (.A(_08655_),
    .Y(_08772_));
 sky130_fd_sc_hd__nor2_2 _11909_ (.A(_08772_),
    .B(_08614_),
    .Y(_08773_));
 sky130_fd_sc_hd__nand2_8 _11910_ (.A(_08773_),
    .B(_08721_),
    .Y(_08774_));
 sky130_fd_sc_hd__buf_12 _11911_ (.A(net49),
    .X(_08775_));
 sky130_fd_sc_hd__clkbuf_16 _11912_ (.A(_08775_),
    .X(_08776_));
 sky130_fd_sc_hd__clkbuf_16 _11913_ (.A(_08776_),
    .X(_08777_));
 sky130_fd_sc_hd__buf_12 _11914_ (.A(_08725_),
    .X(_08778_));
 sky130_fd_sc_hd__o2111ai_1 _11915_ (.A1(net4316),
    .A2(_08774_),
    .B1(_08777_),
    .C1(_08778_),
    .D1(net2713),
    .Y(_08779_));
 sky130_fd_sc_hd__nand3_1 _11916_ (.A(_08682_),
    .B(_08717_),
    .C(_08683_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand3_1 _11917_ (.A(_08702_),
    .B(_08716_),
    .C(_08718_),
    .Y(_08781_));
 sky130_fd_sc_hd__nand2_1 _11918_ (.A(_08689_),
    .B(_08706_),
    .Y(_08782_));
 sky130_fd_sc_hd__nand2_1 _11919_ (.A(_08707_),
    .B(_08690_),
    .Y(_08783_));
 sky130_fd_sc_hd__or3b_1 _11920_ (.A(_08782_),
    .B(_08783_),
    .C_N(_08712_),
    .X(_08784_));
 sky130_fd_sc_hd__or4_2 _11921_ (.A(_08780_),
    .B(_08781_),
    .C(_08675_),
    .D(_08784_),
    .X(_08785_));
 sky130_fd_sc_hd__or2_1 _11922_ (.A(_08772_),
    .B(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__nor2_1 _11923_ (.A(_08725_),
    .B(_08723_),
    .Y(_08787_));
 sky130_fd_sc_hd__o311a_1 _11924_ (.A1(_08661_),
    .A2(_08786_),
    .A3(_08614_),
    .B1(_08633_),
    .C1(_08787_),
    .X(_08788_));
 sky130_fd_sc_hd__inv_2 _11925_ (.A(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__nand2_1 _11926_ (.A(_08779_),
    .B(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__buf_12 _11927_ (.A(_08726_),
    .X(_08791_));
 sky130_fd_sc_hd__nand2_2 _11928_ (.A(net4335),
    .B(net49),
    .Y(_08792_));
 sky130_fd_sc_hd__clkinv_4 _11929_ (.A(_08792_),
    .Y(_08793_));
 sky130_fd_sc_hd__inv_16 _11930_ (.A(_08725_),
    .Y(_08794_));
 sky130_fd_sc_hd__buf_12 _11931_ (.A(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__a31o_1 _11932_ (.A1(_08793_),
    .A2(_08795_),
    .A3(_08791_),
    .B1(net4215),
    .X(_08796_));
 sky130_fd_sc_hd__a21o_1 _11933_ (.A1(_08790_),
    .A2(_08791_),
    .B1(_08796_),
    .X(_02570_));
 sky130_fd_sc_hd__buf_12 _11934_ (.A(_08794_),
    .X(_08797_));
 sky130_fd_sc_hd__o211a_1 _11935_ (.A1(_08797_),
    .A2(net2713),
    .B1(_08723_),
    .C1(_08726_),
    .X(_08798_));
 sky130_fd_sc_hd__nor2_1 _11936_ (.A(net2702),
    .B(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__buf_8 _11937_ (.A(_08775_),
    .X(_08800_));
 sky130_fd_sc_hd__clkbuf_8 _11938_ (.A(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__nor2_1 _11939_ (.A(_08632_),
    .B(_08614_),
    .Y(_08802_));
 sky130_fd_sc_hd__and3_1 _11940_ (.A(_08721_),
    .B(_08791_),
    .C(_08655_),
    .X(_08803_));
 sky130_fd_sc_hd__o2111ai_1 _11941_ (.A1(_08795_),
    .A2(net2713),
    .B1(_08801_),
    .C1(_08802_),
    .D1(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__o21ai_1 _11942_ (.A1(_08724_),
    .A2(_08799_),
    .B1(net2714),
    .Y(_02571_));
 sky130_fd_sc_hd__inv_2 _11943_ (.A(\base_h_fporch[3] ),
    .Y(_08805_));
 sky130_fd_sc_hd__nand2_1 _11944_ (.A(_08539_),
    .B(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand2_1 _11945_ (.A(\base_h_active[3] ),
    .B(\base_h_fporch[3] ),
    .Y(_08807_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(_08806_),
    .B(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__inv_2 _11947_ (.A(\base_h_fporch[2] ),
    .Y(_08809_));
 sky130_fd_sc_hd__nand2_1 _11948_ (.A(_08533_),
    .B(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand2_1 _11949_ (.A(\base_h_active[2] ),
    .B(\base_h_fporch[2] ),
    .Y(_08811_));
 sky130_fd_sc_hd__nand2_1 _11950_ (.A(_08810_),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__nor2_1 _11951_ (.A(_08808_),
    .B(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_1 _11952_ (.A(\base_h_active[0] ),
    .B(\base_h_fporch[0] ),
    .Y(_08814_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(\base_h_active[1] ),
    .B(\base_h_fporch[1] ),
    .Y(_08815_));
 sky130_fd_sc_hd__nand2_1 _11954_ (.A(\base_h_active[1] ),
    .B(\base_h_fporch[1] ),
    .Y(_08816_));
 sky130_fd_sc_hd__o21ai_1 _11955_ (.A1(_08814_),
    .A2(_08815_),
    .B1(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__nand2_1 _11956_ (.A(_08813_),
    .B(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__nor2_1 _11957_ (.A(\base_h_active[3] ),
    .B(\base_h_fporch[3] ),
    .Y(_08819_));
 sky130_fd_sc_hd__o21a_1 _11958_ (.A1(_08811_),
    .A2(_08819_),
    .B1(_08807_),
    .X(_08820_));
 sky130_fd_sc_hd__nand2_1 _11959_ (.A(_08818_),
    .B(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__or2_1 _11960_ (.A(\base_h_active[4] ),
    .B(\base_h_fporch[4] ),
    .X(_08822_));
 sky130_fd_sc_hd__nand2_1 _11961_ (.A(\base_h_active[4] ),
    .B(\base_h_fporch[4] ),
    .Y(_08823_));
 sky130_fd_sc_hd__nand2_1 _11962_ (.A(_08822_),
    .B(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__inv_2 _11963_ (.A(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__nand2_1 _11964_ (.A(_08825_),
    .B(\base_h_active[5] ),
    .Y(_08826_));
 sky130_fd_sc_hd__inv_2 _11965_ (.A(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(_08821_),
    .B(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__nor2_1 _11967_ (.A(_08517_),
    .B(_08823_),
    .Y(_08829_));
 sky130_fd_sc_hd__inv_2 _11968_ (.A(_08829_),
    .Y(_08830_));
 sky130_fd_sc_hd__nand2_1 _11969_ (.A(_08828_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__nand2_1 _11970_ (.A(_08831_),
    .B(\base_h_active[6] ),
    .Y(_08832_));
 sky130_fd_sc_hd__or2_1 _11971_ (.A(_08510_),
    .B(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__inv_2 _11972_ (.A(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__or2_1 _11973_ (.A(\base_h_active[8] ),
    .B(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__nand2_1 _11974_ (.A(_08834_),
    .B(\base_h_active[8] ),
    .Y(_08836_));
 sky130_fd_sc_hd__nand2_1 _11975_ (.A(_08835_),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_08832_),
    .B(_08510_),
    .Y(_08838_));
 sky130_fd_sc_hd__nand2_1 _11977_ (.A(_08833_),
    .B(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__a21oi_2 _11978_ (.A1(_08821_),
    .A2(_08827_),
    .B1(_08829_),
    .Y(_08840_));
 sky130_fd_sc_hd__inv_2 _11979_ (.A(\base_h_active[6] ),
    .Y(_08841_));
 sky130_fd_sc_hd__nand2_1 _11980_ (.A(_08840_),
    .B(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__nand2_1 _11981_ (.A(_08842_),
    .B(_08832_),
    .Y(_08843_));
 sky130_fd_sc_hd__inv_2 _11982_ (.A(\base_h_sync[6] ),
    .Y(_08844_));
 sky130_fd_sc_hd__nand2_1 _11983_ (.A(_08843_),
    .B(_08844_),
    .Y(_08845_));
 sky130_fd_sc_hd__nand3_1 _11984_ (.A(_08842_),
    .B(\base_h_sync[6] ),
    .C(_08832_),
    .Y(_08846_));
 sky130_fd_sc_hd__nand2_1 _11985_ (.A(_08845_),
    .B(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__nor2_1 _11986_ (.A(_08839_),
    .B(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nand2_1 _11987_ (.A(_08821_),
    .B(_08825_),
    .Y(_08849_));
 sky130_fd_sc_hd__nand3_1 _11988_ (.A(_08849_),
    .B(_08517_),
    .C(_08823_),
    .Y(_08850_));
 sky130_fd_sc_hd__nand2_2 _11989_ (.A(_08850_),
    .B(_08840_),
    .Y(_08851_));
 sky130_fd_sc_hd__inv_2 _11990_ (.A(\base_h_sync[5] ),
    .Y(_08852_));
 sky130_fd_sc_hd__nand2_1 _11991_ (.A(_08851_),
    .B(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__nand3_1 _11992_ (.A(_08818_),
    .B(_08820_),
    .C(_08824_),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_1 _11993_ (.A(_08849_),
    .B(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__inv_2 _11994_ (.A(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__nand2_2 _11995_ (.A(_08856_),
    .B(\base_h_sync[4] ),
    .Y(_08857_));
 sky130_fd_sc_hd__inv_2 _11996_ (.A(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__nor2_1 _11997_ (.A(_08852_),
    .B(_08851_),
    .Y(_08859_));
 sky130_fd_sc_hd__a21oi_2 _11998_ (.A1(_08853_),
    .A2(_08858_),
    .B1(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__inv_2 _11999_ (.A(_08860_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand2_1 _12000_ (.A(_08848_),
    .B(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__or2_1 _12001_ (.A(_08846_),
    .B(_08839_),
    .X(_08863_));
 sky130_fd_sc_hd__nand2_1 _12002_ (.A(_08862_),
    .B(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__inv_2 _12003_ (.A(_08814_),
    .Y(_08865_));
 sky130_fd_sc_hd__inv_2 _12004_ (.A(\base_h_fporch[1] ),
    .Y(_08866_));
 sky130_fd_sc_hd__nand2_1 _12005_ (.A(_08529_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__nand3_2 _12006_ (.A(_08865_),
    .B(_08867_),
    .C(_08816_),
    .Y(_08868_));
 sky130_fd_sc_hd__nand2_1 _12007_ (.A(_08866_),
    .B(\base_h_active[1] ),
    .Y(_08869_));
 sky130_fd_sc_hd__nand2_1 _12008_ (.A(_08529_),
    .B(\base_h_fporch[1] ),
    .Y(_08870_));
 sky130_fd_sc_hd__nand3_1 _12009_ (.A(_08869_),
    .B(_08870_),
    .C(_08814_),
    .Y(_08871_));
 sky130_fd_sc_hd__nand2_1 _12010_ (.A(_08868_),
    .B(_08871_),
    .Y(_08872_));
 sky130_fd_sc_hd__inv_2 _12011_ (.A(\base_h_sync[1] ),
    .Y(_08873_));
 sky130_fd_sc_hd__nand2_1 _12012_ (.A(_08872_),
    .B(_08873_),
    .Y(_08874_));
 sky130_fd_sc_hd__nand3_1 _12013_ (.A(_08868_),
    .B(_08871_),
    .C(\base_h_sync[1] ),
    .Y(_08875_));
 sky130_fd_sc_hd__nor2_1 _12014_ (.A(\base_h_active[0] ),
    .B(\base_h_fporch[0] ),
    .Y(_08876_));
 sky130_fd_sc_hd__nor2_1 _12015_ (.A(_08876_),
    .B(_08865_),
    .Y(_08877_));
 sky130_fd_sc_hd__nand2_1 _12016_ (.A(_08877_),
    .B(\base_h_sync[0] ),
    .Y(_08878_));
 sky130_fd_sc_hd__inv_2 _12017_ (.A(_08878_),
    .Y(_08879_));
 sky130_fd_sc_hd__nand3_1 _12018_ (.A(_08874_),
    .B(_08875_),
    .C(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__nand2_1 _12019_ (.A(_08880_),
    .B(_08875_),
    .Y(_08881_));
 sky130_fd_sc_hd__nand3_1 _12020_ (.A(_08868_),
    .B(_08816_),
    .C(_08812_),
    .Y(_08882_));
 sky130_fd_sc_hd__inv_2 _12021_ (.A(_08812_),
    .Y(_08883_));
 sky130_fd_sc_hd__nand2_2 _12022_ (.A(_08817_),
    .B(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__nand2_1 _12023_ (.A(_08882_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__nand2_1 _12024_ (.A(_08885_),
    .B(\base_h_sync[2] ),
    .Y(_08886_));
 sky130_fd_sc_hd__inv_2 _12025_ (.A(\base_h_sync[2] ),
    .Y(_08887_));
 sky130_fd_sc_hd__nand3_1 _12026_ (.A(_08882_),
    .B(_08887_),
    .C(_08884_),
    .Y(_08888_));
 sky130_fd_sc_hd__nand2_1 _12027_ (.A(_08886_),
    .B(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__nand2_2 _12028_ (.A(_08881_),
    .B(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__nand3_2 _12029_ (.A(_08882_),
    .B(\base_h_sync[2] ),
    .C(_08884_),
    .Y(_08891_));
 sky130_fd_sc_hd__nand2_1 _12030_ (.A(_08890_),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__nand2_1 _12031_ (.A(_08884_),
    .B(_08811_),
    .Y(_08893_));
 sky130_fd_sc_hd__inv_2 _12032_ (.A(_08808_),
    .Y(_08894_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_08893_),
    .B(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__nand3_1 _12034_ (.A(_08884_),
    .B(_08808_),
    .C(_08811_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand2_1 _12035_ (.A(_08895_),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__inv_2 _12036_ (.A(\base_h_sync[3] ),
    .Y(_08898_));
 sky130_fd_sc_hd__nand2_1 _12037_ (.A(_08897_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__nand2_1 _12038_ (.A(_08892_),
    .B(_08899_),
    .Y(_08900_));
 sky130_fd_sc_hd__nand3_2 _12039_ (.A(_08895_),
    .B(\base_h_sync[3] ),
    .C(_08896_),
    .Y(_08901_));
 sky130_fd_sc_hd__nand2_1 _12040_ (.A(_08900_),
    .B(_08901_),
    .Y(_08902_));
 sky130_fd_sc_hd__xor2_1 _12041_ (.A(\base_h_sync[4] ),
    .B(_08855_),
    .X(_08903_));
 sky130_fd_sc_hd__inv_2 _12042_ (.A(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__nand2_1 _12043_ (.A(_08851_),
    .B(\base_h_sync[5] ),
    .Y(_08905_));
 sky130_fd_sc_hd__nand3_1 _12044_ (.A(_08850_),
    .B(_08840_),
    .C(_08852_),
    .Y(_08906_));
 sky130_fd_sc_hd__nand2_1 _12045_ (.A(_08905_),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_1 _12046_ (.A(_08904_),
    .B(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__inv_2 _12047_ (.A(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__nand3_1 _12048_ (.A(_08848_),
    .B(_08902_),
    .C(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__inv_2 _12049_ (.A(_08910_),
    .Y(_08911_));
 sky130_fd_sc_hd__nor2_1 _12050_ (.A(_08864_),
    .B(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__or2_1 _12051_ (.A(_08837_),
    .B(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__nand2_1 _12052_ (.A(_08912_),
    .B(_08837_),
    .Y(_08914_));
 sky130_fd_sc_hd__nand2_1 _12053_ (.A(_08913_),
    .B(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__inv_2 _12054_ (.A(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__xor2_1 _12055_ (.A(\base_h_active[9] ),
    .B(_08836_),
    .X(_08917_));
 sky130_fd_sc_hd__inv_2 _12056_ (.A(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__xor2_2 _12057_ (.A(_08918_),
    .B(_08913_),
    .X(_08919_));
 sky130_fd_sc_hd__inv_2 _12058_ (.A(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__inv_2 _12059_ (.A(net2896),
    .Y(_08921_));
 sky130_fd_sc_hd__a22o_1 _12060_ (.A1(_08554_),
    .A2(_08916_),
    .B1(_08920_),
    .B2(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__nand3_1 _12061_ (.A(_08902_),
    .B(_08907_),
    .C(_08904_),
    .Y(_08923_));
 sky130_fd_sc_hd__nand2_1 _12062_ (.A(_08923_),
    .B(_08860_),
    .Y(_08924_));
 sky130_fd_sc_hd__inv_2 _12063_ (.A(_08847_),
    .Y(_08925_));
 sky130_fd_sc_hd__nand2_1 _12064_ (.A(_08924_),
    .B(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__nand3_1 _12065_ (.A(_08926_),
    .B(_08839_),
    .C(_08846_),
    .Y(_08927_));
 sky130_fd_sc_hd__nand2_2 _12066_ (.A(_08927_),
    .B(_08912_),
    .Y(_08928_));
 sky130_fd_sc_hd__inv_2 _12067_ (.A(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__nand2_1 _12068_ (.A(_08929_),
    .B(_08512_),
    .Y(_08930_));
 sky130_fd_sc_hd__nand2_2 _12069_ (.A(_08902_),
    .B(_08904_),
    .Y(_08931_));
 sky130_fd_sc_hd__nand2_1 _12070_ (.A(_08931_),
    .B(_08857_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand2_1 _12071_ (.A(_08932_),
    .B(_08907_),
    .Y(_08933_));
 sky130_fd_sc_hd__inv_2 _12072_ (.A(_08907_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand3_2 _12073_ (.A(_08931_),
    .B(_08934_),
    .C(_08857_),
    .Y(_08935_));
 sky130_fd_sc_hd__nand2_1 _12074_ (.A(_08933_),
    .B(_08935_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand3_1 _12075_ (.A(_08900_),
    .B(_08903_),
    .C(_08901_),
    .Y(_08937_));
 sky130_fd_sc_hd__nand2_1 _12076_ (.A(_08931_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__nand2_1 _12077_ (.A(_08885_),
    .B(_08887_),
    .Y(_08939_));
 sky130_fd_sc_hd__nand2_1 _12078_ (.A(_08939_),
    .B(_08891_),
    .Y(_08940_));
 sky130_fd_sc_hd__a21boi_1 _12079_ (.A1(_08874_),
    .A2(_08879_),
    .B1_N(_08875_),
    .Y(_08941_));
 sky130_fd_sc_hd__nand2_1 _12080_ (.A(_08940_),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(_08890_),
    .B(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand3_1 _12082_ (.A(_08892_),
    .B(_08901_),
    .C(_08899_),
    .Y(_08944_));
 sky130_fd_sc_hd__nand2_1 _12083_ (.A(_08899_),
    .B(_08901_),
    .Y(_08945_));
 sky130_fd_sc_hd__nand3_1 _12084_ (.A(_08945_),
    .B(_08891_),
    .C(_08890_),
    .Y(_08946_));
 sky130_fd_sc_hd__nand2_1 _12085_ (.A(_08944_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(_08872_),
    .B(\base_h_sync[1] ),
    .Y(_08948_));
 sky130_fd_sc_hd__nand3_1 _12087_ (.A(_08868_),
    .B(_08871_),
    .C(_08873_),
    .Y(_08949_));
 sky130_fd_sc_hd__nand3_1 _12088_ (.A(_08948_),
    .B(_08949_),
    .C(_08878_),
    .Y(_08950_));
 sky130_fd_sc_hd__nand2_1 _12089_ (.A(_08880_),
    .B(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__nand2_1 _12090_ (.A(_08951_),
    .B(_08526_),
    .Y(_08952_));
 sky130_fd_sc_hd__or2_1 _12091_ (.A(\base_h_sync[0] ),
    .B(_08877_),
    .X(_08953_));
 sky130_fd_sc_hd__nand2_1 _12092_ (.A(_08953_),
    .B(_08878_),
    .Y(_08954_));
 sky130_fd_sc_hd__inv_2 _12093_ (.A(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__nor2_1 _12094_ (.A(_08526_),
    .B(_08951_),
    .Y(_08956_));
 sky130_fd_sc_hd__a31o_1 _12095_ (.A1(_08952_),
    .A2(_08525_),
    .A3(_08955_),
    .B1(_08956_),
    .X(_08957_));
 sky130_fd_sc_hd__nand2_1 _12096_ (.A(_08943_),
    .B(\base_h_counter[2] ),
    .Y(_08958_));
 sky130_fd_sc_hd__nand2_1 _12097_ (.A(_08957_),
    .B(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__o221ai_1 _12098_ (.A1(\base_h_counter[2] ),
    .A2(_08943_),
    .B1(\base_h_counter[3] ),
    .B2(_08947_),
    .C1(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__nand2_1 _12099_ (.A(_08938_),
    .B(\base_h_counter[4] ),
    .Y(_08961_));
 sky130_fd_sc_hd__nand2_1 _12100_ (.A(_08947_),
    .B(\base_h_counter[3] ),
    .Y(_08962_));
 sky130_fd_sc_hd__nand3_1 _12101_ (.A(_08960_),
    .B(_08961_),
    .C(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__o221ai_2 _12102_ (.A1(\base_h_counter[5] ),
    .A2(_08936_),
    .B1(\base_h_counter[4] ),
    .B2(_08938_),
    .C1(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand3_1 _12103_ (.A(_08923_),
    .B(_08847_),
    .C(_08860_),
    .Y(_08965_));
 sky130_fd_sc_hd__nand2_1 _12104_ (.A(_08926_),
    .B(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__nand2_1 _12105_ (.A(_08966_),
    .B(\base_h_counter[6] ),
    .Y(_08967_));
 sky130_fd_sc_hd__nand2_1 _12106_ (.A(_08936_),
    .B(\base_h_counter[5] ),
    .Y(_08968_));
 sky130_fd_sc_hd__nand3_1 _12107_ (.A(_08964_),
    .B(_08967_),
    .C(_08968_),
    .Y(_08969_));
 sky130_fd_sc_hd__or2_1 _12108_ (.A(\base_h_counter[6] ),
    .B(_08966_),
    .X(_08970_));
 sky130_fd_sc_hd__a22o_1 _12109_ (.A1(\base_h_counter[7] ),
    .A2(_08928_),
    .B1(_08969_),
    .B2(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__o2bb2a_1 _12110_ (.A1_N(_08930_),
    .A2_N(_08971_),
    .B1(_08554_),
    .B2(_08916_),
    .X(_08972_));
 sky130_fd_sc_hd__nand2_1 _12111_ (.A(_08919_),
    .B(\base_h_counter[9] ),
    .Y(_08973_));
 sky130_fd_sc_hd__or2_1 _12112_ (.A(\base_h_counter[8] ),
    .B(_08837_),
    .X(_08974_));
 sky130_fd_sc_hd__a2bb2o_1 _12113_ (.A1_N(\base_h_counter[5] ),
    .A2_N(_08851_),
    .B1(_08522_),
    .B2(_08856_),
    .X(_08975_));
 sky130_fd_sc_hd__and2_1 _12114_ (.A(_08885_),
    .B(\base_h_counter[2] ),
    .X(_08976_));
 sky130_fd_sc_hd__nand2_1 _12115_ (.A(_08872_),
    .B(_08526_),
    .Y(_08977_));
 sky130_fd_sc_hd__and3_1 _12116_ (.A(_08977_),
    .B(_08525_),
    .C(_08877_),
    .X(_08978_));
 sky130_fd_sc_hd__o21ba_1 _12117_ (.A1(_08526_),
    .A2(_08872_),
    .B1_N(_08978_),
    .X(_08979_));
 sky130_fd_sc_hd__or2_1 _12118_ (.A(\base_h_counter[3] ),
    .B(_08897_),
    .X(_08980_));
 sky130_fd_sc_hd__or2_1 _12119_ (.A(\base_h_counter[2] ),
    .B(_08885_),
    .X(_08981_));
 sky130_fd_sc_hd__o211ai_1 _12120_ (.A1(_08976_),
    .A2(_08979_),
    .B1(_08980_),
    .C1(_08981_),
    .Y(_08982_));
 sky130_fd_sc_hd__nand2_1 _12121_ (.A(_08897_),
    .B(\base_h_counter[3] ),
    .Y(_08983_));
 sky130_fd_sc_hd__nand2_1 _12122_ (.A(_08855_),
    .B(\base_h_counter[4] ),
    .Y(_08984_));
 sky130_fd_sc_hd__a21o_1 _12123_ (.A1(_08983_),
    .A2(_08984_),
    .B1(_08975_),
    .X(_08985_));
 sky130_fd_sc_hd__nand2_1 _12124_ (.A(_08851_),
    .B(\base_h_counter[5] ),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_1 _12125_ (.A(_08843_),
    .B(\base_h_counter[6] ),
    .Y(_08987_));
 sky130_fd_sc_hd__o2111ai_1 _12126_ (.A1(_08975_),
    .A2(_08982_),
    .B1(_08985_),
    .C1(_08986_),
    .D1(_08987_),
    .Y(_08988_));
 sky130_fd_sc_hd__or2_1 _12127_ (.A(\base_h_counter[6] ),
    .B(_08843_),
    .X(_08989_));
 sky130_fd_sc_hd__a22o_1 _12128_ (.A1(\base_h_counter[7] ),
    .A2(_08839_),
    .B1(_08988_),
    .B2(_08989_),
    .X(_08990_));
 sky130_fd_sc_hd__or2_1 _12129_ (.A(\base_h_counter[7] ),
    .B(_08839_),
    .X(_08991_));
 sky130_fd_sc_hd__a22o_1 _12130_ (.A1(\base_h_counter[8] ),
    .A2(_08837_),
    .B1(_08990_),
    .B2(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__o211ai_1 _12131_ (.A1(\base_h_counter[9] ),
    .A2(_08917_),
    .B1(_08974_),
    .C1(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__o21ai_1 _12132_ (.A1(_08921_),
    .A2(_08918_),
    .B1(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__o211a_4 _12133_ (.A1(_08922_),
    .A2(_08972_),
    .B1(_08973_),
    .C1(_08994_),
    .X(net92));
 sky130_fd_sc_hd__nand2_1 _12134_ (.A(\base_v_active[0] ),
    .B(\base_v_fporch[0] ),
    .Y(_08995_));
 sky130_fd_sc_hd__inv_2 _12135_ (.A(\base_v_fporch[1] ),
    .Y(_08996_));
 sky130_fd_sc_hd__nand2_1 _12136_ (.A(_08597_),
    .B(_08996_),
    .Y(_08997_));
 sky130_fd_sc_hd__nand2_1 _12137_ (.A(\base_v_active[1] ),
    .B(\base_v_fporch[1] ),
    .Y(_08998_));
 sky130_fd_sc_hd__nand2_1 _12138_ (.A(_08997_),
    .B(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__or2_1 _12139_ (.A(_08995_),
    .B(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__nand2_1 _12140_ (.A(_09000_),
    .B(_08998_),
    .Y(_09001_));
 sky130_fd_sc_hd__or2_1 _12141_ (.A(\base_v_active[2] ),
    .B(\base_v_fporch[2] ),
    .X(_09002_));
 sky130_fd_sc_hd__nand2_1 _12142_ (.A(\base_v_active[2] ),
    .B(\base_v_fporch[2] ),
    .Y(_09003_));
 sky130_fd_sc_hd__nand2_1 _12143_ (.A(_09002_),
    .B(_09003_),
    .Y(_09004_));
 sky130_fd_sc_hd__inv_2 _12144_ (.A(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__nand2_1 _12145_ (.A(_09001_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__and2_1 _12146_ (.A(_09006_),
    .B(_09003_),
    .X(_09007_));
 sky130_fd_sc_hd__nand3b_2 _12147_ (.A_N(_09007_),
    .B(\base_v_active[4] ),
    .C(\base_v_active[3] ),
    .Y(_09008_));
 sky130_fd_sc_hd__nor2_1 _12148_ (.A(_08570_),
    .B(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__inv_2 _12149_ (.A(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__nand2_1 _12150_ (.A(_09008_),
    .B(_08570_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_1 _12151_ (.A(_09010_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__inv_2 _12152_ (.A(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__nand2_1 _12153_ (.A(_09013_),
    .B(_08572_),
    .Y(_09014_));
 sky130_fd_sc_hd__nand2_1 _12154_ (.A(_09012_),
    .B(\base_v_counter[5] ),
    .Y(_09015_));
 sky130_fd_sc_hd__nand2_1 _12155_ (.A(_09014_),
    .B(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__or2_1 _12156_ (.A(_08590_),
    .B(_09007_),
    .X(_09017_));
 sky130_fd_sc_hd__nand2_1 _12157_ (.A(_09017_),
    .B(_08575_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand2_1 _12158_ (.A(_09018_),
    .B(_09008_),
    .Y(_09019_));
 sky130_fd_sc_hd__or2_1 _12159_ (.A(\base_v_counter[4] ),
    .B(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__nand2_1 _12160_ (.A(_09019_),
    .B(\base_v_counter[4] ),
    .Y(_09021_));
 sky130_fd_sc_hd__nand2_1 _12161_ (.A(_09020_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__nand2_1 _12162_ (.A(_09010_),
    .B(_08560_),
    .Y(_09023_));
 sky130_fd_sc_hd__nand2_1 _12163_ (.A(_09009_),
    .B(\base_v_active[6] ),
    .Y(_09024_));
 sky130_fd_sc_hd__nand2_1 _12164_ (.A(_09023_),
    .B(_09024_),
    .Y(_09025_));
 sky130_fd_sc_hd__inv_2 _12165_ (.A(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__nor2_1 _12166_ (.A(_08562_),
    .B(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__nand2_1 _12167_ (.A(_09024_),
    .B(_08567_),
    .Y(_09028_));
 sky130_fd_sc_hd__nand3_1 _12168_ (.A(_09009_),
    .B(\base_v_active[7] ),
    .C(\base_v_active[6] ),
    .Y(_09029_));
 sky130_fd_sc_hd__nand2_1 _12169_ (.A(_09028_),
    .B(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__xor2_1 _12170_ (.A(\base_v_counter[7] ),
    .B(_09030_),
    .X(_09031_));
 sky130_fd_sc_hd__inv_2 _12171_ (.A(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__nand2_1 _12172_ (.A(_09026_),
    .B(_08562_),
    .Y(_09033_));
 sky130_fd_sc_hd__or3b_1 _12173_ (.A(_09027_),
    .B(_09032_),
    .C_N(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__nor3_1 _12174_ (.A(_09016_),
    .B(_09022_),
    .C(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__nand2_1 _12175_ (.A(_08999_),
    .B(_08995_),
    .Y(_09036_));
 sky130_fd_sc_hd__nand2_1 _12176_ (.A(_09000_),
    .B(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__or2_1 _12177_ (.A(\base_v_active[0] ),
    .B(\base_v_fporch[0] ),
    .X(_09038_));
 sky130_fd_sc_hd__nand2_1 _12178_ (.A(_09038_),
    .B(_08995_),
    .Y(_09039_));
 sky130_fd_sc_hd__inv_2 _12179_ (.A(_09037_),
    .Y(_09040_));
 sky130_fd_sc_hd__inv_2 _12180_ (.A(net4312),
    .Y(_09041_));
 sky130_fd_sc_hd__a22o_1 _12181_ (.A1(\base_v_counter[0] ),
    .A2(_09039_),
    .B1(_09040_),
    .B2(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__a21o_1 _12182_ (.A1(\base_v_counter[1] ),
    .A2(_09037_),
    .B1(_09042_),
    .X(_09043_));
 sky130_fd_sc_hd__nand2_1 _12183_ (.A(_09007_),
    .B(_08590_),
    .Y(_09044_));
 sky130_fd_sc_hd__nand2_1 _12184_ (.A(_09017_),
    .B(_09044_),
    .Y(_09045_));
 sky130_fd_sc_hd__nor2_1 _12185_ (.A(\base_v_counter[3] ),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__inv_2 _12186_ (.A(_09045_),
    .Y(_09047_));
 sky130_fd_sc_hd__nor2_1 _12187_ (.A(_08588_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__nor2_1 _12188_ (.A(_09046_),
    .B(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__or2_1 _12189_ (.A(_09005_),
    .B(_09001_),
    .X(_09050_));
 sky130_fd_sc_hd__nand2_1 _12190_ (.A(_09050_),
    .B(_09006_),
    .Y(_09051_));
 sky130_fd_sc_hd__inv_2 _12191_ (.A(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__nand2_1 _12192_ (.A(_09052_),
    .B(_08593_),
    .Y(_09053_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(_09051_),
    .B(\base_v_counter[2] ),
    .Y(_09054_));
 sky130_fd_sc_hd__and3_1 _12194_ (.A(_09049_),
    .B(_09053_),
    .C(_09054_),
    .X(_09055_));
 sky130_fd_sc_hd__or2_1 _12195_ (.A(\base_v_counter[0] ),
    .B(_09039_),
    .X(_09056_));
 sky130_fd_sc_hd__and3b_1 _12196_ (.A_N(_09043_),
    .B(_09055_),
    .C(_09056_),
    .X(_09057_));
 sky130_fd_sc_hd__or2_1 _12197_ (.A(_08582_),
    .B(_09029_),
    .X(_09058_));
 sky130_fd_sc_hd__clkbuf_2 _12198_ (.A(_09058_),
    .X(_09059_));
 sky130_fd_sc_hd__xor2_1 _12199_ (.A(\base_v_counter[9] ),
    .B(_09059_),
    .X(_09060_));
 sky130_fd_sc_hd__nand2_1 _12200_ (.A(_09029_),
    .B(_08582_),
    .Y(_09061_));
 sky130_fd_sc_hd__nand2_1 _12201_ (.A(_09059_),
    .B(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__inv_2 _12202_ (.A(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_1 _12203_ (.A(_09063_),
    .B(_08584_),
    .Y(_09064_));
 sky130_fd_sc_hd__nand2_1 _12204_ (.A(_09062_),
    .B(\base_v_counter[8] ),
    .Y(_09065_));
 sky130_fd_sc_hd__and3_1 _12205_ (.A(_09060_),
    .B(_09064_),
    .C(_09065_),
    .X(_09066_));
 sky130_fd_sc_hd__and3_1 _12206_ (.A(_09035_),
    .B(_09057_),
    .C(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__o21a_1 _12207_ (.A1(_09020_),
    .A2(_09016_),
    .B1(_09014_),
    .X(_09068_));
 sky130_fd_sc_hd__inv_2 _12208_ (.A(_09030_),
    .Y(_09069_));
 sky130_fd_sc_hd__nand2_1 _12209_ (.A(_09069_),
    .B(_08565_),
    .Y(_09070_));
 sky130_fd_sc_hd__o221a_1 _12210_ (.A1(_09033_),
    .A2(_09032_),
    .B1(_09068_),
    .B2(_09034_),
    .C1(_09070_),
    .X(_09071_));
 sky130_fd_sc_hd__o21ai_1 _12211_ (.A1(\base_v_counter[1] ),
    .A2(_09037_),
    .B1(_09043_),
    .Y(_09072_));
 sky130_fd_sc_hd__a31o_1 _12212_ (.A1(_09049_),
    .A2(_08593_),
    .A3(_09052_),
    .B1(_09046_),
    .X(_09073_));
 sky130_fd_sc_hd__a21o_1 _12213_ (.A1(_09055_),
    .A2(_09072_),
    .B1(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__nand2_1 _12214_ (.A(_09035_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(_09071_),
    .B(_09075_),
    .Y(_09076_));
 sky130_fd_sc_hd__nor2_1 _12216_ (.A(\base_v_counter[9] ),
    .B(_09059_),
    .Y(_09077_));
 sky130_fd_sc_hd__a31o_1 _12217_ (.A1(_09060_),
    .A2(_08584_),
    .A3(_09063_),
    .B1(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__a21oi_2 _12218_ (.A1(_09076_),
    .A2(_09066_),
    .B1(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__nand2_1 _12219_ (.A(_09040_),
    .B(\base_v_sync[1] ),
    .Y(_09080_));
 sky130_fd_sc_hd__inv_2 _12220_ (.A(\base_v_sync[0] ),
    .Y(_09081_));
 sky130_fd_sc_hd__or2_1 _12221_ (.A(_09081_),
    .B(_09039_),
    .X(_09082_));
 sky130_fd_sc_hd__inv_2 _12222_ (.A(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__inv_2 _12223_ (.A(\base_v_sync[1] ),
    .Y(_09084_));
 sky130_fd_sc_hd__nand2_1 _12224_ (.A(_09037_),
    .B(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__nand3_1 _12225_ (.A(_09080_),
    .B(_09083_),
    .C(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__nand2_1 _12226_ (.A(_09086_),
    .B(_09080_),
    .Y(_09087_));
 sky130_fd_sc_hd__inv_2 _12227_ (.A(\base_v_sync[2] ),
    .Y(_09088_));
 sky130_fd_sc_hd__nand2_1 _12228_ (.A(_09051_),
    .B(_09088_),
    .Y(_09089_));
 sky130_fd_sc_hd__nand3_2 _12229_ (.A(_09050_),
    .B(\base_v_sync[2] ),
    .C(_09006_),
    .Y(_09090_));
 sky130_fd_sc_hd__nand3_2 _12230_ (.A(_09087_),
    .B(_09089_),
    .C(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__nand2_1 _12231_ (.A(_09091_),
    .B(_09090_),
    .Y(_09092_));
 sky130_fd_sc_hd__nand2_2 _12232_ (.A(_09092_),
    .B(_09047_),
    .Y(_09093_));
 sky130_fd_sc_hd__or2_1 _12233_ (.A(_09019_),
    .B(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__nand2_1 _12234_ (.A(_09093_),
    .B(_09019_),
    .Y(_09095_));
 sky130_fd_sc_hd__nand2_1 _12235_ (.A(_09094_),
    .B(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__inv_2 _12236_ (.A(_09096_),
    .Y(_09097_));
 sky130_fd_sc_hd__nor2_1 _12237_ (.A(_08577_),
    .B(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__nor2_1 _12238_ (.A(\base_v_counter[4] ),
    .B(_09096_),
    .Y(_09099_));
 sky130_fd_sc_hd__nand2_1 _12239_ (.A(_09094_),
    .B(_09012_),
    .Y(_09100_));
 sky130_fd_sc_hd__nand3_1 _12240_ (.A(_09018_),
    .B(\base_v_active[5] ),
    .C(_09008_),
    .Y(_09101_));
 sky130_fd_sc_hd__or2_1 _12241_ (.A(_09101_),
    .B(_09093_),
    .X(_09102_));
 sky130_fd_sc_hd__nand2_1 _12242_ (.A(_09100_),
    .B(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__or2_1 _12243_ (.A(\base_v_counter[5] ),
    .B(_09103_),
    .X(_09104_));
 sky130_fd_sc_hd__nand2_1 _12244_ (.A(_09103_),
    .B(\base_v_counter[5] ),
    .Y(_09105_));
 sky130_fd_sc_hd__nand2_1 _12245_ (.A(_09104_),
    .B(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__or3_1 _12246_ (.A(_09098_),
    .B(_09099_),
    .C(_09106_),
    .X(_09107_));
 sky130_fd_sc_hd__nor2_1 _12247_ (.A(_09025_),
    .B(_09102_),
    .Y(_09108_));
 sky130_fd_sc_hd__inv_2 _12248_ (.A(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand2_1 _12249_ (.A(_09109_),
    .B(_09030_),
    .Y(_09110_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(_09108_),
    .B(_09069_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand2_1 _12251_ (.A(_09110_),
    .B(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__xor2_1 _12252_ (.A(\base_v_counter[7] ),
    .B(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__nand2_1 _12253_ (.A(_09102_),
    .B(_09025_),
    .Y(_09114_));
 sky130_fd_sc_hd__nand2_1 _12254_ (.A(_09109_),
    .B(_09114_),
    .Y(_09115_));
 sky130_fd_sc_hd__nor2_1 _12255_ (.A(\base_v_counter[6] ),
    .B(_09115_),
    .Y(_09116_));
 sky130_fd_sc_hd__inv_2 _12256_ (.A(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__nand2_1 _12257_ (.A(_09115_),
    .B(\base_v_counter[6] ),
    .Y(_09118_));
 sky130_fd_sc_hd__and3_1 _12258_ (.A(_09113_),
    .B(_09117_),
    .C(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__and2b_1 _12259_ (.A_N(_09107_),
    .B(_09119_),
    .X(_09120_));
 sky130_fd_sc_hd__or2_1 _12260_ (.A(_09062_),
    .B(_09111_),
    .X(_09121_));
 sky130_fd_sc_hd__nand2_1 _12261_ (.A(_09121_),
    .B(_09059_),
    .Y(_09122_));
 sky130_fd_sc_hd__xor2_1 _12262_ (.A(_08606_),
    .B(_09122_),
    .X(_09123_));
 sky130_fd_sc_hd__nand2_1 _12263_ (.A(_09111_),
    .B(_09062_),
    .Y(_09124_));
 sky130_fd_sc_hd__nand2_1 _12264_ (.A(_09121_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__inv_2 _12265_ (.A(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__nand2_1 _12266_ (.A(_09126_),
    .B(_08584_),
    .Y(_09127_));
 sky130_fd_sc_hd__nand2_1 _12267_ (.A(_09125_),
    .B(\base_v_counter[8] ),
    .Y(_09128_));
 sky130_fd_sc_hd__and3_1 _12268_ (.A(_09123_),
    .B(_09127_),
    .C(_09128_),
    .X(_09129_));
 sky130_fd_sc_hd__nand2_1 _12269_ (.A(_09039_),
    .B(_09081_),
    .Y(_09130_));
 sky130_fd_sc_hd__nand2_1 _12270_ (.A(_09082_),
    .B(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__inv_2 _12271_ (.A(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__nand2_1 _12272_ (.A(_09080_),
    .B(_09085_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand2_1 _12273_ (.A(_09133_),
    .B(_09082_),
    .Y(_09134_));
 sky130_fd_sc_hd__nand2_1 _12274_ (.A(_09134_),
    .B(_09086_),
    .Y(_09135_));
 sky130_fd_sc_hd__nand2_1 _12275_ (.A(_09135_),
    .B(\base_v_counter[1] ),
    .Y(_09136_));
 sky130_fd_sc_hd__or2_1 _12276_ (.A(\base_v_counter[1] ),
    .B(_09135_),
    .X(_09137_));
 sky130_fd_sc_hd__o211ai_1 _12277_ (.A1(_08581_),
    .A2(_09132_),
    .B1(_09136_),
    .C1(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__nand3_2 _12278_ (.A(_09091_),
    .B(_09045_),
    .C(_09090_),
    .Y(_09139_));
 sky130_fd_sc_hd__nand2_1 _12279_ (.A(_09093_),
    .B(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__or2_1 _12280_ (.A(\base_v_counter[3] ),
    .B(_09140_),
    .X(_09141_));
 sky130_fd_sc_hd__a21o_1 _12281_ (.A1(_09089_),
    .A2(_09090_),
    .B1(_09087_),
    .X(_09142_));
 sky130_fd_sc_hd__nand2_1 _12282_ (.A(_09142_),
    .B(_09091_),
    .Y(_09143_));
 sky130_fd_sc_hd__or2_1 _12283_ (.A(\base_v_counter[2] ),
    .B(_09143_),
    .X(_09144_));
 sky130_fd_sc_hd__nand2_1 _12284_ (.A(_09143_),
    .B(\base_v_counter[2] ),
    .Y(_09145_));
 sky130_fd_sc_hd__nand2_1 _12285_ (.A(_09140_),
    .B(\base_v_counter[3] ),
    .Y(_09146_));
 sky130_fd_sc_hd__and4_1 _12286_ (.A(_09141_),
    .B(_09144_),
    .C(_09145_),
    .D(_09146_),
    .X(_09147_));
 sky130_fd_sc_hd__inv_2 _12287_ (.A(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__a211oi_1 _12288_ (.A1(_08581_),
    .A2(_09132_),
    .B1(_09138_),
    .C1(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__nand3_1 _12289_ (.A(_09120_),
    .B(_09129_),
    .C(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__nand2_1 _12290_ (.A(_09141_),
    .B(_09146_),
    .Y(_09151_));
 sky130_fd_sc_hd__and2_1 _12291_ (.A(_09138_),
    .B(_09137_),
    .X(_09152_));
 sky130_fd_sc_hd__o221ai_2 _12292_ (.A1(_09144_),
    .A2(_09151_),
    .B1(_09152_),
    .B2(_09148_),
    .C1(_09141_),
    .Y(_09153_));
 sky130_fd_sc_hd__nand2_1 _12293_ (.A(_09113_),
    .B(_09116_),
    .Y(_09154_));
 sky130_fd_sc_hd__a21bo_1 _12294_ (.A1(_09099_),
    .A2(_09105_),
    .B1_N(_09104_),
    .X(_09155_));
 sky130_fd_sc_hd__nand2_1 _12295_ (.A(_09119_),
    .B(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__o211ai_1 _12296_ (.A1(\base_v_counter[7] ),
    .A2(_09112_),
    .B1(_09154_),
    .C1(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__a21o_1 _12297_ (.A1(_09153_),
    .A2(_09120_),
    .B1(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__inv_2 _12298_ (.A(_09122_),
    .Y(_09159_));
 sky130_fd_sc_hd__nor2_1 _12299_ (.A(\base_v_counter[9] ),
    .B(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__a31o_1 _12300_ (.A1(_09123_),
    .A2(_08584_),
    .A3(_09126_),
    .B1(_09160_),
    .X(_09161_));
 sky130_fd_sc_hd__a21o_1 _12301_ (.A1(_09158_),
    .A2(_09129_),
    .B1(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__o211ai_4 _12302_ (.A1(_09067_),
    .A2(_09079_),
    .B1(_09150_),
    .C1(_09162_),
    .Y(_09163_));
 sky130_fd_sc_hd__inv_2 _12303_ (.A(_09163_),
    .Y(net134));
 sky130_fd_sc_hd__buf_4 _12304_ (.A(_08776_),
    .X(_09164_));
 sky130_fd_sc_hd__clkbuf_8 _12305_ (.A(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__buf_12 _12306_ (.A(_08727_),
    .X(_09166_));
 sky130_fd_sc_hd__nand2_1 _12307_ (.A(net2787),
    .B(net3791),
    .Y(_09167_));
 sky130_fd_sc_hd__inv_2 _12308_ (.A(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__nor2_1 _12309_ (.A(net2927),
    .B(net4337),
    .Y(_09169_));
 sky130_fd_sc_hd__nand2_1 _12310_ (.A(_09168_),
    .B(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__inv_2 _12311_ (.A(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__nand2_4 _12312_ (.A(net2781),
    .B(\line_cache_idx[2] ),
    .Y(_09172_));
 sky130_fd_sc_hd__inv_2 _12313_ (.A(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__and3_1 _12314_ (.A(_09171_),
    .B(\line_cache_idx[8] ),
    .C(_09173_),
    .X(_09174_));
 sky130_fd_sc_hd__inv_2 _12315_ (.A(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__nor2_1 _12316_ (.A(_09166_),
    .B(_09175_),
    .Y(_09176_));
 sky130_fd_sc_hd__inv_4 _12317_ (.A(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__buf_4 _12318_ (.A(_09177_),
    .X(_09178_));
 sky130_fd_sc_hd__inv_2 _12319_ (.A(net66),
    .Y(_09179_));
 sky130_fd_sc_hd__buf_12 _12320_ (.A(_09179_),
    .X(_09180_));
 sky130_fd_sc_hd__buf_12 _12321_ (.A(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__buf_4 _12322_ (.A(_09177_),
    .X(_09182_));
 sky130_fd_sc_hd__nor2_1 _12323_ (.A(_09181_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__a31o_1 _12324_ (.A1(_09165_),
    .A2(net483),
    .A3(_09178_),
    .B1(_09183_),
    .X(_01944_));
 sky130_fd_sc_hd__clkinv_8 _12325_ (.A(net67),
    .Y(_09184_));
 sky130_fd_sc_hd__buf_12 _12326_ (.A(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__nor2_1 _12327_ (.A(_09185_),
    .B(_09182_),
    .Y(_09186_));
 sky130_fd_sc_hd__a31o_1 _12328_ (.A1(_09165_),
    .A2(net2424),
    .A3(_09178_),
    .B1(_09186_),
    .X(_01945_));
 sky130_fd_sc_hd__inv_4 _12329_ (.A(net68),
    .Y(_09187_));
 sky130_fd_sc_hd__clkbuf_16 _12330_ (.A(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__nor2_1 _12331_ (.A(_09188_),
    .B(_09182_),
    .Y(_09189_));
 sky130_fd_sc_hd__a31o_1 _12332_ (.A1(_09165_),
    .A2(net2026),
    .A3(_09178_),
    .B1(_09189_),
    .X(_01946_));
 sky130_fd_sc_hd__buf_12 _12333_ (.A(_08794_),
    .X(_09190_));
 sky130_fd_sc_hd__nor2_4 _12334_ (.A(_09190_),
    .B(_09175_),
    .Y(_09191_));
 sky130_fd_sc_hd__inv_16 _12335_ (.A(_08726_),
    .Y(_09192_));
 sky130_fd_sc_hd__buf_8 _12336_ (.A(_09192_),
    .X(_09193_));
 sky130_fd_sc_hd__nor2_2 _12337_ (.A(net69),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__buf_12 _12338_ (.A(_09194_),
    .X(_09195_));
 sky130_fd_sc_hd__clkbuf_16 _12339_ (.A(_08800_),
    .X(_09196_));
 sky130_fd_sc_hd__nand2_1 _12340_ (.A(_09196_),
    .B(net2797),
    .Y(_09197_));
 sky130_fd_sc_hd__a22o_1 _12341_ (.A1(_09191_),
    .A2(_09195_),
    .B1(_09177_),
    .B2(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__inv_2 _12342_ (.A(_09198_),
    .Y(_01947_));
 sky130_fd_sc_hd__buf_12 _12343_ (.A(_09192_),
    .X(_09199_));
 sky130_fd_sc_hd__nor2_2 _12344_ (.A(net70),
    .B(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__buf_12 _12345_ (.A(_09200_),
    .X(_09201_));
 sky130_fd_sc_hd__nand2_1 _12346_ (.A(_09196_),
    .B(net2884),
    .Y(_09202_));
 sky130_fd_sc_hd__a22o_1 _12347_ (.A1(_09191_),
    .A2(_09201_),
    .B1(_09177_),
    .B2(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__inv_2 _12348_ (.A(_09203_),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_8 _12349_ (.A(net71),
    .B(_09199_),
    .Y(_09204_));
 sky130_fd_sc_hd__buf_12 _12350_ (.A(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__nand2_1 _12351_ (.A(_09196_),
    .B(net2818),
    .Y(_09206_));
 sky130_fd_sc_hd__a22o_1 _12352_ (.A1(_09191_),
    .A2(_09205_),
    .B1(_09177_),
    .B2(_09206_),
    .X(_09207_));
 sky130_fd_sc_hd__inv_2 _12353_ (.A(_09207_),
    .Y(_01949_));
 sky130_fd_sc_hd__inv_8 _12354_ (.A(net73),
    .Y(_09208_));
 sky130_fd_sc_hd__buf_12 _12355_ (.A(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__nor2_1 _12356_ (.A(_09209_),
    .B(_09182_),
    .Y(_09210_));
 sky130_fd_sc_hd__a31o_1 _12357_ (.A1(_09165_),
    .A2(net2161),
    .A3(_09178_),
    .B1(_09210_),
    .X(_01950_));
 sky130_fd_sc_hd__nor2_8 _12358_ (.A(net74),
    .B(_09199_),
    .Y(_09211_));
 sky130_fd_sc_hd__buf_12 _12359_ (.A(_09211_),
    .X(_09212_));
 sky130_fd_sc_hd__nand2_1 _12360_ (.A(_09196_),
    .B(net3034),
    .Y(_09213_));
 sky130_fd_sc_hd__a22o_1 _12361_ (.A1(_09191_),
    .A2(_09212_),
    .B1(_09177_),
    .B2(_09213_),
    .X(_09214_));
 sky130_fd_sc_hd__inv_2 _12362_ (.A(_09214_),
    .Y(_01951_));
 sky130_fd_sc_hd__inv_2 _12363_ (.A(net57),
    .Y(_09215_));
 sky130_fd_sc_hd__buf_12 _12364_ (.A(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__nor2_1 _12365_ (.A(_09216_),
    .B(_09182_),
    .Y(_09217_));
 sky130_fd_sc_hd__a31o_1 _12366_ (.A1(_09165_),
    .A2(net475),
    .A3(_09178_),
    .B1(_09217_),
    .X(_01936_));
 sky130_fd_sc_hd__nor2_8 _12367_ (.A(net58),
    .B(_09192_),
    .Y(_09218_));
 sky130_fd_sc_hd__buf_12 _12368_ (.A(net146),
    .X(_09219_));
 sky130_fd_sc_hd__nand2_1 _12369_ (.A(_09196_),
    .B(net2783),
    .Y(_09220_));
 sky130_fd_sc_hd__a22o_1 _12370_ (.A1(_09191_),
    .A2(_09219_),
    .B1(_09177_),
    .B2(_09220_),
    .X(_09221_));
 sky130_fd_sc_hd__inv_2 _12371_ (.A(_09221_),
    .Y(_01937_));
 sky130_fd_sc_hd__buf_12 _12372_ (.A(_08775_),
    .X(_09222_));
 sky130_fd_sc_hd__buf_8 _12373_ (.A(_09222_),
    .X(_09223_));
 sky130_fd_sc_hd__clkbuf_8 _12374_ (.A(_09223_),
    .X(_09224_));
 sky130_fd_sc_hd__inv_12 _12375_ (.A(_08727_),
    .Y(_09225_));
 sky130_fd_sc_hd__buf_12 _12376_ (.A(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__clkbuf_8 _12377_ (.A(_09226_),
    .X(_09227_));
 sky130_fd_sc_hd__and3_1 _12378_ (.A(_09174_),
    .B(net59),
    .C(_09227_),
    .X(_09228_));
 sky130_fd_sc_hd__a31o_1 _12379_ (.A1(_09178_),
    .A2(_09224_),
    .A3(net1039),
    .B1(_09228_),
    .X(_01938_));
 sky130_fd_sc_hd__inv_8 _12380_ (.A(net60),
    .Y(_09229_));
 sky130_fd_sc_hd__clkbuf_16 _12381_ (.A(_09229_),
    .X(_09230_));
 sky130_fd_sc_hd__nor2_1 _12382_ (.A(_09230_),
    .B(_09182_),
    .Y(_09231_));
 sky130_fd_sc_hd__a31o_1 _12383_ (.A1(_09165_),
    .A2(net2401),
    .A3(_09178_),
    .B1(_09231_),
    .X(_01939_));
 sky130_fd_sc_hd__inv_8 _12384_ (.A(net62),
    .Y(_09232_));
 sky130_fd_sc_hd__buf_8 _12385_ (.A(_09232_),
    .X(_09233_));
 sky130_fd_sc_hd__nor2_1 _12386_ (.A(_09233_),
    .B(_09182_),
    .Y(_09234_));
 sky130_fd_sc_hd__a31o_1 _12387_ (.A1(_09165_),
    .A2(net779),
    .A3(_09178_),
    .B1(_09234_),
    .X(_01940_));
 sky130_fd_sc_hd__inv_8 _12388_ (.A(net63),
    .Y(_09235_));
 sky130_fd_sc_hd__buf_12 _12389_ (.A(_09235_),
    .X(_09236_));
 sky130_fd_sc_hd__nor2_1 _12390_ (.A(_09236_),
    .B(_09182_),
    .Y(_09237_));
 sky130_fd_sc_hd__a31o_1 _12391_ (.A1(_09165_),
    .A2(net1812),
    .A3(_09178_),
    .B1(_09237_),
    .X(_01941_));
 sky130_fd_sc_hd__nor2_4 _12392_ (.A(net64),
    .B(_09199_),
    .Y(_09238_));
 sky130_fd_sc_hd__buf_12 _12393_ (.A(_09238_),
    .X(_09239_));
 sky130_fd_sc_hd__nand2_1 _12394_ (.A(_09196_),
    .B(net2824),
    .Y(_09240_));
 sky130_fd_sc_hd__a22o_1 _12395_ (.A1(_09191_),
    .A2(_09239_),
    .B1(_09177_),
    .B2(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__inv_2 _12396_ (.A(_09241_),
    .Y(_01942_));
 sky130_fd_sc_hd__inv_6 _12397_ (.A(net65),
    .Y(_09242_));
 sky130_fd_sc_hd__clkbuf_16 _12398_ (.A(_09242_),
    .X(_09243_));
 sky130_fd_sc_hd__nor2_1 _12399_ (.A(_09243_),
    .B(_09182_),
    .Y(_09244_));
 sky130_fd_sc_hd__a31o_1 _12400_ (.A1(_09165_),
    .A2(net1693),
    .A3(_09178_),
    .B1(_09244_),
    .X(_01943_));
 sky130_fd_sc_hd__inv_2 _12401_ (.A(net81),
    .Y(_09245_));
 sky130_fd_sc_hd__clkbuf_16 _12402_ (.A(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__nor2_1 _12403_ (.A(_09246_),
    .B(_09182_),
    .Y(_09247_));
 sky130_fd_sc_hd__a31o_1 _12404_ (.A1(_09165_),
    .A2(net671),
    .A3(_09178_),
    .B1(_09247_),
    .X(_01928_));
 sky130_fd_sc_hd__nor2_8 _12405_ (.A(net82),
    .B(_09199_),
    .Y(_09248_));
 sky130_fd_sc_hd__buf_12 _12406_ (.A(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__nand2_1 _12407_ (.A(_09196_),
    .B(net2865),
    .Y(_09250_));
 sky130_fd_sc_hd__a22o_1 _12408_ (.A1(_09191_),
    .A2(_09249_),
    .B1(_09177_),
    .B2(_09250_),
    .X(_09251_));
 sky130_fd_sc_hd__inv_2 _12409_ (.A(_09251_),
    .Y(_01929_));
 sky130_fd_sc_hd__inv_4 _12410_ (.A(net51),
    .Y(_09252_));
 sky130_fd_sc_hd__clkbuf_16 _12411_ (.A(_09252_),
    .X(_09253_));
 sky130_fd_sc_hd__nor2_1 _12412_ (.A(_09253_),
    .B(_09182_),
    .Y(_09254_));
 sky130_fd_sc_hd__a31o_1 _12413_ (.A1(_09165_),
    .A2(net2070),
    .A3(_09178_),
    .B1(_09254_),
    .X(_01930_));
 sky130_fd_sc_hd__nor2_8 _12414_ (.A(net52),
    .B(_09199_),
    .Y(_09255_));
 sky130_fd_sc_hd__buf_12 _12415_ (.A(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__nand2_1 _12416_ (.A(_09196_),
    .B(net3059),
    .Y(_09257_));
 sky130_fd_sc_hd__a22o_1 _12417_ (.A1(_09191_),
    .A2(_09256_),
    .B1(_09177_),
    .B2(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__inv_2 _12418_ (.A(_09258_),
    .Y(_01931_));
 sky130_fd_sc_hd__inv_8 _12419_ (.A(net53),
    .Y(_09259_));
 sky130_fd_sc_hd__clkbuf_16 _12420_ (.A(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__nor2_1 _12421_ (.A(_09260_),
    .B(_09182_),
    .Y(_09261_));
 sky130_fd_sc_hd__a31o_1 _12422_ (.A1(_09165_),
    .A2(net1131),
    .A3(_09182_),
    .B1(_09261_),
    .X(_01932_));
 sky130_fd_sc_hd__nor2_4 _12423_ (.A(net54),
    .B(_09192_),
    .Y(_09262_));
 sky130_fd_sc_hd__clkbuf_16 _12424_ (.A(net145),
    .X(_09263_));
 sky130_fd_sc_hd__nand2_1 _12425_ (.A(_09196_),
    .B(net2983),
    .Y(_09264_));
 sky130_fd_sc_hd__a22o_1 _12426_ (.A1(_09191_),
    .A2(_09263_),
    .B1(_09177_),
    .B2(_09264_),
    .X(_09265_));
 sky130_fd_sc_hd__inv_2 _12427_ (.A(_09265_),
    .Y(_01933_));
 sky130_fd_sc_hd__buf_8 _12428_ (.A(net55),
    .X(_09266_));
 sky130_fd_sc_hd__and3_1 _12429_ (.A(_09174_),
    .B(_09266_),
    .C(_09227_),
    .X(_09267_));
 sky130_fd_sc_hd__a31o_1 _12430_ (.A1(_09178_),
    .A2(_09224_),
    .A3(net2516),
    .B1(_09267_),
    .X(_01934_));
 sky130_fd_sc_hd__nor2_8 _12431_ (.A(net56),
    .B(_09192_),
    .Y(_09268_));
 sky130_fd_sc_hd__buf_12 _12432_ (.A(net144),
    .X(_09269_));
 sky130_fd_sc_hd__buf_4 _12433_ (.A(_08800_),
    .X(_09270_));
 sky130_fd_sc_hd__nand2_1 _12434_ (.A(_09270_),
    .B(net3169),
    .Y(_09271_));
 sky130_fd_sc_hd__a22o_1 _12435_ (.A1(_09191_),
    .A2(_09269_),
    .B1(_09177_),
    .B2(_09271_),
    .X(_09272_));
 sky130_fd_sc_hd__inv_2 _12436_ (.A(_09272_),
    .Y(_01935_));
 sky130_fd_sc_hd__clkbuf_8 _12437_ (.A(_09223_),
    .X(_09273_));
 sky130_fd_sc_hd__buf_8 _12438_ (.A(net50),
    .X(_09274_));
 sky130_fd_sc_hd__and3_1 _12439_ (.A(_09174_),
    .B(_09274_),
    .C(_09227_),
    .X(_09275_));
 sky130_fd_sc_hd__a31o_1 _12440_ (.A1(_09178_),
    .A2(_09273_),
    .A3(net2700),
    .B1(_09275_),
    .X(_01920_));
 sky130_fd_sc_hd__inv_6 _12441_ (.A(net61),
    .Y(_09276_));
 sky130_fd_sc_hd__clkbuf_16 _12442_ (.A(_09276_),
    .X(_09277_));
 sky130_fd_sc_hd__nor2_1 _12443_ (.A(_09277_),
    .B(_09182_),
    .Y(_09278_));
 sky130_fd_sc_hd__a31o_1 _12444_ (.A1(_09165_),
    .A2(net1852),
    .A3(_09182_),
    .B1(_09278_),
    .X(_01921_));
 sky130_fd_sc_hd__nor2_2 _12445_ (.A(net72),
    .B(_09193_),
    .Y(_09279_));
 sky130_fd_sc_hd__buf_12 _12446_ (.A(_09279_),
    .X(_09280_));
 sky130_fd_sc_hd__nand2_1 _12447_ (.A(_09270_),
    .B(net3258),
    .Y(_09281_));
 sky130_fd_sc_hd__a22o_1 _12448_ (.A1(_09191_),
    .A2(_09280_),
    .B1(_09177_),
    .B2(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__inv_2 _12449_ (.A(_09282_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_8 _12450_ (.A(net76),
    .B(_09199_),
    .Y(_09283_));
 sky130_fd_sc_hd__clkbuf_16 _12451_ (.A(_09283_),
    .X(_09284_));
 sky130_fd_sc_hd__nand2_1 _12452_ (.A(_09270_),
    .B(net3217),
    .Y(_09285_));
 sky130_fd_sc_hd__a22o_1 _12453_ (.A1(_09191_),
    .A2(_09284_),
    .B1(_09177_),
    .B2(_09285_),
    .X(_09286_));
 sky130_fd_sc_hd__inv_2 _12454_ (.A(_09286_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_4 _12455_ (.A(net77),
    .B(_09199_),
    .Y(_09287_));
 sky130_fd_sc_hd__buf_12 _12456_ (.A(net139),
    .X(_09288_));
 sky130_fd_sc_hd__nand2_1 _12457_ (.A(_09270_),
    .B(net3089),
    .Y(_09289_));
 sky130_fd_sc_hd__a22o_1 _12458_ (.A1(_09191_),
    .A2(_09288_),
    .B1(_09177_),
    .B2(_09289_),
    .X(_09290_));
 sky130_fd_sc_hd__inv_2 _12459_ (.A(_09290_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _12460_ (.A(_08801_),
    .B(net3626),
    .Y(_09291_));
 sky130_fd_sc_hd__or2_1 _12461_ (.A(net78),
    .B(_09166_),
    .X(_09292_));
 sky130_fd_sc_hd__clkbuf_4 _12462_ (.A(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__clkbuf_16 _12463_ (.A(_09293_),
    .X(_09294_));
 sky130_fd_sc_hd__o2bb2a_1 _12464_ (.A1_N(_09291_),
    .A2_N(_09178_),
    .B1(_09175_),
    .B2(_09294_),
    .X(_01925_));
 sky130_fd_sc_hd__nand2_1 _12465_ (.A(_08801_),
    .B(net3723),
    .Y(_09295_));
 sky130_fd_sc_hd__nor2_8 _12466_ (.A(net79),
    .B(_09166_),
    .Y(_09296_));
 sky130_fd_sc_hd__inv_6 _12467_ (.A(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__buf_6 _12468_ (.A(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__o2bb2a_1 _12469_ (.A1_N(_09295_),
    .A2_N(_09178_),
    .B1(_09175_),
    .B2(_09298_),
    .X(_01926_));
 sky130_fd_sc_hd__inv_8 _12470_ (.A(net80),
    .Y(_09299_));
 sky130_fd_sc_hd__buf_12 _12471_ (.A(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__nor2_1 _12472_ (.A(_09300_),
    .B(_09177_),
    .Y(_09301_));
 sky130_fd_sc_hd__a31o_1 _12473_ (.A1(_09165_),
    .A2(net2327),
    .A3(_09182_),
    .B1(_09301_),
    .X(_01927_));
 sky130_fd_sc_hd__buf_6 _12474_ (.A(_09222_),
    .X(_09302_));
 sky130_fd_sc_hd__clkbuf_8 _12475_ (.A(_09302_),
    .X(_09303_));
 sky130_fd_sc_hd__buf_12 _12476_ (.A(_08727_),
    .X(_09304_));
 sky130_fd_sc_hd__nor2_2 _12477_ (.A(net4336),
    .B(_08744_),
    .Y(_09305_));
 sky130_fd_sc_hd__and3_2 _12478_ (.A(_09171_),
    .B(\line_cache_idx[8] ),
    .C(_09305_),
    .X(_09306_));
 sky130_fd_sc_hd__inv_2 _12479_ (.A(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__nor2_1 _12480_ (.A(_09304_),
    .B(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__inv_2 _12481_ (.A(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__buf_4 _12482_ (.A(_09309_),
    .X(_09310_));
 sky130_fd_sc_hd__buf_4 _12483_ (.A(_09309_),
    .X(_09311_));
 sky130_fd_sc_hd__nor2_1 _12484_ (.A(_09181_),
    .B(_09311_),
    .Y(_09312_));
 sky130_fd_sc_hd__a31o_1 _12485_ (.A1(_09303_),
    .A2(net2699),
    .A3(_09310_),
    .B1(_09312_),
    .X(_01912_));
 sky130_fd_sc_hd__nor2_4 _12486_ (.A(_08795_),
    .B(_09307_),
    .Y(_09313_));
 sky130_fd_sc_hd__nor2_8 _12487_ (.A(net67),
    .B(_09192_),
    .Y(_09314_));
 sky130_fd_sc_hd__buf_12 _12488_ (.A(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__nand2_1 _12489_ (.A(_09270_),
    .B(net3403),
    .Y(_09316_));
 sky130_fd_sc_hd__a22o_1 _12490_ (.A1(_09313_),
    .A2(_09315_),
    .B1(_09311_),
    .B2(_09316_),
    .X(_09317_));
 sky130_fd_sc_hd__inv_2 _12491_ (.A(_09317_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _12492_ (.A(_09188_),
    .B(_09311_),
    .Y(_09318_));
 sky130_fd_sc_hd__a31o_1 _12493_ (.A1(_09303_),
    .A2(net697),
    .A3(_09310_),
    .B1(_09318_),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_1 _12494_ (.A(_09270_),
    .B(net2971),
    .Y(_09319_));
 sky130_fd_sc_hd__a22o_1 _12495_ (.A1(_09313_),
    .A2(_09195_),
    .B1(_09311_),
    .B2(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__inv_2 _12496_ (.A(_09320_),
    .Y(_01915_));
 sky130_fd_sc_hd__buf_8 _12497_ (.A(net70),
    .X(_09321_));
 sky130_fd_sc_hd__and3_1 _12498_ (.A(_09306_),
    .B(_09321_),
    .C(_09227_),
    .X(_09322_));
 sky130_fd_sc_hd__a31o_1 _12499_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net1435),
    .B1(_09322_),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_1 _12500_ (.A(_09270_),
    .B(net3418),
    .Y(_09323_));
 sky130_fd_sc_hd__a22o_1 _12501_ (.A1(_09313_),
    .A2(_09205_),
    .B1(_09311_),
    .B2(_09323_),
    .X(_09324_));
 sky130_fd_sc_hd__inv_2 _12502_ (.A(_09324_),
    .Y(_01917_));
 sky130_fd_sc_hd__nor2_1 _12503_ (.A(_09209_),
    .B(_09311_),
    .Y(_09325_));
 sky130_fd_sc_hd__a31o_1 _12504_ (.A1(_09303_),
    .A2(net829),
    .A3(_09310_),
    .B1(_09325_),
    .X(_01918_));
 sky130_fd_sc_hd__clkbuf_16 _12505_ (.A(net74),
    .X(_09326_));
 sky130_fd_sc_hd__and3_1 _12506_ (.A(_09306_),
    .B(_09326_),
    .C(_09227_),
    .X(_09327_));
 sky130_fd_sc_hd__a31o_1 _12507_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net2087),
    .B1(_09327_),
    .X(_01919_));
 sky130_fd_sc_hd__nor2_1 _12508_ (.A(_09216_),
    .B(_09311_),
    .Y(_09328_));
 sky130_fd_sc_hd__a31o_1 _12509_ (.A1(_09303_),
    .A2(net575),
    .A3(_09310_),
    .B1(_09328_),
    .X(_01904_));
 sky130_fd_sc_hd__nand2_1 _12510_ (.A(_09270_),
    .B(net2976),
    .Y(_09329_));
 sky130_fd_sc_hd__a22o_1 _12511_ (.A1(_09313_),
    .A2(_09219_),
    .B1(_09309_),
    .B2(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__inv_2 _12512_ (.A(_09330_),
    .Y(_01905_));
 sky130_fd_sc_hd__nor2_8 _12513_ (.A(net59),
    .B(_09192_),
    .Y(_09331_));
 sky130_fd_sc_hd__clkbuf_16 _12514_ (.A(_09331_),
    .X(_09332_));
 sky130_fd_sc_hd__nand2_1 _12515_ (.A(_09270_),
    .B(net3262),
    .Y(_09333_));
 sky130_fd_sc_hd__a22o_1 _12516_ (.A1(_09313_),
    .A2(_09332_),
    .B1(_09309_),
    .B2(_09333_),
    .X(_09334_));
 sky130_fd_sc_hd__inv_2 _12517_ (.A(_09334_),
    .Y(_01906_));
 sky130_fd_sc_hd__nor2_1 _12518_ (.A(_09230_),
    .B(_09311_),
    .Y(_09335_));
 sky130_fd_sc_hd__a31o_1 _12519_ (.A1(_09303_),
    .A2(net1796),
    .A3(_09310_),
    .B1(_09335_),
    .X(_01907_));
 sky130_fd_sc_hd__nor2_1 _12520_ (.A(_09233_),
    .B(_09311_),
    .Y(_09336_));
 sky130_fd_sc_hd__a31o_1 _12521_ (.A1(_09303_),
    .A2(net2058),
    .A3(_09311_),
    .B1(_09336_),
    .X(_01908_));
 sky130_fd_sc_hd__nor2_8 _12522_ (.A(net63),
    .B(_09199_),
    .Y(_09337_));
 sky130_fd_sc_hd__buf_12 _12523_ (.A(_09337_),
    .X(_09338_));
 sky130_fd_sc_hd__nand2_1 _12524_ (.A(_09270_),
    .B(net3132),
    .Y(_09339_));
 sky130_fd_sc_hd__a22o_1 _12525_ (.A1(_09313_),
    .A2(_09338_),
    .B1(_09309_),
    .B2(_09339_),
    .X(_09340_));
 sky130_fd_sc_hd__inv_2 _12526_ (.A(_09340_),
    .Y(_01909_));
 sky130_fd_sc_hd__clkbuf_16 _12527_ (.A(net64),
    .X(_09341_));
 sky130_fd_sc_hd__and3_1 _12528_ (.A(_09306_),
    .B(_09341_),
    .C(_09227_),
    .X(_09342_));
 sky130_fd_sc_hd__a31o_1 _12529_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net1141),
    .B1(_09342_),
    .X(_01910_));
 sky130_fd_sc_hd__nor2_1 _12530_ (.A(_09243_),
    .B(_09311_),
    .Y(_09343_));
 sky130_fd_sc_hd__a31o_1 _12531_ (.A1(_09303_),
    .A2(net1614),
    .A3(_09311_),
    .B1(_09343_),
    .X(_01911_));
 sky130_fd_sc_hd__nor2_1 _12532_ (.A(_09246_),
    .B(_09311_),
    .Y(_09344_));
 sky130_fd_sc_hd__a31o_1 _12533_ (.A1(_09303_),
    .A2(net745),
    .A3(_09311_),
    .B1(_09344_),
    .X(_01896_));
 sky130_fd_sc_hd__buf_8 _12534_ (.A(net82),
    .X(_09345_));
 sky130_fd_sc_hd__and3_1 _12535_ (.A(_09306_),
    .B(_09345_),
    .C(_09227_),
    .X(_09346_));
 sky130_fd_sc_hd__a31o_1 _12536_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net2184),
    .B1(_09346_),
    .X(_01897_));
 sky130_fd_sc_hd__nor2_8 _12537_ (.A(net51),
    .B(_09192_),
    .Y(_09347_));
 sky130_fd_sc_hd__buf_12 _12538_ (.A(_09347_),
    .X(_09348_));
 sky130_fd_sc_hd__nand2_1 _12539_ (.A(_09270_),
    .B(net3487),
    .Y(_09349_));
 sky130_fd_sc_hd__a22o_1 _12540_ (.A1(_09313_),
    .A2(_09348_),
    .B1(_09309_),
    .B2(_09349_),
    .X(_09350_));
 sky130_fd_sc_hd__inv_2 _12541_ (.A(_09350_),
    .Y(_01898_));
 sky130_fd_sc_hd__buf_8 _12542_ (.A(net52),
    .X(_09351_));
 sky130_fd_sc_hd__and3_1 _12543_ (.A(_09306_),
    .B(_09351_),
    .C(_09227_),
    .X(_09352_));
 sky130_fd_sc_hd__a31o_1 _12544_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net2085),
    .B1(_09352_),
    .X(_01899_));
 sky130_fd_sc_hd__nor2_4 _12545_ (.A(net53),
    .B(_09199_),
    .Y(_09353_));
 sky130_fd_sc_hd__buf_12 _12546_ (.A(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__nand2_1 _12547_ (.A(_09270_),
    .B(net3275),
    .Y(_09355_));
 sky130_fd_sc_hd__a22o_1 _12548_ (.A1(_09313_),
    .A2(_09354_),
    .B1(_09309_),
    .B2(_09355_),
    .X(_09356_));
 sky130_fd_sc_hd__inv_2 _12549_ (.A(_09356_),
    .Y(_01900_));
 sky130_fd_sc_hd__nand2_1 _12550_ (.A(_09270_),
    .B(net3540),
    .Y(_09357_));
 sky130_fd_sc_hd__a22o_1 _12551_ (.A1(_09313_),
    .A2(_09263_),
    .B1(_09309_),
    .B2(_09357_),
    .X(_09358_));
 sky130_fd_sc_hd__inv_2 _12552_ (.A(_09358_),
    .Y(_01901_));
 sky130_fd_sc_hd__clkbuf_16 _12553_ (.A(_09225_),
    .X(_09359_));
 sky130_fd_sc_hd__buf_4 _12554_ (.A(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__and3_1 _12555_ (.A(_09306_),
    .B(_09266_),
    .C(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__a31o_1 _12556_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net1377),
    .B1(_09361_),
    .X(_01902_));
 sky130_fd_sc_hd__nand2_1 _12557_ (.A(_09270_),
    .B(net3758),
    .Y(_09362_));
 sky130_fd_sc_hd__a22o_1 _12558_ (.A1(_09313_),
    .A2(_09269_),
    .B1(_09309_),
    .B2(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__inv_2 _12559_ (.A(_09363_),
    .Y(_01903_));
 sky130_fd_sc_hd__and3_1 _12560_ (.A(_09306_),
    .B(_09274_),
    .C(_09360_),
    .X(_09364_));
 sky130_fd_sc_hd__a31o_1 _12561_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net1973),
    .B1(_09364_),
    .X(_01888_));
 sky130_fd_sc_hd__nor2_8 _12562_ (.A(net61),
    .B(_09192_),
    .Y(_09365_));
 sky130_fd_sc_hd__buf_12 _12563_ (.A(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__nand2_1 _12564_ (.A(_09270_),
    .B(net3696),
    .Y(_09367_));
 sky130_fd_sc_hd__a22o_1 _12565_ (.A1(_09313_),
    .A2(_09366_),
    .B1(_09309_),
    .B2(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__inv_2 _12566_ (.A(_09368_),
    .Y(_01889_));
 sky130_fd_sc_hd__buf_8 _12567_ (.A(net72),
    .X(_09369_));
 sky130_fd_sc_hd__and3_1 _12568_ (.A(_09306_),
    .B(_09369_),
    .C(_09360_),
    .X(_09370_));
 sky130_fd_sc_hd__a31o_1 _12569_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net1641),
    .B1(_09370_),
    .X(_01890_));
 sky130_fd_sc_hd__nand2_1 _12570_ (.A(_09270_),
    .B(net3342),
    .Y(_09371_));
 sky130_fd_sc_hd__a22o_1 _12571_ (.A1(_09313_),
    .A2(_09284_),
    .B1(_09309_),
    .B2(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__inv_2 _12572_ (.A(_09372_),
    .Y(_01891_));
 sky130_fd_sc_hd__buf_8 _12573_ (.A(net77),
    .X(_09373_));
 sky130_fd_sc_hd__and3_1 _12574_ (.A(_09306_),
    .B(_09373_),
    .C(_09360_),
    .X(_09374_));
 sky130_fd_sc_hd__a31o_1 _12575_ (.A1(_09310_),
    .A2(_09273_),
    .A3(net1173),
    .B1(_09374_),
    .X(_01892_));
 sky130_fd_sc_hd__buf_8 _12576_ (.A(_09222_),
    .X(_09375_));
 sky130_fd_sc_hd__clkbuf_8 _12577_ (.A(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__nand2_1 _12578_ (.A(_09376_),
    .B(net3668),
    .Y(_09377_));
 sky130_fd_sc_hd__o2bb2a_1 _12579_ (.A1_N(_09377_),
    .A2_N(_09310_),
    .B1(_09294_),
    .B2(_09307_),
    .X(_01893_));
 sky130_fd_sc_hd__nand2_1 _12580_ (.A(_09376_),
    .B(net3756),
    .Y(_09378_));
 sky130_fd_sc_hd__o2bb2a_1 _12581_ (.A1_N(_09378_),
    .A2_N(_09310_),
    .B1(_09298_),
    .B2(_09307_),
    .X(_01894_));
 sky130_fd_sc_hd__nor2_1 _12582_ (.A(_09300_),
    .B(_09311_),
    .Y(_09379_));
 sky130_fd_sc_hd__a31o_1 _12583_ (.A1(_09303_),
    .A2(net817),
    .A3(_09311_),
    .B1(_09379_),
    .X(_01895_));
 sky130_fd_sc_hd__nor2_2 _12584_ (.A(net2781),
    .B(_08747_),
    .Y(_09380_));
 sky130_fd_sc_hd__and3_2 _12585_ (.A(_09171_),
    .B(_08736_),
    .C(_09380_),
    .X(_09381_));
 sky130_fd_sc_hd__inv_2 _12586_ (.A(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__nor2_1 _12587_ (.A(_09166_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__clkinv_4 _12588_ (.A(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__buf_4 _12589_ (.A(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__buf_4 _12590_ (.A(_09384_),
    .X(_09386_));
 sky130_fd_sc_hd__nor2_1 _12591_ (.A(_09181_),
    .B(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__a31o_1 _12592_ (.A1(_09303_),
    .A2(net2638),
    .A3(_09385_),
    .B1(_09387_),
    .X(_01880_));
 sky130_fd_sc_hd__nor2_1 _12593_ (.A(_09185_),
    .B(_09386_),
    .Y(_09388_));
 sky130_fd_sc_hd__a31o_1 _12594_ (.A1(_09303_),
    .A2(net1089),
    .A3(_09385_),
    .B1(_09388_),
    .X(_01881_));
 sky130_fd_sc_hd__nor2_1 _12595_ (.A(_09188_),
    .B(_09386_),
    .Y(_09389_));
 sky130_fd_sc_hd__a31o_1 _12596_ (.A1(_09303_),
    .A2(net1209),
    .A3(_09385_),
    .B1(_09389_),
    .X(_01882_));
 sky130_fd_sc_hd__nor2_4 _12597_ (.A(_08795_),
    .B(_09382_),
    .Y(_09390_));
 sky130_fd_sc_hd__buf_4 _12598_ (.A(_08800_),
    .X(_09391_));
 sky130_fd_sc_hd__nand2_1 _12599_ (.A(_09391_),
    .B(net3128),
    .Y(_09392_));
 sky130_fd_sc_hd__a22o_1 _12600_ (.A1(_09390_),
    .A2(_09195_),
    .B1(_09384_),
    .B2(_09392_),
    .X(_09393_));
 sky130_fd_sc_hd__inv_2 _12601_ (.A(_09393_),
    .Y(_01883_));
 sky130_fd_sc_hd__and3_1 _12602_ (.A(_09381_),
    .B(_09321_),
    .C(_09360_),
    .X(_09394_));
 sky130_fd_sc_hd__a31o_1 _12603_ (.A1(_09385_),
    .A2(_09273_),
    .A3(net1415),
    .B1(_09394_),
    .X(_01884_));
 sky130_fd_sc_hd__buf_8 _12604_ (.A(net71),
    .X(_09395_));
 sky130_fd_sc_hd__and3_1 _12605_ (.A(_09381_),
    .B(_09395_),
    .C(_09360_),
    .X(_09396_));
 sky130_fd_sc_hd__a31o_1 _12606_ (.A1(_09385_),
    .A2(_09273_),
    .A3(net2513),
    .B1(_09396_),
    .X(_01885_));
 sky130_fd_sc_hd__nor2_2 _12607_ (.A(net73),
    .B(_09199_),
    .Y(_09397_));
 sky130_fd_sc_hd__buf_12 _12608_ (.A(_09397_),
    .X(_09398_));
 sky130_fd_sc_hd__nand2_1 _12609_ (.A(_09391_),
    .B(net3747),
    .Y(_09399_));
 sky130_fd_sc_hd__a22o_1 _12610_ (.A1(_09390_),
    .A2(_09398_),
    .B1(_09384_),
    .B2(_09399_),
    .X(_09400_));
 sky130_fd_sc_hd__inv_2 _12611_ (.A(_09400_),
    .Y(_01886_));
 sky130_fd_sc_hd__and3_1 _12612_ (.A(_09381_),
    .B(_09326_),
    .C(_09360_),
    .X(_09401_));
 sky130_fd_sc_hd__a31o_1 _12613_ (.A1(_09385_),
    .A2(_09273_),
    .A3(net2389),
    .B1(_09401_),
    .X(_01887_));
 sky130_fd_sc_hd__nor2_1 _12614_ (.A(_09216_),
    .B(_09386_),
    .Y(_09402_));
 sky130_fd_sc_hd__a31o_1 _12615_ (.A1(_09303_),
    .A2(net1695),
    .A3(_09385_),
    .B1(_09402_),
    .X(_01872_));
 sky130_fd_sc_hd__nand2_1 _12616_ (.A(_09391_),
    .B(net3644),
    .Y(_09403_));
 sky130_fd_sc_hd__a22o_1 _12617_ (.A1(_09390_),
    .A2(_09219_),
    .B1(_09384_),
    .B2(_09403_),
    .X(_09404_));
 sky130_fd_sc_hd__inv_2 _12618_ (.A(_09404_),
    .Y(_01873_));
 sky130_fd_sc_hd__nand2_1 _12619_ (.A(_09391_),
    .B(net4136),
    .Y(_09405_));
 sky130_fd_sc_hd__a22o_1 _12620_ (.A1(_09390_),
    .A2(_09332_),
    .B1(_09384_),
    .B2(_09405_),
    .X(_09406_));
 sky130_fd_sc_hd__inv_2 _12621_ (.A(_09406_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _12622_ (.A(_09230_),
    .B(_09386_),
    .Y(_09407_));
 sky130_fd_sc_hd__a31o_1 _12623_ (.A1(_09303_),
    .A2(net1357),
    .A3(_09385_),
    .B1(_09407_),
    .X(_01875_));
 sky130_fd_sc_hd__nor2_1 _12624_ (.A(_09233_),
    .B(_09386_),
    .Y(_09408_));
 sky130_fd_sc_hd__a31o_1 _12625_ (.A1(_09303_),
    .A2(net1624),
    .A3(_09386_),
    .B1(_09408_),
    .X(_01876_));
 sky130_fd_sc_hd__nor2_1 _12626_ (.A(_09236_),
    .B(_09386_),
    .Y(_09409_));
 sky130_fd_sc_hd__a31o_1 _12627_ (.A1(_09303_),
    .A2(net1469),
    .A3(_09386_),
    .B1(_09409_),
    .X(_01877_));
 sky130_fd_sc_hd__nand2_1 _12628_ (.A(_09391_),
    .B(net3612),
    .Y(_09410_));
 sky130_fd_sc_hd__a22o_1 _12629_ (.A1(_09390_),
    .A2(_09239_),
    .B1(_09384_),
    .B2(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__inv_2 _12630_ (.A(_09411_),
    .Y(_01878_));
 sky130_fd_sc_hd__buf_4 _12631_ (.A(_09302_),
    .X(_09412_));
 sky130_fd_sc_hd__nor2_1 _12632_ (.A(_09243_),
    .B(_09386_),
    .Y(_09413_));
 sky130_fd_sc_hd__a31o_1 _12633_ (.A1(_09412_),
    .A2(net1047),
    .A3(_09386_),
    .B1(_09413_),
    .X(_01879_));
 sky130_fd_sc_hd__nor2_8 _12634_ (.A(net81),
    .B(_09199_),
    .Y(_09414_));
 sky130_fd_sc_hd__buf_12 _12635_ (.A(net137),
    .X(_09415_));
 sky130_fd_sc_hd__nand2_1 _12636_ (.A(_09391_),
    .B(net3896),
    .Y(_09416_));
 sky130_fd_sc_hd__a22o_1 _12637_ (.A1(_09390_),
    .A2(_09415_),
    .B1(_09384_),
    .B2(_09416_),
    .X(_09417_));
 sky130_fd_sc_hd__inv_2 _12638_ (.A(_09417_),
    .Y(_01856_));
 sky130_fd_sc_hd__and3_1 _12639_ (.A(_09381_),
    .B(_09345_),
    .C(_09360_),
    .X(_09418_));
 sky130_fd_sc_hd__a31o_1 _12640_ (.A1(_09385_),
    .A2(_09273_),
    .A3(net2412),
    .B1(_09418_),
    .X(_01857_));
 sky130_fd_sc_hd__nor2_1 _12641_ (.A(_09253_),
    .B(_09386_),
    .Y(_09419_));
 sky130_fd_sc_hd__a31o_1 _12642_ (.A1(_09412_),
    .A2(net1019),
    .A3(_09386_),
    .B1(_09419_),
    .X(_01858_));
 sky130_fd_sc_hd__and3_1 _12643_ (.A(_09381_),
    .B(_09351_),
    .C(_09360_),
    .X(_09420_));
 sky130_fd_sc_hd__a31o_1 _12644_ (.A1(_09385_),
    .A2(_09273_),
    .A3(net2383),
    .B1(_09420_),
    .X(_01859_));
 sky130_fd_sc_hd__nor2_1 _12645_ (.A(_09260_),
    .B(_09386_),
    .Y(_09421_));
 sky130_fd_sc_hd__a31o_1 _12646_ (.A1(_09412_),
    .A2(net1313),
    .A3(_09386_),
    .B1(_09421_),
    .X(_01860_));
 sky130_fd_sc_hd__nand2_1 _12647_ (.A(_09391_),
    .B(net3746),
    .Y(_09422_));
 sky130_fd_sc_hd__a22o_1 _12648_ (.A1(_09390_),
    .A2(_09263_),
    .B1(_09384_),
    .B2(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__inv_2 _12649_ (.A(_09423_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_8 _12650_ (.A(net55),
    .B(_09199_),
    .Y(_09424_));
 sky130_fd_sc_hd__buf_12 _12651_ (.A(_09424_),
    .X(_09425_));
 sky130_fd_sc_hd__nand2_1 _12652_ (.A(_09391_),
    .B(net3194),
    .Y(_09426_));
 sky130_fd_sc_hd__a22o_1 _12653_ (.A1(_09390_),
    .A2(_09425_),
    .B1(_09384_),
    .B2(_09426_),
    .X(_09427_));
 sky130_fd_sc_hd__inv_2 _12654_ (.A(_09427_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_1 _12655_ (.A(_09391_),
    .B(net3414),
    .Y(_09428_));
 sky130_fd_sc_hd__a22o_1 _12656_ (.A1(_09390_),
    .A2(_09269_),
    .B1(_09384_),
    .B2(_09428_),
    .X(_09429_));
 sky130_fd_sc_hd__inv_2 _12657_ (.A(_09429_),
    .Y(_01863_));
 sky130_fd_sc_hd__and3_1 _12658_ (.A(_09381_),
    .B(_09274_),
    .C(_09360_),
    .X(_09430_));
 sky130_fd_sc_hd__a31o_1 _12659_ (.A1(_09385_),
    .A2(_09273_),
    .A3(net2342),
    .B1(_09430_),
    .X(_01848_));
 sky130_fd_sc_hd__nor2_1 _12660_ (.A(_09277_),
    .B(_09384_),
    .Y(_09431_));
 sky130_fd_sc_hd__a31o_1 _12661_ (.A1(_09412_),
    .A2(net1305),
    .A3(_09386_),
    .B1(_09431_),
    .X(_01849_));
 sky130_fd_sc_hd__clkbuf_8 _12662_ (.A(_09223_),
    .X(_09432_));
 sky130_fd_sc_hd__and3_1 _12663_ (.A(_09381_),
    .B(_09369_),
    .C(_09360_),
    .X(_09433_));
 sky130_fd_sc_hd__a31o_1 _12664_ (.A1(_09385_),
    .A2(_09432_),
    .A3(net2351),
    .B1(_09433_),
    .X(_01850_));
 sky130_fd_sc_hd__nand2_1 _12665_ (.A(_09391_),
    .B(net3074),
    .Y(_09434_));
 sky130_fd_sc_hd__a22o_1 _12666_ (.A1(_09390_),
    .A2(_09284_),
    .B1(_09384_),
    .B2(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__inv_2 _12667_ (.A(_09435_),
    .Y(_01851_));
 sky130_fd_sc_hd__and3_1 _12668_ (.A(_09381_),
    .B(_09373_),
    .C(_09360_),
    .X(_09436_));
 sky130_fd_sc_hd__a31o_1 _12669_ (.A1(_09385_),
    .A2(_09432_),
    .A3(net1605),
    .B1(_09436_),
    .X(_01852_));
 sky130_fd_sc_hd__nand2_1 _12670_ (.A(_09376_),
    .B(net3777),
    .Y(_09437_));
 sky130_fd_sc_hd__o2bb2a_1 _12671_ (.A1_N(_09437_),
    .A2_N(_09385_),
    .B1(_09294_),
    .B2(_09382_),
    .X(_01853_));
 sky130_fd_sc_hd__nand2_1 _12672_ (.A(_09376_),
    .B(net3674),
    .Y(_09438_));
 sky130_fd_sc_hd__o2bb2a_1 _12673_ (.A1_N(_09438_),
    .A2_N(_09385_),
    .B1(_09298_),
    .B2(_09382_),
    .X(_01854_));
 sky130_fd_sc_hd__nand2_1 _12674_ (.A(_09376_),
    .B(net3682),
    .Y(_09439_));
 sky130_fd_sc_hd__nor2_8 _12675_ (.A(net80),
    .B(_08727_),
    .Y(_09440_));
 sky130_fd_sc_hd__inv_6 _12676_ (.A(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__buf_8 _12677_ (.A(_09441_),
    .X(_09442_));
 sky130_fd_sc_hd__o2bb2a_1 _12678_ (.A1_N(_09439_),
    .A2_N(_09385_),
    .B1(_09382_),
    .B2(_09442_),
    .X(_01855_));
 sky130_fd_sc_hd__inv_2 _12679_ (.A(\line_cache_idx[8] ),
    .Y(_09443_));
 sky130_fd_sc_hd__buf_8 _12680_ (.A(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__nor2_2 _12681_ (.A(net2781),
    .B(net4297),
    .Y(_09445_));
 sky130_fd_sc_hd__nand2_1 _12682_ (.A(_09171_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__nor2_2 _12683_ (.A(_09444_),
    .B(_09446_),
    .Y(_09447_));
 sky130_fd_sc_hd__inv_2 _12684_ (.A(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__nor2_4 _12685_ (.A(_09190_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__nor2_2 _12686_ (.A(net66),
    .B(_09192_),
    .Y(_09450_));
 sky130_fd_sc_hd__buf_12 _12687_ (.A(_09450_),
    .X(_09451_));
 sky130_fd_sc_hd__nor2_1 _12688_ (.A(_09166_),
    .B(_09448_),
    .Y(_09452_));
 sky130_fd_sc_hd__inv_2 _12689_ (.A(_09452_),
    .Y(_09453_));
 sky130_fd_sc_hd__buf_4 _12690_ (.A(_09453_),
    .X(_09454_));
 sky130_fd_sc_hd__nand2_1 _12691_ (.A(_09391_),
    .B(net3303),
    .Y(_09455_));
 sky130_fd_sc_hd__a22o_1 _12692_ (.A1(_09449_),
    .A2(_09451_),
    .B1(_09454_),
    .B2(_09455_),
    .X(_09456_));
 sky130_fd_sc_hd__inv_2 _12693_ (.A(_09456_),
    .Y(_01840_));
 sky130_fd_sc_hd__buf_4 _12694_ (.A(_09453_),
    .X(_09457_));
 sky130_fd_sc_hd__nor2_1 _12695_ (.A(_09185_),
    .B(_09454_),
    .Y(_09458_));
 sky130_fd_sc_hd__a31o_1 _12696_ (.A1(_09412_),
    .A2(net1005),
    .A3(_09457_),
    .B1(_09458_),
    .X(_01841_));
 sky130_fd_sc_hd__nor2_8 _12697_ (.A(net68),
    .B(_09192_),
    .Y(_09459_));
 sky130_fd_sc_hd__buf_12 _12698_ (.A(_09459_),
    .X(_09460_));
 sky130_fd_sc_hd__nand2_1 _12699_ (.A(_09391_),
    .B(net3138),
    .Y(_09461_));
 sky130_fd_sc_hd__a22o_1 _12700_ (.A1(_09449_),
    .A2(_09460_),
    .B1(_09454_),
    .B2(_09461_),
    .X(_09462_));
 sky130_fd_sc_hd__inv_2 _12701_ (.A(_09462_),
    .Y(_01842_));
 sky130_fd_sc_hd__buf_8 _12702_ (.A(net69),
    .X(_09463_));
 sky130_fd_sc_hd__and3_1 _12703_ (.A(_09447_),
    .B(_09463_),
    .C(_09360_),
    .X(_09464_));
 sky130_fd_sc_hd__a31o_1 _12704_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net1037),
    .B1(_09464_),
    .X(_01843_));
 sky130_fd_sc_hd__and3_1 _12705_ (.A(_09447_),
    .B(_09321_),
    .C(_09360_),
    .X(_09465_));
 sky130_fd_sc_hd__a31o_1 _12706_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net729),
    .B1(_09465_),
    .X(_01844_));
 sky130_fd_sc_hd__and3_1 _12707_ (.A(_09447_),
    .B(_09395_),
    .C(_09360_),
    .X(_09466_));
 sky130_fd_sc_hd__a31o_1 _12708_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net1741),
    .B1(_09466_),
    .X(_01845_));
 sky130_fd_sc_hd__nor2_1 _12709_ (.A(_09209_),
    .B(_09454_),
    .Y(_09467_));
 sky130_fd_sc_hd__a31o_1 _12710_ (.A1(_09412_),
    .A2(net2168),
    .A3(_09457_),
    .B1(_09467_),
    .X(_01846_));
 sky130_fd_sc_hd__nand2_1 _12711_ (.A(_09391_),
    .B(net3192),
    .Y(_09468_));
 sky130_fd_sc_hd__a22o_1 _12712_ (.A1(_09449_),
    .A2(_09212_),
    .B1(_09454_),
    .B2(_09468_),
    .X(_09469_));
 sky130_fd_sc_hd__inv_2 _12713_ (.A(_09469_),
    .Y(_01847_));
 sky130_fd_sc_hd__nor2_1 _12714_ (.A(_09216_),
    .B(_09454_),
    .Y(_09470_));
 sky130_fd_sc_hd__a31o_1 _12715_ (.A1(_09412_),
    .A2(net971),
    .A3(_09457_),
    .B1(_09470_),
    .X(_01832_));
 sky130_fd_sc_hd__nand2_1 _12716_ (.A(_09391_),
    .B(net3528),
    .Y(_09471_));
 sky130_fd_sc_hd__a22o_1 _12717_ (.A1(_09449_),
    .A2(_09219_),
    .B1(_09454_),
    .B2(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__inv_2 _12718_ (.A(_09472_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _12719_ (.A(_09391_),
    .B(net3369),
    .Y(_09473_));
 sky130_fd_sc_hd__a22o_1 _12720_ (.A1(_09449_),
    .A2(_09332_),
    .B1(_09453_),
    .B2(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__inv_2 _12721_ (.A(_09474_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _12722_ (.A(_09230_),
    .B(_09454_),
    .Y(_09475_));
 sky130_fd_sc_hd__a31o_1 _12723_ (.A1(_09412_),
    .A2(net1575),
    .A3(_09457_),
    .B1(_09475_),
    .X(_01835_));
 sky130_fd_sc_hd__nor2_1 _12724_ (.A(_09233_),
    .B(_09454_),
    .Y(_09476_));
 sky130_fd_sc_hd__a31o_1 _12725_ (.A1(_09412_),
    .A2(net739),
    .A3(_09457_),
    .B1(_09476_),
    .X(_01836_));
 sky130_fd_sc_hd__nor2_1 _12726_ (.A(_09236_),
    .B(_09454_),
    .Y(_09477_));
 sky130_fd_sc_hd__a31o_1 _12727_ (.A1(_09412_),
    .A2(net1546),
    .A3(_09457_),
    .B1(_09477_),
    .X(_01837_));
 sky130_fd_sc_hd__and3_1 _12728_ (.A(_09447_),
    .B(_09341_),
    .C(_09360_),
    .X(_09478_));
 sky130_fd_sc_hd__a31o_1 _12729_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net1874),
    .B1(_09478_),
    .X(_01838_));
 sky130_fd_sc_hd__nor2_1 _12730_ (.A(_09243_),
    .B(_09454_),
    .Y(_09479_));
 sky130_fd_sc_hd__a31o_1 _12731_ (.A1(_09412_),
    .A2(net1403),
    .A3(_09454_),
    .B1(_09479_),
    .X(_01839_));
 sky130_fd_sc_hd__nand2_1 _12732_ (.A(_09391_),
    .B(net3311),
    .Y(_09480_));
 sky130_fd_sc_hd__a22o_1 _12733_ (.A1(_09449_),
    .A2(_09415_),
    .B1(_09453_),
    .B2(_09480_),
    .X(_09481_));
 sky130_fd_sc_hd__inv_2 _12734_ (.A(_09481_),
    .Y(_01824_));
 sky130_fd_sc_hd__buf_4 _12735_ (.A(_09359_),
    .X(_09482_));
 sky130_fd_sc_hd__and3_1 _12736_ (.A(_09447_),
    .B(_09345_),
    .C(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__a31o_1 _12737_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net2418),
    .B1(_09483_),
    .X(_01825_));
 sky130_fd_sc_hd__clkbuf_8 _12738_ (.A(_08800_),
    .X(_09484_));
 sky130_fd_sc_hd__nand2_1 _12739_ (.A(_09484_),
    .B(net3012),
    .Y(_09485_));
 sky130_fd_sc_hd__a22o_1 _12740_ (.A1(_09449_),
    .A2(_09348_),
    .B1(_09453_),
    .B2(_09485_),
    .X(_09486_));
 sky130_fd_sc_hd__inv_2 _12741_ (.A(_09486_),
    .Y(_01826_));
 sky130_fd_sc_hd__and3_1 _12742_ (.A(_09447_),
    .B(_09351_),
    .C(_09482_),
    .X(_09487_));
 sky130_fd_sc_hd__a31o_1 _12743_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net2534),
    .B1(_09487_),
    .X(_01827_));
 sky130_fd_sc_hd__nor2_1 _12744_ (.A(_09260_),
    .B(_09454_),
    .Y(_09488_));
 sky130_fd_sc_hd__a31o_1 _12745_ (.A1(_09412_),
    .A2(net2052),
    .A3(_09454_),
    .B1(_09488_),
    .X(_01828_));
 sky130_fd_sc_hd__nand2_1 _12746_ (.A(_09484_),
    .B(net3180),
    .Y(_09489_));
 sky130_fd_sc_hd__a22o_1 _12747_ (.A1(_09449_),
    .A2(_09263_),
    .B1(_09453_),
    .B2(_09489_),
    .X(_09490_));
 sky130_fd_sc_hd__inv_2 _12748_ (.A(_09490_),
    .Y(_01829_));
 sky130_fd_sc_hd__and3_1 _12749_ (.A(_09447_),
    .B(_09266_),
    .C(_09482_),
    .X(_09491_));
 sky130_fd_sc_hd__a31o_1 _12750_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net2186),
    .B1(_09491_),
    .X(_01830_));
 sky130_fd_sc_hd__nand2_1 _12751_ (.A(_09484_),
    .B(net3111),
    .Y(_09492_));
 sky130_fd_sc_hd__a22o_1 _12752_ (.A1(_09449_),
    .A2(_09269_),
    .B1(_09453_),
    .B2(_09492_),
    .X(_09493_));
 sky130_fd_sc_hd__inv_2 _12753_ (.A(_09493_),
    .Y(_01831_));
 sky130_fd_sc_hd__nor2_4 _12754_ (.A(net50),
    .B(_09192_),
    .Y(_09494_));
 sky130_fd_sc_hd__buf_12 _12755_ (.A(net141),
    .X(_09495_));
 sky130_fd_sc_hd__nand2_1 _12756_ (.A(_09484_),
    .B(net2817),
    .Y(_09496_));
 sky130_fd_sc_hd__a22o_1 _12757_ (.A1(_09449_),
    .A2(_09495_),
    .B1(_09453_),
    .B2(_09496_),
    .X(_09497_));
 sky130_fd_sc_hd__inv_2 _12758_ (.A(_09497_),
    .Y(_01816_));
 sky130_fd_sc_hd__nor2_1 _12759_ (.A(_09277_),
    .B(_09454_),
    .Y(_09498_));
 sky130_fd_sc_hd__a31o_1 _12760_ (.A1(_09412_),
    .A2(net1337),
    .A3(_09454_),
    .B1(_09498_),
    .X(_01817_));
 sky130_fd_sc_hd__and3_1 _12761_ (.A(_09447_),
    .B(_09369_),
    .C(_09482_),
    .X(_09499_));
 sky130_fd_sc_hd__a31o_1 _12762_ (.A1(_09457_),
    .A2(_09432_),
    .A3(net1971),
    .B1(_09499_),
    .X(_01818_));
 sky130_fd_sc_hd__nand2_1 _12763_ (.A(_09484_),
    .B(net3134),
    .Y(_09500_));
 sky130_fd_sc_hd__a22o_1 _12764_ (.A1(_09449_),
    .A2(_09284_),
    .B1(_09453_),
    .B2(_09500_),
    .X(_09501_));
 sky130_fd_sc_hd__inv_2 _12765_ (.A(_09501_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _12766_ (.A(_09484_),
    .B(net2951),
    .Y(_09502_));
 sky130_fd_sc_hd__a22o_1 _12767_ (.A1(_09449_),
    .A2(_09288_),
    .B1(_09453_),
    .B2(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__inv_2 _12768_ (.A(_09503_),
    .Y(_01820_));
 sky130_fd_sc_hd__nor2_8 _12769_ (.A(net78),
    .B(_09193_),
    .Y(_09504_));
 sky130_fd_sc_hd__nand2_1 _12770_ (.A(_09484_),
    .B(net3435),
    .Y(_09505_));
 sky130_fd_sc_hd__a22o_1 _12771_ (.A1(_09449_),
    .A2(_09504_),
    .B1(_09453_),
    .B2(_09505_),
    .X(_09506_));
 sky130_fd_sc_hd__inv_2 _12772_ (.A(_09506_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _12773_ (.A(_09376_),
    .B(net3670),
    .Y(_09507_));
 sky130_fd_sc_hd__o2bb2a_1 _12774_ (.A1_N(_09507_),
    .A2_N(_09457_),
    .B1(_09298_),
    .B2(_09448_),
    .X(_01822_));
 sky130_fd_sc_hd__nand2_1 _12775_ (.A(_09376_),
    .B(net3815),
    .Y(_09508_));
 sky130_fd_sc_hd__o2bb2a_1 _12776_ (.A1_N(_09508_),
    .A2_N(_09457_),
    .B1(_09442_),
    .B2(_09448_),
    .X(_01823_));
 sky130_fd_sc_hd__nor2_8 _12777_ (.A(net3791),
    .B(_08758_),
    .Y(_09509_));
 sky130_fd_sc_hd__nand2_1 _12778_ (.A(_09509_),
    .B(_09169_),
    .Y(_09510_));
 sky130_fd_sc_hd__inv_2 _12779_ (.A(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_1 _12780_ (.A(_09511_),
    .B(_09173_),
    .Y(_09512_));
 sky130_fd_sc_hd__nor2_4 _12781_ (.A(_09444_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__inv_2 _12782_ (.A(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__nor2_1 _12783_ (.A(_08727_),
    .B(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__clkinv_4 _12784_ (.A(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__buf_4 _12785_ (.A(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__buf_4 _12786_ (.A(_09516_),
    .X(_09518_));
 sky130_fd_sc_hd__nor2_1 _12787_ (.A(_09181_),
    .B(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__a31o_1 _12788_ (.A1(_09412_),
    .A2(net865),
    .A3(_09517_),
    .B1(_09519_),
    .X(_01808_));
 sky130_fd_sc_hd__nor2_1 _12789_ (.A(_09185_),
    .B(_09518_),
    .Y(_09520_));
 sky130_fd_sc_hd__a31o_1 _12790_ (.A1(_09412_),
    .A2(net727),
    .A3(_09517_),
    .B1(_09520_),
    .X(_01809_));
 sky130_fd_sc_hd__nor2_1 _12791_ (.A(_09188_),
    .B(_09518_),
    .Y(_09521_));
 sky130_fd_sc_hd__a31o_1 _12792_ (.A1(_09412_),
    .A2(net1143),
    .A3(_09517_),
    .B1(_09521_),
    .X(_01810_));
 sky130_fd_sc_hd__nor2_4 _12793_ (.A(_08795_),
    .B(_09514_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand2_1 _12794_ (.A(_09484_),
    .B(net2961),
    .Y(_09523_));
 sky130_fd_sc_hd__a22o_1 _12795_ (.A1(_09522_),
    .A2(_09195_),
    .B1(_09518_),
    .B2(_09523_),
    .X(_09524_));
 sky130_fd_sc_hd__inv_2 _12796_ (.A(_09524_),
    .Y(_01811_));
 sky130_fd_sc_hd__and3_1 _12797_ (.A(_09513_),
    .B(_09321_),
    .C(_09482_),
    .X(_09525_));
 sky130_fd_sc_hd__a31o_1 _12798_ (.A1(_09517_),
    .A2(_09432_),
    .A3(net1839),
    .B1(_09525_),
    .X(_01812_));
 sky130_fd_sc_hd__and3_1 _12799_ (.A(_09513_),
    .B(_09395_),
    .C(_09482_),
    .X(_09526_));
 sky130_fd_sc_hd__a31o_1 _12800_ (.A1(_09517_),
    .A2(_09432_),
    .A3(net1947),
    .B1(_09526_),
    .X(_01813_));
 sky130_fd_sc_hd__buf_4 _12801_ (.A(_09302_),
    .X(_09527_));
 sky130_fd_sc_hd__nor2_1 _12802_ (.A(_09209_),
    .B(_09518_),
    .Y(_09528_));
 sky130_fd_sc_hd__a31o_1 _12803_ (.A1(_09527_),
    .A2(net985),
    .A3(_09517_),
    .B1(_09528_),
    .X(_01814_));
 sky130_fd_sc_hd__and3_1 _12804_ (.A(_09513_),
    .B(_09326_),
    .C(_09482_),
    .X(_09529_));
 sky130_fd_sc_hd__a31o_1 _12805_ (.A1(_09517_),
    .A2(_09432_),
    .A3(net1387),
    .B1(_09529_),
    .X(_01815_));
 sky130_fd_sc_hd__nor2_8 _12806_ (.A(net57),
    .B(_09199_),
    .Y(_09530_));
 sky130_fd_sc_hd__buf_12 _12807_ (.A(_09530_),
    .X(_09531_));
 sky130_fd_sc_hd__nand2_1 _12808_ (.A(_09484_),
    .B(net3880),
    .Y(_09532_));
 sky130_fd_sc_hd__a22o_1 _12809_ (.A1(_09522_),
    .A2(_09531_),
    .B1(_09516_),
    .B2(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__inv_2 _12810_ (.A(_09533_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2_1 _12811_ (.A(_09484_),
    .B(net2802),
    .Y(_09534_));
 sky130_fd_sc_hd__a22o_1 _12812_ (.A1(_09522_),
    .A2(_09219_),
    .B1(_09516_),
    .B2(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__inv_2 _12813_ (.A(_09535_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _12814_ (.A(_09484_),
    .B(net2814),
    .Y(_09536_));
 sky130_fd_sc_hd__a22o_1 _12815_ (.A1(_09522_),
    .A2(_09332_),
    .B1(_09516_),
    .B2(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__inv_2 _12816_ (.A(_09537_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _12817_ (.A(_09230_),
    .B(_09518_),
    .Y(_09538_));
 sky130_fd_sc_hd__a31o_1 _12818_ (.A1(_09527_),
    .A2(net1968),
    .A3(_09517_),
    .B1(_09538_),
    .X(_01803_));
 sky130_fd_sc_hd__nor2_1 _12819_ (.A(_09233_),
    .B(_09518_),
    .Y(_09539_));
 sky130_fd_sc_hd__a31o_1 _12820_ (.A1(_09527_),
    .A2(net553),
    .A3(_09518_),
    .B1(_09539_),
    .X(_01804_));
 sky130_fd_sc_hd__nand2_1 _12821_ (.A(_09484_),
    .B(net2877),
    .Y(_09540_));
 sky130_fd_sc_hd__a22o_1 _12822_ (.A1(_09522_),
    .A2(_09338_),
    .B1(_09516_),
    .B2(_09540_),
    .X(_09541_));
 sky130_fd_sc_hd__inv_2 _12823_ (.A(_09541_),
    .Y(_01805_));
 sky130_fd_sc_hd__and3_1 _12824_ (.A(_09513_),
    .B(_09341_),
    .C(_09482_),
    .X(_09542_));
 sky130_fd_sc_hd__a31o_1 _12825_ (.A1(_09517_),
    .A2(_09432_),
    .A3(net1021),
    .B1(_09542_),
    .X(_01806_));
 sky130_fd_sc_hd__nor2_1 _12826_ (.A(_09243_),
    .B(_09518_),
    .Y(_09543_));
 sky130_fd_sc_hd__a31o_1 _12827_ (.A1(_09527_),
    .A2(net563),
    .A3(_09518_),
    .B1(_09543_),
    .X(_01807_));
 sky130_fd_sc_hd__nor2_1 _12828_ (.A(_09246_),
    .B(_09518_),
    .Y(_09544_));
 sky130_fd_sc_hd__a31o_1 _12829_ (.A1(_09527_),
    .A2(net1961),
    .A3(_09518_),
    .B1(_09544_),
    .X(_01792_));
 sky130_fd_sc_hd__and3_1 _12830_ (.A(_09513_),
    .B(_09345_),
    .C(_09482_),
    .X(_09545_));
 sky130_fd_sc_hd__a31o_1 _12831_ (.A1(_09517_),
    .A2(_09432_),
    .A3(net2027),
    .B1(_09545_),
    .X(_01793_));
 sky130_fd_sc_hd__nor2_1 _12832_ (.A(_09253_),
    .B(_09518_),
    .Y(_09546_));
 sky130_fd_sc_hd__a31o_1 _12833_ (.A1(_09527_),
    .A2(net1259),
    .A3(_09518_),
    .B1(_09546_),
    .X(_01794_));
 sky130_fd_sc_hd__and3_1 _12834_ (.A(_09513_),
    .B(_09351_),
    .C(_09482_),
    .X(_09547_));
 sky130_fd_sc_hd__a31o_1 _12835_ (.A1(_09517_),
    .A2(_09432_),
    .A3(net2081),
    .B1(_09547_),
    .X(_01795_));
 sky130_fd_sc_hd__nand2_1 _12836_ (.A(_09484_),
    .B(net3425),
    .Y(_09548_));
 sky130_fd_sc_hd__a22o_1 _12837_ (.A1(_09522_),
    .A2(_09354_),
    .B1(_09516_),
    .B2(_09548_),
    .X(_09549_));
 sky130_fd_sc_hd__inv_2 _12838_ (.A(_09549_),
    .Y(_01796_));
 sky130_fd_sc_hd__nand2_1 _12839_ (.A(_09484_),
    .B(net3280),
    .Y(_09550_));
 sky130_fd_sc_hd__a22o_1 _12840_ (.A1(_09522_),
    .A2(_09263_),
    .B1(_09516_),
    .B2(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__inv_2 _12841_ (.A(_09551_),
    .Y(_01797_));
 sky130_fd_sc_hd__clkbuf_8 _12842_ (.A(_09223_),
    .X(_09552_));
 sky130_fd_sc_hd__and3_1 _12843_ (.A(_09513_),
    .B(_09266_),
    .C(_09482_),
    .X(_09553_));
 sky130_fd_sc_hd__a31o_1 _12844_ (.A1(_09517_),
    .A2(_09552_),
    .A3(net2448),
    .B1(_09553_),
    .X(_01798_));
 sky130_fd_sc_hd__nand2_1 _12845_ (.A(_09484_),
    .B(net3079),
    .Y(_09554_));
 sky130_fd_sc_hd__a22o_1 _12846_ (.A1(_09522_),
    .A2(_09269_),
    .B1(_09516_),
    .B2(_09554_),
    .X(_09555_));
 sky130_fd_sc_hd__inv_2 _12847_ (.A(_09555_),
    .Y(_01799_));
 sky130_fd_sc_hd__nand2_1 _12848_ (.A(_09484_),
    .B(net3378),
    .Y(_09556_));
 sky130_fd_sc_hd__a22o_1 _12849_ (.A1(_09522_),
    .A2(_09495_),
    .B1(_09516_),
    .B2(_09556_),
    .X(_09557_));
 sky130_fd_sc_hd__inv_2 _12850_ (.A(_09557_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _12851_ (.A(_09277_),
    .B(_09518_),
    .Y(_09558_));
 sky130_fd_sc_hd__a31o_1 _12852_ (.A1(_09527_),
    .A2(net2436),
    .A3(_09518_),
    .B1(_09558_),
    .X(_01785_));
 sky130_fd_sc_hd__and3_1 _12853_ (.A(_09513_),
    .B(_09369_),
    .C(_09482_),
    .X(_09559_));
 sky130_fd_sc_hd__a31o_1 _12854_ (.A1(_09517_),
    .A2(_09552_),
    .A3(net1942),
    .B1(_09559_),
    .X(_01786_));
 sky130_fd_sc_hd__buf_4 _12855_ (.A(_08800_),
    .X(_09560_));
 sky130_fd_sc_hd__nand2_1 _12856_ (.A(_09560_),
    .B(net3344),
    .Y(_09561_));
 sky130_fd_sc_hd__a22o_1 _12857_ (.A1(_09522_),
    .A2(_09284_),
    .B1(_09516_),
    .B2(_09561_),
    .X(_09562_));
 sky130_fd_sc_hd__inv_2 _12858_ (.A(_09562_),
    .Y(_01787_));
 sky130_fd_sc_hd__nand2_1 _12859_ (.A(_09560_),
    .B(net3543),
    .Y(_09563_));
 sky130_fd_sc_hd__a22o_1 _12860_ (.A1(_09522_),
    .A2(_09288_),
    .B1(_09516_),
    .B2(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__inv_2 _12861_ (.A(_09564_),
    .Y(_01788_));
 sky130_fd_sc_hd__nand2_1 _12862_ (.A(_09376_),
    .B(net3567),
    .Y(_09565_));
 sky130_fd_sc_hd__o2bb2a_1 _12863_ (.A1_N(_09565_),
    .A2_N(_09517_),
    .B1(_09294_),
    .B2(_09514_),
    .X(_01789_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(_09376_),
    .B(net3609),
    .Y(_09566_));
 sky130_fd_sc_hd__o2bb2a_1 _12865_ (.A1_N(_09566_),
    .A2_N(_09517_),
    .B1(_09298_),
    .B2(_09514_),
    .X(_01790_));
 sky130_fd_sc_hd__nand2_1 _12866_ (.A(_09376_),
    .B(net3778),
    .Y(_09567_));
 sky130_fd_sc_hd__o2bb2a_1 _12867_ (.A1_N(_09567_),
    .A2_N(_09517_),
    .B1(_09442_),
    .B2(_09514_),
    .X(_01791_));
 sky130_fd_sc_hd__and3_4 _12868_ (.A(_09511_),
    .B(\line_cache_idx[8] ),
    .C(_09305_),
    .X(_09568_));
 sky130_fd_sc_hd__inv_2 _12869_ (.A(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__nor2_1 _12870_ (.A(_09166_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__clkinv_4 _12871_ (.A(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__buf_4 _12872_ (.A(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__buf_4 _12873_ (.A(_09571_),
    .X(_09573_));
 sky130_fd_sc_hd__nor2_1 _12874_ (.A(_09181_),
    .B(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__a31o_1 _12875_ (.A1(_09527_),
    .A2(net787),
    .A3(_09572_),
    .B1(_09574_),
    .X(_01760_));
 sky130_fd_sc_hd__nor2_1 _12876_ (.A(_09185_),
    .B(_09573_),
    .Y(_09575_));
 sky130_fd_sc_hd__a31o_1 _12877_ (.A1(_09527_),
    .A2(net2360),
    .A3(_09572_),
    .B1(_09575_),
    .X(_01761_));
 sky130_fd_sc_hd__nor2_1 _12878_ (.A(_09188_),
    .B(_09573_),
    .Y(_09576_));
 sky130_fd_sc_hd__a31o_1 _12879_ (.A1(_09527_),
    .A2(net1207),
    .A3(_09572_),
    .B1(_09576_),
    .X(_01762_));
 sky130_fd_sc_hd__and3_1 _12880_ (.A(_09568_),
    .B(_09463_),
    .C(_09482_),
    .X(_09577_));
 sky130_fd_sc_hd__a31o_1 _12881_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net1702),
    .B1(_09577_),
    .X(_01763_));
 sky130_fd_sc_hd__and3_1 _12882_ (.A(_09568_),
    .B(_09321_),
    .C(_09482_),
    .X(_09578_));
 sky130_fd_sc_hd__a31o_1 _12883_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net1919),
    .B1(_09578_),
    .X(_01764_));
 sky130_fd_sc_hd__and3_1 _12884_ (.A(_09568_),
    .B(_09395_),
    .C(_09482_),
    .X(_09579_));
 sky130_fd_sc_hd__a31o_1 _12885_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net2299),
    .B1(_09579_),
    .X(_01765_));
 sky130_fd_sc_hd__nor2_1 _12886_ (.A(_09209_),
    .B(_09573_),
    .Y(_09580_));
 sky130_fd_sc_hd__a31o_1 _12887_ (.A1(_09527_),
    .A2(net1273),
    .A3(_09572_),
    .B1(_09580_),
    .X(_01766_));
 sky130_fd_sc_hd__and3_1 _12888_ (.A(_09568_),
    .B(_09326_),
    .C(_09482_),
    .X(_09581_));
 sky130_fd_sc_hd__a31o_1 _12889_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net2191),
    .B1(_09581_),
    .X(_01767_));
 sky130_fd_sc_hd__nor2_1 _12890_ (.A(_09216_),
    .B(_09573_),
    .Y(_09582_));
 sky130_fd_sc_hd__a31o_1 _12891_ (.A1(_09527_),
    .A2(net2158),
    .A3(_09573_),
    .B1(_09582_),
    .X(_01752_));
 sky130_fd_sc_hd__nor2_4 _12892_ (.A(_08795_),
    .B(_09569_),
    .Y(_09583_));
 sky130_fd_sc_hd__nand2_1 _12893_ (.A(_09560_),
    .B(net3573),
    .Y(_09584_));
 sky130_fd_sc_hd__a22o_1 _12894_ (.A1(_09583_),
    .A2(_09219_),
    .B1(_09571_),
    .B2(_09584_),
    .X(_09585_));
 sky130_fd_sc_hd__inv_2 _12895_ (.A(_09585_),
    .Y(_01753_));
 sky130_fd_sc_hd__nand2_1 _12896_ (.A(_09560_),
    .B(net3478),
    .Y(_09586_));
 sky130_fd_sc_hd__a22o_1 _12897_ (.A1(_09583_),
    .A2(_09332_),
    .B1(_09571_),
    .B2(_09586_),
    .X(_09587_));
 sky130_fd_sc_hd__inv_2 _12898_ (.A(_09587_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_8 _12899_ (.A(net60),
    .B(_09199_),
    .Y(_09588_));
 sky130_fd_sc_hd__buf_12 _12900_ (.A(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__nand2_1 _12901_ (.A(_09560_),
    .B(net3061),
    .Y(_09590_));
 sky130_fd_sc_hd__a22o_1 _12902_ (.A1(_09583_),
    .A2(_09589_),
    .B1(_09571_),
    .B2(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__inv_2 _12903_ (.A(_09591_),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_8 _12904_ (.A(net62),
    .B(_09199_),
    .Y(_09592_));
 sky130_fd_sc_hd__buf_12 _12905_ (.A(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__nand2_1 _12906_ (.A(_09560_),
    .B(net3212),
    .Y(_09594_));
 sky130_fd_sc_hd__a22o_1 _12907_ (.A1(_09583_),
    .A2(_09593_),
    .B1(_09571_),
    .B2(_09594_),
    .X(_09595_));
 sky130_fd_sc_hd__inv_2 _12908_ (.A(_09595_),
    .Y(_01756_));
 sky130_fd_sc_hd__nor2_1 _12909_ (.A(_09236_),
    .B(_09573_),
    .Y(_09596_));
 sky130_fd_sc_hd__a31o_1 _12910_ (.A1(_09527_),
    .A2(net1776),
    .A3(_09573_),
    .B1(_09596_),
    .X(_01757_));
 sky130_fd_sc_hd__nand2_1 _12911_ (.A(_09560_),
    .B(net3672),
    .Y(_09597_));
 sky130_fd_sc_hd__a22o_1 _12912_ (.A1(_09583_),
    .A2(_09239_),
    .B1(_09571_),
    .B2(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__inv_2 _12913_ (.A(_09598_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _12914_ (.A(_09243_),
    .B(_09573_),
    .Y(_09599_));
 sky130_fd_sc_hd__a31o_1 _12915_ (.A1(_09527_),
    .A2(net657),
    .A3(_09573_),
    .B1(_09599_),
    .X(_01759_));
 sky130_fd_sc_hd__nand2_1 _12916_ (.A(_09560_),
    .B(net3562),
    .Y(_09600_));
 sky130_fd_sc_hd__a22o_1 _12917_ (.A1(_09583_),
    .A2(_09415_),
    .B1(_09571_),
    .B2(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__inv_2 _12918_ (.A(_09601_),
    .Y(_01744_));
 sky130_fd_sc_hd__buf_4 _12919_ (.A(_09359_),
    .X(_09602_));
 sky130_fd_sc_hd__and3_1 _12920_ (.A(_09568_),
    .B(_09345_),
    .C(_09602_),
    .X(_09603_));
 sky130_fd_sc_hd__a31o_1 _12921_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net1848),
    .B1(_09603_),
    .X(_01745_));
 sky130_fd_sc_hd__nor2_1 _12922_ (.A(_09253_),
    .B(_09573_),
    .Y(_09604_));
 sky130_fd_sc_hd__a31o_1 _12923_ (.A1(_09527_),
    .A2(net1175),
    .A3(_09573_),
    .B1(_09604_),
    .X(_01746_));
 sky130_fd_sc_hd__and3_1 _12924_ (.A(_09568_),
    .B(_09351_),
    .C(_09602_),
    .X(_09605_));
 sky130_fd_sc_hd__a31o_1 _12925_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net1739),
    .B1(_09605_),
    .X(_01747_));
 sky130_fd_sc_hd__nor2_1 _12926_ (.A(_09260_),
    .B(_09573_),
    .Y(_09606_));
 sky130_fd_sc_hd__a31o_1 _12927_ (.A1(_09527_),
    .A2(net789),
    .A3(_09573_),
    .B1(_09606_),
    .X(_01748_));
 sky130_fd_sc_hd__nand2_1 _12928_ (.A(_09560_),
    .B(net3404),
    .Y(_09607_));
 sky130_fd_sc_hd__a22o_1 _12929_ (.A1(_09583_),
    .A2(_09263_),
    .B1(_09571_),
    .B2(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__inv_2 _12930_ (.A(_09608_),
    .Y(_01749_));
 sky130_fd_sc_hd__and3_1 _12931_ (.A(_09568_),
    .B(_09266_),
    .C(_09602_),
    .X(_09609_));
 sky130_fd_sc_hd__a31o_1 _12932_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net1737),
    .B1(_09609_),
    .X(_01750_));
 sky130_fd_sc_hd__nand2_1 _12933_ (.A(_09560_),
    .B(net3864),
    .Y(_09610_));
 sky130_fd_sc_hd__a22o_1 _12934_ (.A1(_09583_),
    .A2(_09269_),
    .B1(_09571_),
    .B2(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__inv_2 _12935_ (.A(_09611_),
    .Y(_01751_));
 sky130_fd_sc_hd__and3_1 _12936_ (.A(_09568_),
    .B(_09274_),
    .C(_09602_),
    .X(_09612_));
 sky130_fd_sc_hd__a31o_1 _12937_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net2210),
    .B1(_09612_),
    .X(_01736_));
 sky130_fd_sc_hd__clkbuf_8 _12938_ (.A(_09302_),
    .X(_09613_));
 sky130_fd_sc_hd__nor2_1 _12939_ (.A(_09277_),
    .B(_09571_),
    .Y(_09614_));
 sky130_fd_sc_hd__a31o_1 _12940_ (.A1(_09613_),
    .A2(net1649),
    .A3(_09573_),
    .B1(_09614_),
    .X(_01737_));
 sky130_fd_sc_hd__and3_1 _12941_ (.A(_09568_),
    .B(_09369_),
    .C(_09602_),
    .X(_09615_));
 sky130_fd_sc_hd__a31o_1 _12942_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net2287),
    .B1(_09615_),
    .X(_01738_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(_09560_),
    .B(net3355),
    .Y(_09616_));
 sky130_fd_sc_hd__a22o_1 _12944_ (.A1(_09583_),
    .A2(_09284_),
    .B1(_09571_),
    .B2(_09616_),
    .X(_09617_));
 sky130_fd_sc_hd__inv_2 _12945_ (.A(_09617_),
    .Y(_01739_));
 sky130_fd_sc_hd__and3_1 _12946_ (.A(_09568_),
    .B(_09373_),
    .C(_09602_),
    .X(_09618_));
 sky130_fd_sc_hd__a31o_1 _12947_ (.A1(_09572_),
    .A2(_09552_),
    .A3(net2234),
    .B1(_09618_),
    .X(_01740_));
 sky130_fd_sc_hd__nand2_1 _12948_ (.A(_09376_),
    .B(net3709),
    .Y(_09619_));
 sky130_fd_sc_hd__o2bb2a_1 _12949_ (.A1_N(_09619_),
    .A2_N(_09572_),
    .B1(_09294_),
    .B2(_09569_),
    .X(_01741_));
 sky130_fd_sc_hd__nand2_1 _12950_ (.A(_09376_),
    .B(net3808),
    .Y(_09620_));
 sky130_fd_sc_hd__o2bb2a_1 _12951_ (.A1_N(_09620_),
    .A2_N(_09572_),
    .B1(_09298_),
    .B2(_09569_),
    .X(_01742_));
 sky130_fd_sc_hd__nor2_1 _12952_ (.A(_09300_),
    .B(_09571_),
    .Y(_09621_));
 sky130_fd_sc_hd__a31o_1 _12953_ (.A1(_09613_),
    .A2(net2408),
    .A3(_09573_),
    .B1(_09621_),
    .X(_01743_));
 sky130_fd_sc_hd__and3_4 _12954_ (.A(_09511_),
    .B(_08736_),
    .C(_09380_),
    .X(_09622_));
 sky130_fd_sc_hd__inv_2 _12955_ (.A(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__nor2_4 _12956_ (.A(_09190_),
    .B(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__buf_12 _12957_ (.A(_08727_),
    .X(_09625_));
 sky130_fd_sc_hd__nor2_1 _12958_ (.A(_09625_),
    .B(_09623_),
    .Y(_09626_));
 sky130_fd_sc_hd__inv_2 _12959_ (.A(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__buf_4 _12960_ (.A(_09627_),
    .X(_09628_));
 sky130_fd_sc_hd__nand2_1 _12961_ (.A(_09560_),
    .B(net3200),
    .Y(_09629_));
 sky130_fd_sc_hd__a22o_1 _12962_ (.A1(_09624_),
    .A2(_09451_),
    .B1(_09628_),
    .B2(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__inv_2 _12963_ (.A(_09630_),
    .Y(_01728_));
 sky130_fd_sc_hd__buf_4 _12964_ (.A(_09627_),
    .X(_09631_));
 sky130_fd_sc_hd__nor2_1 _12965_ (.A(_09185_),
    .B(_09628_),
    .Y(_09632_));
 sky130_fd_sc_hd__a31o_1 _12966_ (.A1(_09613_),
    .A2(net847),
    .A3(_09631_),
    .B1(_09632_),
    .X(_01729_));
 sky130_fd_sc_hd__nor2_1 _12967_ (.A(_09188_),
    .B(_09628_),
    .Y(_09633_));
 sky130_fd_sc_hd__a31o_1 _12968_ (.A1(_09613_),
    .A2(net1674),
    .A3(_09631_),
    .B1(_09633_),
    .X(_01730_));
 sky130_fd_sc_hd__and3_1 _12969_ (.A(_09622_),
    .B(_09463_),
    .C(_09602_),
    .X(_09634_));
 sky130_fd_sc_hd__a31o_1 _12970_ (.A1(_09631_),
    .A2(_09552_),
    .A3(net1725),
    .B1(_09634_),
    .X(_01731_));
 sky130_fd_sc_hd__and3_1 _12971_ (.A(_09622_),
    .B(_09321_),
    .C(_09602_),
    .X(_09635_));
 sky130_fd_sc_hd__a31o_1 _12972_ (.A1(_09631_),
    .A2(_09552_),
    .A3(net2268),
    .B1(_09635_),
    .X(_01732_));
 sky130_fd_sc_hd__and3_1 _12973_ (.A(_09622_),
    .B(_09395_),
    .C(_09602_),
    .X(_09636_));
 sky130_fd_sc_hd__a31o_1 _12974_ (.A1(_09631_),
    .A2(_09552_),
    .A3(net2142),
    .B1(_09636_),
    .X(_01733_));
 sky130_fd_sc_hd__nand2_1 _12975_ (.A(_09560_),
    .B(net2908),
    .Y(_09637_));
 sky130_fd_sc_hd__a22o_1 _12976_ (.A1(_09624_),
    .A2(_09398_),
    .B1(_09628_),
    .B2(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__inv_2 _12977_ (.A(_09638_),
    .Y(_01734_));
 sky130_fd_sc_hd__and3_1 _12978_ (.A(_09622_),
    .B(_09326_),
    .C(_09602_),
    .X(_09639_));
 sky130_fd_sc_hd__a31o_1 _12979_ (.A1(_09631_),
    .A2(_09552_),
    .A3(net2289),
    .B1(_09639_),
    .X(_01735_));
 sky130_fd_sc_hd__nand2_1 _12980_ (.A(_09560_),
    .B(net3283),
    .Y(_09640_));
 sky130_fd_sc_hd__a22o_1 _12981_ (.A1(_09624_),
    .A2(_09531_),
    .B1(_09628_),
    .B2(_09640_),
    .X(_09641_));
 sky130_fd_sc_hd__inv_2 _12982_ (.A(_09641_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _12983_ (.A(_09560_),
    .B(net2942),
    .Y(_09642_));
 sky130_fd_sc_hd__a22o_1 _12984_ (.A1(_09624_),
    .A2(_09219_),
    .B1(_09628_),
    .B2(_09642_),
    .X(_09643_));
 sky130_fd_sc_hd__inv_2 _12985_ (.A(_09643_),
    .Y(_01721_));
 sky130_fd_sc_hd__nand2_1 _12986_ (.A(_09560_),
    .B(net2920),
    .Y(_09644_));
 sky130_fd_sc_hd__a22o_1 _12987_ (.A1(_09624_),
    .A2(_09332_),
    .B1(_09628_),
    .B2(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__inv_2 _12988_ (.A(_09645_),
    .Y(_01722_));
 sky130_fd_sc_hd__buf_4 _12989_ (.A(_08800_),
    .X(_09646_));
 sky130_fd_sc_hd__nand2_1 _12990_ (.A(_09646_),
    .B(net3714),
    .Y(_09647_));
 sky130_fd_sc_hd__a22o_1 _12991_ (.A1(_09624_),
    .A2(_09589_),
    .B1(_09627_),
    .B2(_09647_),
    .X(_09648_));
 sky130_fd_sc_hd__inv_2 _12992_ (.A(_09648_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_1 _12993_ (.A(_09646_),
    .B(net3126),
    .Y(_09649_));
 sky130_fd_sc_hd__a22o_1 _12994_ (.A1(_09624_),
    .A2(_09593_),
    .B1(_09627_),
    .B2(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__inv_2 _12995_ (.A(_09650_),
    .Y(_01724_));
 sky130_fd_sc_hd__nor2_1 _12996_ (.A(_09236_),
    .B(_09628_),
    .Y(_09651_));
 sky130_fd_sc_hd__a31o_1 _12997_ (.A1(_09613_),
    .A2(net999),
    .A3(_09631_),
    .B1(_09651_),
    .X(_01725_));
 sky130_fd_sc_hd__nand2_1 _12998_ (.A(_09646_),
    .B(net3614),
    .Y(_09652_));
 sky130_fd_sc_hd__a22o_1 _12999_ (.A1(_09624_),
    .A2(_09239_),
    .B1(_09627_),
    .B2(_09652_),
    .X(_09653_));
 sky130_fd_sc_hd__inv_2 _13000_ (.A(_09653_),
    .Y(_01726_));
 sky130_fd_sc_hd__nor2_1 _13001_ (.A(_09243_),
    .B(_09628_),
    .Y(_09654_));
 sky130_fd_sc_hd__a31o_1 _13002_ (.A1(_09613_),
    .A2(net1059),
    .A3(_09631_),
    .B1(_09654_),
    .X(_01727_));
 sky130_fd_sc_hd__nor2_1 _13003_ (.A(_09246_),
    .B(_09628_),
    .Y(_09655_));
 sky130_fd_sc_hd__a31o_1 _13004_ (.A1(_09613_),
    .A2(net1419),
    .A3(_09631_),
    .B1(_09655_),
    .X(_01712_));
 sky130_fd_sc_hd__clkbuf_8 _13005_ (.A(_09223_),
    .X(_09656_));
 sky130_fd_sc_hd__and3_1 _13006_ (.A(_09622_),
    .B(_09345_),
    .C(_09602_),
    .X(_09657_));
 sky130_fd_sc_hd__a31o_1 _13007_ (.A1(_09631_),
    .A2(_09656_),
    .A3(net2231),
    .B1(_09657_),
    .X(_01713_));
 sky130_fd_sc_hd__nor2_1 _13008_ (.A(_09253_),
    .B(_09628_),
    .Y(_09658_));
 sky130_fd_sc_hd__a31o_1 _13009_ (.A1(_09613_),
    .A2(net977),
    .A3(_09628_),
    .B1(_09658_),
    .X(_01714_));
 sky130_fd_sc_hd__and3_1 _13010_ (.A(_09622_),
    .B(_09351_),
    .C(_09602_),
    .X(_09659_));
 sky130_fd_sc_hd__a31o_1 _13011_ (.A1(_09631_),
    .A2(_09656_),
    .A3(net1655),
    .B1(_09659_),
    .X(_01715_));
 sky130_fd_sc_hd__nor2_1 _13012_ (.A(_09260_),
    .B(_09628_),
    .Y(_09660_));
 sky130_fd_sc_hd__a31o_1 _13013_ (.A1(_09613_),
    .A2(net2056),
    .A3(_09628_),
    .B1(_09660_),
    .X(_01716_));
 sky130_fd_sc_hd__nand2_1 _13014_ (.A(_09646_),
    .B(net3867),
    .Y(_09661_));
 sky130_fd_sc_hd__a22o_1 _13015_ (.A1(_09624_),
    .A2(_09263_),
    .B1(_09627_),
    .B2(_09661_),
    .X(_09662_));
 sky130_fd_sc_hd__inv_2 _13016_ (.A(_09662_),
    .Y(_01717_));
 sky130_fd_sc_hd__and3_1 _13017_ (.A(_09622_),
    .B(_09266_),
    .C(_09602_),
    .X(_09663_));
 sky130_fd_sc_hd__a31o_1 _13018_ (.A1(_09631_),
    .A2(_09656_),
    .A3(net2156),
    .B1(_09663_),
    .X(_01718_));
 sky130_fd_sc_hd__nand2_1 _13019_ (.A(_09646_),
    .B(net3776),
    .Y(_09664_));
 sky130_fd_sc_hd__a22o_1 _13020_ (.A1(_09624_),
    .A2(_09269_),
    .B1(_09627_),
    .B2(_09664_),
    .X(_09665_));
 sky130_fd_sc_hd__inv_2 _13021_ (.A(_09665_),
    .Y(_01719_));
 sky130_fd_sc_hd__and3_1 _13022_ (.A(_09622_),
    .B(_09274_),
    .C(_09602_),
    .X(_09666_));
 sky130_fd_sc_hd__a31o_1 _13023_ (.A1(_09631_),
    .A2(_09656_),
    .A3(net2315),
    .B1(_09666_),
    .X(_01704_));
 sky130_fd_sc_hd__nor2_1 _13024_ (.A(_09277_),
    .B(_09628_),
    .Y(_09667_));
 sky130_fd_sc_hd__a31o_1 _13025_ (.A1(_09613_),
    .A2(net571),
    .A3(_09628_),
    .B1(_09667_),
    .X(_01705_));
 sky130_fd_sc_hd__nand2_1 _13026_ (.A(_09646_),
    .B(net3564),
    .Y(_09668_));
 sky130_fd_sc_hd__a22o_1 _13027_ (.A1(_09624_),
    .A2(_09280_),
    .B1(_09627_),
    .B2(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__inv_2 _13028_ (.A(_09669_),
    .Y(_01706_));
 sky130_fd_sc_hd__nand2_1 _13029_ (.A(_09646_),
    .B(net3740),
    .Y(_09670_));
 sky130_fd_sc_hd__a22o_1 _13030_ (.A1(_09624_),
    .A2(_09284_),
    .B1(_09627_),
    .B2(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__inv_2 _13031_ (.A(_09671_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _13032_ (.A(_09646_),
    .B(net3665),
    .Y(_09672_));
 sky130_fd_sc_hd__a22o_1 _13033_ (.A1(_09624_),
    .A2(_09288_),
    .B1(_09627_),
    .B2(_09672_),
    .X(_09673_));
 sky130_fd_sc_hd__inv_2 _13034_ (.A(_09673_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand2_1 _13035_ (.A(_09376_),
    .B(net3675),
    .Y(_09674_));
 sky130_fd_sc_hd__o2bb2a_1 _13036_ (.A1_N(_09674_),
    .A2_N(_09631_),
    .B1(_09294_),
    .B2(_09623_),
    .X(_01709_));
 sky130_fd_sc_hd__nand2_1 _13037_ (.A(_09376_),
    .B(net3529),
    .Y(_09675_));
 sky130_fd_sc_hd__o2bb2a_1 _13038_ (.A1_N(_09675_),
    .A2_N(_09631_),
    .B1(_09298_),
    .B2(_09623_),
    .X(_01710_));
 sky130_fd_sc_hd__nand2_1 _13039_ (.A(_09376_),
    .B(net3794),
    .Y(_09676_));
 sky130_fd_sc_hd__o2bb2a_1 _13040_ (.A1_N(_09676_),
    .A2_N(_09631_),
    .B1(_09442_),
    .B2(_09623_),
    .X(_01711_));
 sky130_fd_sc_hd__nand2_2 _13041_ (.A(_09511_),
    .B(_09445_),
    .Y(_09677_));
 sky130_fd_sc_hd__nor2_4 _13042_ (.A(_09443_),
    .B(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__inv_2 _13043_ (.A(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__nor2_4 _13044_ (.A(_08795_),
    .B(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__nor2_1 _13045_ (.A(_09304_),
    .B(_09679_),
    .Y(_09681_));
 sky130_fd_sc_hd__inv_2 _13046_ (.A(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__buf_4 _13047_ (.A(_09682_),
    .X(_09683_));
 sky130_fd_sc_hd__nand2_1 _13048_ (.A(_09646_),
    .B(net3297),
    .Y(_09684_));
 sky130_fd_sc_hd__a22o_1 _13049_ (.A1(_09680_),
    .A2(_09451_),
    .B1(_09683_),
    .B2(_09684_),
    .X(_09685_));
 sky130_fd_sc_hd__inv_2 _13050_ (.A(_09685_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _13051_ (.A(_09646_),
    .B(net3328),
    .Y(_09686_));
 sky130_fd_sc_hd__a22o_1 _13052_ (.A1(_09680_),
    .A2(_09315_),
    .B1(_09683_),
    .B2(_09686_),
    .X(_09687_));
 sky130_fd_sc_hd__inv_2 _13053_ (.A(_09687_),
    .Y(_01697_));
 sky130_fd_sc_hd__nand2_1 _13054_ (.A(_09646_),
    .B(net3223),
    .Y(_09688_));
 sky130_fd_sc_hd__a22o_1 _13055_ (.A1(_09680_),
    .A2(_09460_),
    .B1(_09683_),
    .B2(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__inv_2 _13056_ (.A(_09689_),
    .Y(_01698_));
 sky130_fd_sc_hd__buf_4 _13057_ (.A(_09682_),
    .X(_09690_));
 sky130_fd_sc_hd__and3_1 _13058_ (.A(_09678_),
    .B(_09463_),
    .C(_09602_),
    .X(_09691_));
 sky130_fd_sc_hd__a31o_1 _13059_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net2159),
    .B1(_09691_),
    .X(_01699_));
 sky130_fd_sc_hd__nand2_1 _13060_ (.A(_09646_),
    .B(net3293),
    .Y(_09692_));
 sky130_fd_sc_hd__a22o_1 _13061_ (.A1(_09680_),
    .A2(_09201_),
    .B1(_09682_),
    .B2(_09692_),
    .X(_09693_));
 sky130_fd_sc_hd__inv_2 _13062_ (.A(_09693_),
    .Y(_01700_));
 sky130_fd_sc_hd__and3_1 _13063_ (.A(_09678_),
    .B(_09395_),
    .C(_09602_),
    .X(_09694_));
 sky130_fd_sc_hd__a31o_1 _13064_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net2040),
    .B1(_09694_),
    .X(_01701_));
 sky130_fd_sc_hd__nor2_1 _13065_ (.A(_09209_),
    .B(_09683_),
    .Y(_09695_));
 sky130_fd_sc_hd__a31o_1 _13066_ (.A1(_09613_),
    .A2(net2339),
    .A3(_09690_),
    .B1(_09695_),
    .X(_01702_));
 sky130_fd_sc_hd__buf_4 _13067_ (.A(_09359_),
    .X(_09696_));
 sky130_fd_sc_hd__and3_1 _13068_ (.A(_09678_),
    .B(_09326_),
    .C(_09696_),
    .X(_09697_));
 sky130_fd_sc_hd__a31o_1 _13069_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net1826),
    .B1(_09697_),
    .X(_01703_));
 sky130_fd_sc_hd__nor2_1 _13070_ (.A(_09216_),
    .B(_09683_),
    .Y(_09698_));
 sky130_fd_sc_hd__a31o_1 _13071_ (.A1(_09613_),
    .A2(net1483),
    .A3(_09690_),
    .B1(_09698_),
    .X(_01688_));
 sky130_fd_sc_hd__nand2_1 _13072_ (.A(_09646_),
    .B(net3734),
    .Y(_09699_));
 sky130_fd_sc_hd__a22o_1 _13073_ (.A1(_09680_),
    .A2(_09219_),
    .B1(_09682_),
    .B2(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__inv_2 _13074_ (.A(_09700_),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _13075_ (.A(_09646_),
    .B(net3484),
    .Y(_09701_));
 sky130_fd_sc_hd__a22o_1 _13076_ (.A1(_09680_),
    .A2(_09332_),
    .B1(_09682_),
    .B2(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__inv_2 _13077_ (.A(_09702_),
    .Y(_01690_));
 sky130_fd_sc_hd__nor2_1 _13078_ (.A(_09230_),
    .B(_09683_),
    .Y(_09703_));
 sky130_fd_sc_hd__a31o_1 _13079_ (.A1(_09613_),
    .A2(net1211),
    .A3(_09690_),
    .B1(_09703_),
    .X(_01691_));
 sky130_fd_sc_hd__nand2_1 _13080_ (.A(_09646_),
    .B(net3049),
    .Y(_09704_));
 sky130_fd_sc_hd__a22o_1 _13081_ (.A1(_09680_),
    .A2(_09593_),
    .B1(_09682_),
    .B2(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__inv_2 _13082_ (.A(_09705_),
    .Y(_01692_));
 sky130_fd_sc_hd__nor2_1 _13083_ (.A(_09236_),
    .B(_09683_),
    .Y(_09706_));
 sky130_fd_sc_hd__a31o_1 _13084_ (.A1(_09613_),
    .A2(net1003),
    .A3(_09690_),
    .B1(_09706_),
    .X(_01693_));
 sky130_fd_sc_hd__and3_1 _13085_ (.A(_09678_),
    .B(_09341_),
    .C(_09696_),
    .X(_09707_));
 sky130_fd_sc_hd__a31o_1 _13086_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net1696),
    .B1(_09707_),
    .X(_01694_));
 sky130_fd_sc_hd__nor2_1 _13087_ (.A(_09243_),
    .B(_09683_),
    .Y(_09708_));
 sky130_fd_sc_hd__a31o_1 _13088_ (.A1(_09613_),
    .A2(net2367),
    .A3(_09690_),
    .B1(_09708_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_1 _13089_ (.A(_09246_),
    .B(_09683_),
    .Y(_09709_));
 sky130_fd_sc_hd__a31o_1 _13090_ (.A1(_09613_),
    .A2(net2183),
    .A3(_09683_),
    .B1(_09709_),
    .X(_01672_));
 sky130_fd_sc_hd__nand2_1 _13091_ (.A(_09646_),
    .B(net3401),
    .Y(_09710_));
 sky130_fd_sc_hd__a22o_1 _13092_ (.A1(_09680_),
    .A2(_09249_),
    .B1(_09682_),
    .B2(_09710_),
    .X(_09711_));
 sky130_fd_sc_hd__inv_2 _13093_ (.A(_09711_),
    .Y(_01673_));
 sky130_fd_sc_hd__clkbuf_8 _13094_ (.A(_09302_),
    .X(_09712_));
 sky130_fd_sc_hd__nor2_1 _13095_ (.A(_09253_),
    .B(_09683_),
    .Y(_09713_));
 sky130_fd_sc_hd__a31o_1 _13096_ (.A1(_09712_),
    .A2(net1794),
    .A3(_09683_),
    .B1(_09713_),
    .X(_01674_));
 sky130_fd_sc_hd__and3_1 _13097_ (.A(_09678_),
    .B(_09351_),
    .C(_09696_),
    .X(_09714_));
 sky130_fd_sc_hd__a31o_1 _13098_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net1908),
    .B1(_09714_),
    .X(_01675_));
 sky130_fd_sc_hd__nor2_1 _13099_ (.A(_09260_),
    .B(_09683_),
    .Y(_09715_));
 sky130_fd_sc_hd__a31o_1 _13100_ (.A1(_09712_),
    .A2(net1473),
    .A3(_09683_),
    .B1(_09715_),
    .X(_01676_));
 sky130_fd_sc_hd__clkbuf_4 _13101_ (.A(_09222_),
    .X(_09716_));
 sky130_fd_sc_hd__clkbuf_8 _13102_ (.A(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__nand2_1 _13103_ (.A(_09717_),
    .B(net3857),
    .Y(_09718_));
 sky130_fd_sc_hd__a22o_1 _13104_ (.A1(_09680_),
    .A2(_09263_),
    .B1(_09682_),
    .B2(_09718_),
    .X(_09719_));
 sky130_fd_sc_hd__inv_2 _13105_ (.A(_09719_),
    .Y(_01677_));
 sky130_fd_sc_hd__and3_1 _13106_ (.A(_09678_),
    .B(_09266_),
    .C(_09696_),
    .X(_09720_));
 sky130_fd_sc_hd__a31o_1 _13107_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net1507),
    .B1(_09720_),
    .X(_01678_));
 sky130_fd_sc_hd__nand2_1 _13108_ (.A(_09717_),
    .B(net3803),
    .Y(_09721_));
 sky130_fd_sc_hd__a22o_1 _13109_ (.A1(_09680_),
    .A2(_09269_),
    .B1(_09682_),
    .B2(_09721_),
    .X(_09722_));
 sky130_fd_sc_hd__inv_2 _13110_ (.A(_09722_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _13111_ (.A(_09717_),
    .B(net3337),
    .Y(_09723_));
 sky130_fd_sc_hd__a22o_1 _13112_ (.A1(_09680_),
    .A2(_09495_),
    .B1(_09682_),
    .B2(_09723_),
    .X(_09724_));
 sky130_fd_sc_hd__inv_2 _13113_ (.A(_09724_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_1 _13114_ (.A(_09277_),
    .B(_09683_),
    .Y(_09725_));
 sky130_fd_sc_hd__a31o_1 _13115_ (.A1(_09712_),
    .A2(net861),
    .A3(_09683_),
    .B1(_09725_),
    .X(_01665_));
 sky130_fd_sc_hd__and3_1 _13116_ (.A(_09678_),
    .B(_09369_),
    .C(_09696_),
    .X(_09726_));
 sky130_fd_sc_hd__a31o_1 _13117_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net2474),
    .B1(_09726_),
    .X(_01666_));
 sky130_fd_sc_hd__nand2_1 _13118_ (.A(_09717_),
    .B(net3650),
    .Y(_09727_));
 sky130_fd_sc_hd__a22o_1 _13119_ (.A1(_09680_),
    .A2(_09284_),
    .B1(_09682_),
    .B2(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__inv_2 _13120_ (.A(_09728_),
    .Y(_01667_));
 sky130_fd_sc_hd__and3_1 _13121_ (.A(_09678_),
    .B(_09373_),
    .C(_09696_),
    .X(_09729_));
 sky130_fd_sc_hd__a31o_1 _13122_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net2294),
    .B1(_09729_),
    .X(_01668_));
 sky130_fd_sc_hd__buf_8 _13123_ (.A(net78),
    .X(_09730_));
 sky130_fd_sc_hd__and3_1 _13124_ (.A(_09678_),
    .B(_09730_),
    .C(_09696_),
    .X(_09731_));
 sky130_fd_sc_hd__a31o_1 _13125_ (.A1(_09690_),
    .A2(_09656_),
    .A3(net1769),
    .B1(_09731_),
    .X(_01669_));
 sky130_fd_sc_hd__nand2_1 _13126_ (.A(_09376_),
    .B(net3549),
    .Y(_09732_));
 sky130_fd_sc_hd__o2bb2a_1 _13127_ (.A1_N(_09732_),
    .A2_N(_09690_),
    .B1(_09298_),
    .B2(_09679_),
    .X(_01670_));
 sky130_fd_sc_hd__buf_6 _13128_ (.A(_09375_),
    .X(_09733_));
 sky130_fd_sc_hd__nand2_1 _13129_ (.A(_09733_),
    .B(net3580),
    .Y(_09734_));
 sky130_fd_sc_hd__o2bb2a_1 _13130_ (.A1_N(_09734_),
    .A2_N(_09690_),
    .B1(_09442_),
    .B2(_09679_),
    .X(_01671_));
 sky130_fd_sc_hd__nor2_8 _13131_ (.A(net2787),
    .B(_08756_),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_1 _13132_ (.A(_09735_),
    .B(_09169_),
    .Y(_09736_));
 sky130_fd_sc_hd__inv_2 _13133_ (.A(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__nand2_2 _13134_ (.A(_09737_),
    .B(_09173_),
    .Y(_09738_));
 sky130_fd_sc_hd__nor2_4 _13135_ (.A(_09444_),
    .B(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__inv_2 _13136_ (.A(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nor2_1 _13137_ (.A(_09166_),
    .B(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__clkinv_4 _13138_ (.A(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__buf_4 _13139_ (.A(_09742_),
    .X(_09743_));
 sky130_fd_sc_hd__buf_4 _13140_ (.A(_09742_),
    .X(_09744_));
 sky130_fd_sc_hd__nor2_1 _13141_ (.A(_09181_),
    .B(_09744_),
    .Y(_09745_));
 sky130_fd_sc_hd__a31o_1 _13142_ (.A1(_09712_),
    .A2(net2698),
    .A3(_09743_),
    .B1(_09745_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_4 _13143_ (.A(_08795_),
    .B(_09740_),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_1 _13144_ (.A(_09717_),
    .B(net4328),
    .Y(_09747_));
 sky130_fd_sc_hd__a22o_1 _13145_ (.A1(_09746_),
    .A2(_09315_),
    .B1(_09742_),
    .B2(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__inv_2 _13146_ (.A(_09748_),
    .Y(_01657_));
 sky130_fd_sc_hd__nor2_1 _13147_ (.A(_09188_),
    .B(_09744_),
    .Y(_09749_));
 sky130_fd_sc_hd__a31o_1 _13148_ (.A1(_09712_),
    .A2(net2721),
    .A3(_09743_),
    .B1(_09749_),
    .X(_01658_));
 sky130_fd_sc_hd__and3_1 _13149_ (.A(_09739_),
    .B(_09463_),
    .C(_09696_),
    .X(_09750_));
 sky130_fd_sc_hd__a31o_1 _13150_ (.A1(_09743_),
    .A2(_09656_),
    .A3(net2704),
    .B1(_09750_),
    .X(_01659_));
 sky130_fd_sc_hd__and3_1 _13151_ (.A(_09739_),
    .B(_09321_),
    .C(_09696_),
    .X(_09751_));
 sky130_fd_sc_hd__a31o_1 _13152_ (.A1(_09743_),
    .A2(_09656_),
    .A3(net2706),
    .B1(_09751_),
    .X(_01660_));
 sky130_fd_sc_hd__and3_1 _13153_ (.A(_09739_),
    .B(_09395_),
    .C(_09696_),
    .X(_09752_));
 sky130_fd_sc_hd__a31o_1 _13154_ (.A1(_09743_),
    .A2(_09656_),
    .A3(net2711),
    .B1(_09752_),
    .X(_01661_));
 sky130_fd_sc_hd__nand2_1 _13155_ (.A(_09717_),
    .B(net4326),
    .Y(_09753_));
 sky130_fd_sc_hd__a22o_1 _13156_ (.A1(_09746_),
    .A2(_09398_),
    .B1(_09742_),
    .B2(_09753_),
    .X(_09754_));
 sky130_fd_sc_hd__inv_2 _13157_ (.A(_09754_),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_1 _13158_ (.A(_09717_),
    .B(net4329),
    .Y(_09755_));
 sky130_fd_sc_hd__a22o_1 _13159_ (.A1(_09746_),
    .A2(_09212_),
    .B1(_09742_),
    .B2(_09755_),
    .X(_09756_));
 sky130_fd_sc_hd__inv_2 _13160_ (.A(_09756_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor2_1 _13161_ (.A(_09216_),
    .B(_09744_),
    .Y(_09757_));
 sky130_fd_sc_hd__a31o_1 _13162_ (.A1(_09712_),
    .A2(net2582),
    .A3(_09743_),
    .B1(_09757_),
    .X(_01648_));
 sky130_fd_sc_hd__nand2_1 _13163_ (.A(_09717_),
    .B(net3775),
    .Y(_09758_));
 sky130_fd_sc_hd__a22o_1 _13164_ (.A1(_09746_),
    .A2(_09219_),
    .B1(_09742_),
    .B2(_09758_),
    .X(_09759_));
 sky130_fd_sc_hd__inv_2 _13165_ (.A(_09759_),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_1 _13166_ (.A(_09717_),
    .B(net3584),
    .Y(_09760_));
 sky130_fd_sc_hd__a22o_1 _13167_ (.A1(_09746_),
    .A2(_09332_),
    .B1(_09742_),
    .B2(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__inv_2 _13168_ (.A(_09761_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _13169_ (.A(_09230_),
    .B(_09744_),
    .Y(_09762_));
 sky130_fd_sc_hd__a31o_1 _13170_ (.A1(_09712_),
    .A2(net2604),
    .A3(_09743_),
    .B1(_09762_),
    .X(_01651_));
 sky130_fd_sc_hd__nor2_1 _13171_ (.A(_09233_),
    .B(_09744_),
    .Y(_09763_));
 sky130_fd_sc_hd__a31o_1 _13172_ (.A1(_09712_),
    .A2(net2615),
    .A3(_09743_),
    .B1(_09763_),
    .X(_01652_));
 sky130_fd_sc_hd__nor2_1 _13173_ (.A(_09236_),
    .B(_09744_),
    .Y(_09764_));
 sky130_fd_sc_hd__a31o_1 _13174_ (.A1(_09712_),
    .A2(net2538),
    .A3(_09743_),
    .B1(_09764_),
    .X(_01653_));
 sky130_fd_sc_hd__nand2_1 _13175_ (.A(_09717_),
    .B(net3835),
    .Y(_09765_));
 sky130_fd_sc_hd__a22o_1 _13176_ (.A1(_09746_),
    .A2(_09239_),
    .B1(_09742_),
    .B2(_09765_),
    .X(_09766_));
 sky130_fd_sc_hd__inv_2 _13177_ (.A(_09766_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_8 _13178_ (.A(net65),
    .B(_09192_),
    .Y(_09767_));
 sky130_fd_sc_hd__buf_12 _13179_ (.A(_09767_),
    .X(_09768_));
 sky130_fd_sc_hd__nand2_1 _13180_ (.A(_09717_),
    .B(net4098),
    .Y(_09769_));
 sky130_fd_sc_hd__a22o_1 _13181_ (.A1(_09746_),
    .A2(_09768_),
    .B1(_09742_),
    .B2(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__inv_2 _13182_ (.A(_09770_),
    .Y(_01655_));
 sky130_fd_sc_hd__nor2_1 _13183_ (.A(_09246_),
    .B(_09744_),
    .Y(_09771_));
 sky130_fd_sc_hd__a31o_1 _13184_ (.A1(_09712_),
    .A2(net2539),
    .A3(_09744_),
    .B1(_09771_),
    .X(_01640_));
 sky130_fd_sc_hd__nand2_1 _13185_ (.A(_09717_),
    .B(net3677),
    .Y(_09772_));
 sky130_fd_sc_hd__a22o_1 _13186_ (.A1(_09746_),
    .A2(_09249_),
    .B1(_09742_),
    .B2(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__inv_2 _13187_ (.A(_09773_),
    .Y(_01641_));
 sky130_fd_sc_hd__nor2_1 _13188_ (.A(_09253_),
    .B(_09744_),
    .Y(_09774_));
 sky130_fd_sc_hd__a31o_1 _13189_ (.A1(_09712_),
    .A2(net2537),
    .A3(_09744_),
    .B1(_09774_),
    .X(_01642_));
 sky130_fd_sc_hd__buf_4 _13190_ (.A(_09223_),
    .X(_09775_));
 sky130_fd_sc_hd__and3_1 _13191_ (.A(_09739_),
    .B(_09351_),
    .C(_09696_),
    .X(_09776_));
 sky130_fd_sc_hd__a31o_1 _13192_ (.A1(_09743_),
    .A2(_09775_),
    .A3(net2171),
    .B1(_09776_),
    .X(_01643_));
 sky130_fd_sc_hd__nor2_1 _13193_ (.A(_09260_),
    .B(_09744_),
    .Y(_09777_));
 sky130_fd_sc_hd__a31o_1 _13194_ (.A1(_09712_),
    .A2(net2222),
    .A3(_09744_),
    .B1(_09777_),
    .X(_01644_));
 sky130_fd_sc_hd__nand2_1 _13195_ (.A(_09717_),
    .B(net3216),
    .Y(_09778_));
 sky130_fd_sc_hd__a22o_1 _13196_ (.A1(_09746_),
    .A2(_09263_),
    .B1(_09742_),
    .B2(_09778_),
    .X(_09779_));
 sky130_fd_sc_hd__inv_2 _13197_ (.A(_09779_),
    .Y(_01645_));
 sky130_fd_sc_hd__and3_1 _13198_ (.A(_09739_),
    .B(_09266_),
    .C(_09696_),
    .X(_09780_));
 sky130_fd_sc_hd__a31o_1 _13199_ (.A1(_09743_),
    .A2(_09775_),
    .A3(net1457),
    .B1(_09780_),
    .X(_01646_));
 sky130_fd_sc_hd__nand2_1 _13200_ (.A(_09717_),
    .B(net3125),
    .Y(_09781_));
 sky130_fd_sc_hd__a22o_1 _13201_ (.A1(_09746_),
    .A2(_09269_),
    .B1(_09742_),
    .B2(_09781_),
    .X(_09782_));
 sky130_fd_sc_hd__inv_2 _13202_ (.A(_09782_),
    .Y(_01647_));
 sky130_fd_sc_hd__and3_1 _13203_ (.A(_09739_),
    .B(_09274_),
    .C(_09696_),
    .X(_09783_));
 sky130_fd_sc_hd__a31o_1 _13204_ (.A1(_09743_),
    .A2(_09775_),
    .A3(net2301),
    .B1(_09783_),
    .X(_01632_));
 sky130_fd_sc_hd__nor2_1 _13205_ (.A(_09277_),
    .B(_09744_),
    .Y(_09784_));
 sky130_fd_sc_hd__a31o_1 _13206_ (.A1(_09712_),
    .A2(net2119),
    .A3(_09744_),
    .B1(_09784_),
    .X(_01633_));
 sky130_fd_sc_hd__and3_1 _13207_ (.A(_09739_),
    .B(_09369_),
    .C(_09696_),
    .X(_09785_));
 sky130_fd_sc_hd__a31o_1 _13208_ (.A1(_09743_),
    .A2(_09775_),
    .A3(net2619),
    .B1(_09785_),
    .X(_01634_));
 sky130_fd_sc_hd__nand2_1 _13209_ (.A(_09717_),
    .B(net3022),
    .Y(_09786_));
 sky130_fd_sc_hd__a22o_1 _13210_ (.A1(_09746_),
    .A2(_09284_),
    .B1(_09742_),
    .B2(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__inv_2 _13211_ (.A(_09787_),
    .Y(_01635_));
 sky130_fd_sc_hd__and3_1 _13212_ (.A(_09739_),
    .B(_09373_),
    .C(_09696_),
    .X(_09788_));
 sky130_fd_sc_hd__a31o_1 _13213_ (.A1(_09743_),
    .A2(_09775_),
    .A3(net1673),
    .B1(_09788_),
    .X(_01636_));
 sky130_fd_sc_hd__and3_1 _13214_ (.A(_09739_),
    .B(_09730_),
    .C(_09696_),
    .X(_09789_));
 sky130_fd_sc_hd__a31o_1 _13215_ (.A1(_09743_),
    .A2(_09775_),
    .A3(net1618),
    .B1(_09789_),
    .X(_01637_));
 sky130_fd_sc_hd__nand2_1 _13216_ (.A(_09733_),
    .B(net3610),
    .Y(_09790_));
 sky130_fd_sc_hd__o2bb2a_1 _13217_ (.A1_N(_09790_),
    .A2_N(_09743_),
    .B1(_09298_),
    .B2(_09740_),
    .X(_01638_));
 sky130_fd_sc_hd__nor2_1 _13218_ (.A(_09300_),
    .B(_09744_),
    .Y(_09791_));
 sky130_fd_sc_hd__a31o_1 _13219_ (.A1(_09712_),
    .A2(net1887),
    .A3(_09744_),
    .B1(_09791_),
    .X(_01639_));
 sky130_fd_sc_hd__and3_4 _13220_ (.A(_09737_),
    .B(_08736_),
    .C(_09305_),
    .X(_09792_));
 sky130_fd_sc_hd__inv_2 _13221_ (.A(_09792_),
    .Y(_09793_));
 sky130_fd_sc_hd__nor2_1 _13222_ (.A(_08794_),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__buf_4 _13223_ (.A(_09794_),
    .X(_09795_));
 sky130_fd_sc_hd__nor2_1 _13224_ (.A(_08728_),
    .B(_09793_),
    .Y(_09796_));
 sky130_fd_sc_hd__inv_2 _13225_ (.A(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__buf_4 _13226_ (.A(_09797_),
    .X(_09798_));
 sky130_fd_sc_hd__nand2_1 _13227_ (.A(_09717_),
    .B(net3313),
    .Y(_09799_));
 sky130_fd_sc_hd__a22o_1 _13228_ (.A1(_09795_),
    .A2(_09451_),
    .B1(_09798_),
    .B2(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__inv_2 _13229_ (.A(_09800_),
    .Y(_01624_));
 sky130_fd_sc_hd__buf_4 _13230_ (.A(_09716_),
    .X(_09801_));
 sky130_fd_sc_hd__nand2_1 _13231_ (.A(_09801_),
    .B(net3228),
    .Y(_09802_));
 sky130_fd_sc_hd__a22o_1 _13232_ (.A1(_09795_),
    .A2(_09315_),
    .B1(_09798_),
    .B2(_09802_),
    .X(_09803_));
 sky130_fd_sc_hd__inv_2 _13233_ (.A(_09803_),
    .Y(_01625_));
 sky130_fd_sc_hd__nand2_1 _13234_ (.A(_09801_),
    .B(net3190),
    .Y(_09804_));
 sky130_fd_sc_hd__a22o_1 _13235_ (.A1(_09795_),
    .A2(_09460_),
    .B1(_09798_),
    .B2(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__inv_2 _13236_ (.A(_09805_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _13237_ (.A(_09801_),
    .B(net3266),
    .Y(_09806_));
 sky130_fd_sc_hd__a22o_1 _13238_ (.A1(_09795_),
    .A2(_09195_),
    .B1(_09798_),
    .B2(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__inv_2 _13239_ (.A(_09807_),
    .Y(_01627_));
 sky130_fd_sc_hd__nand2_1 _13240_ (.A(_09801_),
    .B(net3315),
    .Y(_09808_));
 sky130_fd_sc_hd__a22o_1 _13241_ (.A1(_09795_),
    .A2(_09201_),
    .B1(_09798_),
    .B2(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__inv_2 _13242_ (.A(_09809_),
    .Y(_01628_));
 sky130_fd_sc_hd__nand2_1 _13243_ (.A(_09801_),
    .B(net3537),
    .Y(_09810_));
 sky130_fd_sc_hd__a22o_1 _13244_ (.A1(_09795_),
    .A2(_09205_),
    .B1(_09798_),
    .B2(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__inv_2 _13245_ (.A(_09811_),
    .Y(_01629_));
 sky130_fd_sc_hd__nand2_1 _13246_ (.A(_09801_),
    .B(net2901),
    .Y(_09812_));
 sky130_fd_sc_hd__a22o_1 _13247_ (.A1(_09795_),
    .A2(_09398_),
    .B1(_09798_),
    .B2(_09812_),
    .X(_09813_));
 sky130_fd_sc_hd__inv_2 _13248_ (.A(_09813_),
    .Y(_01630_));
 sky130_fd_sc_hd__nand2_1 _13249_ (.A(_09801_),
    .B(net3058),
    .Y(_09814_));
 sky130_fd_sc_hd__a22o_1 _13250_ (.A1(_09795_),
    .A2(_09212_),
    .B1(_09798_),
    .B2(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__inv_2 _13251_ (.A(_09815_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand2_1 _13252_ (.A(_09801_),
    .B(net3901),
    .Y(_09816_));
 sky130_fd_sc_hd__a22o_1 _13253_ (.A1(_09795_),
    .A2(_09531_),
    .B1(_09798_),
    .B2(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__inv_2 _13254_ (.A(_09817_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _13255_ (.A(_09801_),
    .B(net3122),
    .Y(_09818_));
 sky130_fd_sc_hd__a22o_1 _13256_ (.A1(_09795_),
    .A2(_09219_),
    .B1(_09798_),
    .B2(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__inv_2 _13257_ (.A(_09819_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand2_1 _13258_ (.A(_09801_),
    .B(net3103),
    .Y(_09820_));
 sky130_fd_sc_hd__a22o_1 _13259_ (.A1(_09795_),
    .A2(_09332_),
    .B1(_09798_),
    .B2(_09820_),
    .X(_09821_));
 sky130_fd_sc_hd__inv_2 _13260_ (.A(_09821_),
    .Y(_01618_));
 sky130_fd_sc_hd__buf_4 _13261_ (.A(_09797_),
    .X(_09822_));
 sky130_fd_sc_hd__nor2_1 _13262_ (.A(_09230_),
    .B(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__a31o_1 _13263_ (.A1(_09712_),
    .A2(net1261),
    .A3(_09822_),
    .B1(_09823_),
    .X(_01619_));
 sky130_fd_sc_hd__nand2_1 _13264_ (.A(_09801_),
    .B(net3538),
    .Y(_09824_));
 sky130_fd_sc_hd__a22o_1 _13265_ (.A1(_09795_),
    .A2(_09593_),
    .B1(_09798_),
    .B2(_09824_),
    .X(_09825_));
 sky130_fd_sc_hd__inv_2 _13266_ (.A(_09825_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _13267_ (.A(_09236_),
    .B(_09822_),
    .Y(_09826_));
 sky130_fd_sc_hd__a31o_1 _13268_ (.A1(_09712_),
    .A2(net877),
    .A3(_09822_),
    .B1(_09826_),
    .X(_01621_));
 sky130_fd_sc_hd__nand2_1 _13269_ (.A(_09801_),
    .B(net3001),
    .Y(_09827_));
 sky130_fd_sc_hd__a22o_1 _13270_ (.A1(_09795_),
    .A2(_09239_),
    .B1(_09798_),
    .B2(_09827_),
    .X(_09828_));
 sky130_fd_sc_hd__inv_2 _13271_ (.A(_09828_),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _13272_ (.A(_09801_),
    .B(net3201),
    .Y(_09829_));
 sky130_fd_sc_hd__a22o_1 _13273_ (.A1(_09795_),
    .A2(_09768_),
    .B1(_09797_),
    .B2(_09829_),
    .X(_09830_));
 sky130_fd_sc_hd__inv_2 _13274_ (.A(_09830_),
    .Y(_01623_));
 sky130_fd_sc_hd__clkbuf_8 _13275_ (.A(_09302_),
    .X(_09831_));
 sky130_fd_sc_hd__nor2_1 _13276_ (.A(_09246_),
    .B(_09822_),
    .Y(_09832_));
 sky130_fd_sc_hd__a31o_1 _13277_ (.A1(_09831_),
    .A2(net709),
    .A3(_09822_),
    .B1(_09832_),
    .X(_01608_));
 sky130_fd_sc_hd__buf_4 _13278_ (.A(_09359_),
    .X(_09833_));
 sky130_fd_sc_hd__and3_1 _13279_ (.A(_09792_),
    .B(_09345_),
    .C(_09833_),
    .X(_09834_));
 sky130_fd_sc_hd__a31o_1 _13280_ (.A1(_09822_),
    .A2(_09775_),
    .A3(net2570),
    .B1(_09834_),
    .X(_01609_));
 sky130_fd_sc_hd__nor2_1 _13281_ (.A(_09253_),
    .B(_09798_),
    .Y(_09835_));
 sky130_fd_sc_hd__a31o_1 _13282_ (.A1(_09831_),
    .A2(net1475),
    .A3(_09822_),
    .B1(_09835_),
    .X(_01610_));
 sky130_fd_sc_hd__and3_1 _13283_ (.A(_09792_),
    .B(_09351_),
    .C(_09833_),
    .X(_09836_));
 sky130_fd_sc_hd__a31o_1 _13284_ (.A1(_09822_),
    .A2(_09775_),
    .A3(net2575),
    .B1(_09836_),
    .X(_01611_));
 sky130_fd_sc_hd__nand2_1 _13285_ (.A(_09801_),
    .B(net3182),
    .Y(_09837_));
 sky130_fd_sc_hd__a22o_1 _13286_ (.A1(_09795_),
    .A2(_09354_),
    .B1(_09797_),
    .B2(_09837_),
    .X(_09838_));
 sky130_fd_sc_hd__inv_2 _13287_ (.A(_09838_),
    .Y(_01612_));
 sky130_fd_sc_hd__nand2_1 _13288_ (.A(_09801_),
    .B(net3860),
    .Y(_09839_));
 sky130_fd_sc_hd__a22o_1 _13289_ (.A1(_09795_),
    .A2(_09263_),
    .B1(_09797_),
    .B2(_09839_),
    .X(_09840_));
 sky130_fd_sc_hd__inv_2 _13290_ (.A(_09840_),
    .Y(_01613_));
 sky130_fd_sc_hd__and3_1 _13291_ (.A(_09792_),
    .B(_09266_),
    .C(_09833_),
    .X(_09841_));
 sky130_fd_sc_hd__a31o_1 _13292_ (.A1(_09822_),
    .A2(_09775_),
    .A3(net1815),
    .B1(_09841_),
    .X(_01614_));
 sky130_fd_sc_hd__nand2_1 _13293_ (.A(_09801_),
    .B(net3184),
    .Y(_09842_));
 sky130_fd_sc_hd__a22o_1 _13294_ (.A1(_09794_),
    .A2(_09269_),
    .B1(_09797_),
    .B2(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__inv_2 _13295_ (.A(_09843_),
    .Y(_01615_));
 sky130_fd_sc_hd__and3_1 _13296_ (.A(_09792_),
    .B(_09274_),
    .C(_09833_),
    .X(_09844_));
 sky130_fd_sc_hd__a31o_1 _13297_ (.A1(_09822_),
    .A2(_09775_),
    .A3(net2195),
    .B1(_09844_),
    .X(_01600_));
 sky130_fd_sc_hd__nor2_1 _13298_ (.A(_09277_),
    .B(_09798_),
    .Y(_09845_));
 sky130_fd_sc_hd__a31o_1 _13299_ (.A1(_09831_),
    .A2(net1409),
    .A3(_09822_),
    .B1(_09845_),
    .X(_01601_));
 sky130_fd_sc_hd__buf_4 _13300_ (.A(_09716_),
    .X(_09846_));
 sky130_fd_sc_hd__nand2_1 _13301_ (.A(_09846_),
    .B(net3495),
    .Y(_09847_));
 sky130_fd_sc_hd__a22o_1 _13302_ (.A1(_09794_),
    .A2(_09280_),
    .B1(_09797_),
    .B2(_09847_),
    .X(_09848_));
 sky130_fd_sc_hd__inv_2 _13303_ (.A(net3496),
    .Y(_01602_));
 sky130_fd_sc_hd__nand2_1 _13304_ (.A(_09846_),
    .B(net2975),
    .Y(_09849_));
 sky130_fd_sc_hd__a22o_1 _13305_ (.A1(_09794_),
    .A2(_09284_),
    .B1(_09797_),
    .B2(_09849_),
    .X(_09850_));
 sky130_fd_sc_hd__inv_2 _13306_ (.A(_09850_),
    .Y(_01603_));
 sky130_fd_sc_hd__and3_1 _13307_ (.A(_09792_),
    .B(_09373_),
    .C(_09833_),
    .X(_09851_));
 sky130_fd_sc_hd__a31o_1 _13308_ (.A1(_09822_),
    .A2(_09775_),
    .A3(net2597),
    .B1(_09851_),
    .X(_01604_));
 sky130_fd_sc_hd__nand2_1 _13309_ (.A(_09733_),
    .B(net3427),
    .Y(_09852_));
 sky130_fd_sc_hd__o2bb2a_1 _13310_ (.A1_N(_09852_),
    .A2_N(_09822_),
    .B1(_09294_),
    .B2(_09793_),
    .X(_01605_));
 sky130_fd_sc_hd__nand2_1 _13311_ (.A(_09733_),
    .B(net3716),
    .Y(_09853_));
 sky130_fd_sc_hd__o2bb2a_1 _13312_ (.A1_N(_09853_),
    .A2_N(_09822_),
    .B1(_09298_),
    .B2(_09793_),
    .X(_01606_));
 sky130_fd_sc_hd__nor2_1 _13313_ (.A(_09300_),
    .B(_09798_),
    .Y(_09854_));
 sky130_fd_sc_hd__a31o_1 _13314_ (.A1(_09831_),
    .A2(net873),
    .A3(_09822_),
    .B1(_09854_),
    .X(_01607_));
 sky130_fd_sc_hd__and3_2 _13315_ (.A(_09737_),
    .B(_08736_),
    .C(_09380_),
    .X(_09855_));
 sky130_fd_sc_hd__inv_2 _13316_ (.A(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__nor2_4 _13317_ (.A(_08794_),
    .B(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__buf_4 _13318_ (.A(_09857_),
    .X(_09858_));
 sky130_fd_sc_hd__nor2_1 _13319_ (.A(_09625_),
    .B(_09856_),
    .Y(_09859_));
 sky130_fd_sc_hd__inv_2 _13320_ (.A(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__buf_4 _13321_ (.A(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__nand2_1 _13322_ (.A(_09846_),
    .B(net3507),
    .Y(_09862_));
 sky130_fd_sc_hd__a22o_1 _13323_ (.A1(_09858_),
    .A2(_09451_),
    .B1(_09861_),
    .B2(_09862_),
    .X(_09863_));
 sky130_fd_sc_hd__inv_2 _13324_ (.A(_09863_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _13325_ (.A(_09846_),
    .B(net3637),
    .Y(_09864_));
 sky130_fd_sc_hd__a22o_1 _13326_ (.A1(_09858_),
    .A2(_09315_),
    .B1(_09861_),
    .B2(_09864_),
    .X(_09865_));
 sky130_fd_sc_hd__inv_2 _13327_ (.A(_09865_),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _13328_ (.A(_09846_),
    .B(net3613),
    .Y(_09866_));
 sky130_fd_sc_hd__a22o_1 _13329_ (.A1(_09858_),
    .A2(_09460_),
    .B1(_09861_),
    .B2(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__inv_2 _13330_ (.A(_09867_),
    .Y(_01586_));
 sky130_fd_sc_hd__nand2_1 _13331_ (.A(_09846_),
    .B(net3343),
    .Y(_09868_));
 sky130_fd_sc_hd__a22o_1 _13332_ (.A1(_09858_),
    .A2(_09195_),
    .B1(_09861_),
    .B2(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__inv_2 _13333_ (.A(_09869_),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _13334_ (.A(_09846_),
    .B(net3100),
    .Y(_09870_));
 sky130_fd_sc_hd__a22o_1 _13335_ (.A1(_09858_),
    .A2(_09201_),
    .B1(_09861_),
    .B2(_09870_),
    .X(_09871_));
 sky130_fd_sc_hd__inv_2 _13336_ (.A(_09871_),
    .Y(_01588_));
 sky130_fd_sc_hd__nand2_1 _13337_ (.A(_09846_),
    .B(net3288),
    .Y(_09872_));
 sky130_fd_sc_hd__a22o_1 _13338_ (.A1(_09858_),
    .A2(_09205_),
    .B1(_09861_),
    .B2(_09872_),
    .X(_09873_));
 sky130_fd_sc_hd__inv_2 _13339_ (.A(_09873_),
    .Y(_01589_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_09846_),
    .B(net2977),
    .Y(_09874_));
 sky130_fd_sc_hd__a22o_1 _13341_ (.A1(_09858_),
    .A2(_09398_),
    .B1(_09861_),
    .B2(_09874_),
    .X(_09875_));
 sky130_fd_sc_hd__inv_2 _13342_ (.A(_09875_),
    .Y(_01590_));
 sky130_fd_sc_hd__nand2_1 _13343_ (.A(_09846_),
    .B(net3339),
    .Y(_09876_));
 sky130_fd_sc_hd__a22o_1 _13344_ (.A1(_09858_),
    .A2(_09212_),
    .B1(_09861_),
    .B2(_09876_),
    .X(_09877_));
 sky130_fd_sc_hd__inv_2 _13345_ (.A(_09877_),
    .Y(_01591_));
 sky130_fd_sc_hd__nand2_1 _13346_ (.A(_09846_),
    .B(net3362),
    .Y(_09878_));
 sky130_fd_sc_hd__a22o_1 _13347_ (.A1(_09858_),
    .A2(_09531_),
    .B1(_09861_),
    .B2(_09878_),
    .X(_09879_));
 sky130_fd_sc_hd__inv_2 _13348_ (.A(_09879_),
    .Y(_01576_));
 sky130_fd_sc_hd__nand2_1 _13349_ (.A(_09846_),
    .B(net3092),
    .Y(_09880_));
 sky130_fd_sc_hd__a22o_1 _13350_ (.A1(_09858_),
    .A2(_09219_),
    .B1(_09861_),
    .B2(_09880_),
    .X(_09881_));
 sky130_fd_sc_hd__inv_2 _13351_ (.A(_09881_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand2_1 _13352_ (.A(_09846_),
    .B(net3259),
    .Y(_09882_));
 sky130_fd_sc_hd__a22o_1 _13353_ (.A1(_09858_),
    .A2(_09332_),
    .B1(_09861_),
    .B2(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__inv_2 _13354_ (.A(_09883_),
    .Y(_01578_));
 sky130_fd_sc_hd__nand2_1 _13355_ (.A(_09846_),
    .B(net2845),
    .Y(_09884_));
 sky130_fd_sc_hd__a22o_1 _13356_ (.A1(_09858_),
    .A2(_09589_),
    .B1(_09861_),
    .B2(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__inv_2 _13357_ (.A(_09885_),
    .Y(_01579_));
 sky130_fd_sc_hd__nand2_1 _13358_ (.A(_09846_),
    .B(net2850),
    .Y(_09886_));
 sky130_fd_sc_hd__a22o_1 _13359_ (.A1(_09858_),
    .A2(_09593_),
    .B1(_09861_),
    .B2(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__inv_2 _13360_ (.A(_09887_),
    .Y(_01580_));
 sky130_fd_sc_hd__buf_4 _13361_ (.A(_09860_),
    .X(_09888_));
 sky130_fd_sc_hd__nand2_1 _13362_ (.A(_09846_),
    .B(net3347),
    .Y(_09889_));
 sky130_fd_sc_hd__a22o_1 _13363_ (.A1(_09858_),
    .A2(_09338_),
    .B1(_09888_),
    .B2(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__inv_2 _13364_ (.A(_09890_),
    .Y(_01581_));
 sky130_fd_sc_hd__buf_4 _13365_ (.A(_09716_),
    .X(_09891_));
 sky130_fd_sc_hd__nand2_1 _13366_ (.A(_09891_),
    .B(net3179),
    .Y(_09892_));
 sky130_fd_sc_hd__a22o_1 _13367_ (.A1(_09858_),
    .A2(_09239_),
    .B1(_09888_),
    .B2(_09892_),
    .X(_09893_));
 sky130_fd_sc_hd__inv_2 _13368_ (.A(_09893_),
    .Y(_01582_));
 sky130_fd_sc_hd__nand2_1 _13369_ (.A(_09891_),
    .B(net3655),
    .Y(_09894_));
 sky130_fd_sc_hd__a22o_1 _13370_ (.A1(_09858_),
    .A2(_09768_),
    .B1(_09888_),
    .B2(_09894_),
    .X(_09895_));
 sky130_fd_sc_hd__inv_2 _13371_ (.A(_09895_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _13372_ (.A(_09891_),
    .B(net3178),
    .Y(_09896_));
 sky130_fd_sc_hd__a22o_1 _13373_ (.A1(_09857_),
    .A2(_09415_),
    .B1(_09888_),
    .B2(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__inv_2 _13374_ (.A(_09897_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand2_1 _13375_ (.A(_09891_),
    .B(net3158),
    .Y(_09898_));
 sky130_fd_sc_hd__a22o_1 _13376_ (.A1(_09857_),
    .A2(_09249_),
    .B1(_09888_),
    .B2(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__inv_2 _13377_ (.A(_09899_),
    .Y(_01569_));
 sky130_fd_sc_hd__nand2_1 _13378_ (.A(_09891_),
    .B(net3367),
    .Y(_09900_));
 sky130_fd_sc_hd__a22o_1 _13379_ (.A1(_09857_),
    .A2(_09348_),
    .B1(_09888_),
    .B2(_09900_),
    .X(_09901_));
 sky130_fd_sc_hd__inv_2 _13380_ (.A(_09901_),
    .Y(_01570_));
 sky130_fd_sc_hd__nand2_1 _13381_ (.A(_09891_),
    .B(net3360),
    .Y(_09902_));
 sky130_fd_sc_hd__a22o_1 _13382_ (.A1(_09857_),
    .A2(_09256_),
    .B1(_09888_),
    .B2(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__inv_2 _13383_ (.A(_09903_),
    .Y(_01571_));
 sky130_fd_sc_hd__nand2_1 _13384_ (.A(_09891_),
    .B(net3047),
    .Y(_09904_));
 sky130_fd_sc_hd__a22o_1 _13385_ (.A1(_09857_),
    .A2(_09354_),
    .B1(_09888_),
    .B2(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__inv_2 _13386_ (.A(_09905_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_1 _13387_ (.A(_09891_),
    .B(net3852),
    .Y(_09906_));
 sky130_fd_sc_hd__a22o_1 _13388_ (.A1(_09857_),
    .A2(_09263_),
    .B1(_09888_),
    .B2(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__inv_2 _13389_ (.A(_09907_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand2_1 _13390_ (.A(_09891_),
    .B(net3933),
    .Y(_09908_));
 sky130_fd_sc_hd__a22o_1 _13391_ (.A1(_09857_),
    .A2(_09425_),
    .B1(_09888_),
    .B2(_09908_),
    .X(_09909_));
 sky130_fd_sc_hd__inv_2 _13392_ (.A(_09909_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _13393_ (.A(_09891_),
    .B(net3453),
    .Y(_09910_));
 sky130_fd_sc_hd__a22o_1 _13394_ (.A1(_09857_),
    .A2(_09269_),
    .B1(_09888_),
    .B2(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__inv_2 _13395_ (.A(_09911_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2_1 _13396_ (.A(_09891_),
    .B(net3648),
    .Y(_09912_));
 sky130_fd_sc_hd__a22o_1 _13397_ (.A1(_09857_),
    .A2(_09495_),
    .B1(_09888_),
    .B2(_09912_),
    .X(_09913_));
 sky130_fd_sc_hd__inv_2 _13398_ (.A(_09913_),
    .Y(_01560_));
 sky130_fd_sc_hd__nand2_1 _13399_ (.A(_09891_),
    .B(net3477),
    .Y(_09914_));
 sky130_fd_sc_hd__a22o_1 _13400_ (.A1(_09857_),
    .A2(_09366_),
    .B1(_09888_),
    .B2(_09914_),
    .X(_09915_));
 sky130_fd_sc_hd__inv_2 _13401_ (.A(_09915_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _13402_ (.A(_09891_),
    .B(net3043),
    .Y(_09916_));
 sky130_fd_sc_hd__a22o_1 _13403_ (.A1(_09857_),
    .A2(_09280_),
    .B1(_09888_),
    .B2(_09916_),
    .X(_09917_));
 sky130_fd_sc_hd__inv_2 _13404_ (.A(_09917_),
    .Y(_01562_));
 sky130_fd_sc_hd__nand2_1 _13405_ (.A(_09891_),
    .B(net2954),
    .Y(_09918_));
 sky130_fd_sc_hd__a22o_1 _13406_ (.A1(_09857_),
    .A2(_09284_),
    .B1(_09888_),
    .B2(_09918_),
    .X(_09919_));
 sky130_fd_sc_hd__inv_2 _13407_ (.A(_09919_),
    .Y(_01563_));
 sky130_fd_sc_hd__nand2_1 _13408_ (.A(_09891_),
    .B(net3406),
    .Y(_09920_));
 sky130_fd_sc_hd__a22o_1 _13409_ (.A1(_09857_),
    .A2(_09288_),
    .B1(_09888_),
    .B2(_09920_),
    .X(_09921_));
 sky130_fd_sc_hd__inv_2 _13410_ (.A(_09921_),
    .Y(_01564_));
 sky130_fd_sc_hd__nand2_1 _13411_ (.A(_09733_),
    .B(net3692),
    .Y(_09922_));
 sky130_fd_sc_hd__o2bb2a_1 _13412_ (.A1_N(_09922_),
    .A2_N(_09861_),
    .B1(_09294_),
    .B2(_09856_),
    .X(_01565_));
 sky130_fd_sc_hd__nand2_1 _13413_ (.A(_09733_),
    .B(net3725),
    .Y(_09923_));
 sky130_fd_sc_hd__o2bb2a_1 _13414_ (.A1_N(_09923_),
    .A2_N(_09861_),
    .B1(_09298_),
    .B2(_09856_),
    .X(_01566_));
 sky130_fd_sc_hd__nand2_1 _13415_ (.A(_09733_),
    .B(net3601),
    .Y(_09924_));
 sky130_fd_sc_hd__o2bb2a_1 _13416_ (.A1_N(_09924_),
    .A2_N(_09861_),
    .B1(_09442_),
    .B2(_09856_),
    .X(_01567_));
 sky130_fd_sc_hd__nand2_2 _13417_ (.A(_09737_),
    .B(_09445_),
    .Y(_09925_));
 sky130_fd_sc_hd__nor2_4 _13418_ (.A(_09444_),
    .B(_09925_),
    .Y(_09926_));
 sky130_fd_sc_hd__inv_2 _13419_ (.A(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__nor2_1 _13420_ (.A(_09625_),
    .B(_09927_),
    .Y(_09928_));
 sky130_fd_sc_hd__inv_2 _13421_ (.A(_09928_),
    .Y(_09929_));
 sky130_fd_sc_hd__buf_4 _13422_ (.A(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__buf_4 _13423_ (.A(_09929_),
    .X(_09931_));
 sky130_fd_sc_hd__nor2_1 _13424_ (.A(_09181_),
    .B(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__a31o_1 _13425_ (.A1(_09831_),
    .A2(net859),
    .A3(_09930_),
    .B1(_09932_),
    .X(_01552_));
 sky130_fd_sc_hd__nor2_1 _13426_ (.A(_09185_),
    .B(_09931_),
    .Y(_09933_));
 sky130_fd_sc_hd__a31o_1 _13427_ (.A1(_09831_),
    .A2(net1626),
    .A3(_09930_),
    .B1(_09933_),
    .X(_01553_));
 sky130_fd_sc_hd__nor2_1 _13428_ (.A(_09188_),
    .B(_09931_),
    .Y(_09934_));
 sky130_fd_sc_hd__a31o_1 _13429_ (.A1(_09831_),
    .A2(net2594),
    .A3(_09930_),
    .B1(_09934_),
    .X(_01554_));
 sky130_fd_sc_hd__nor2_8 _13430_ (.A(_08797_),
    .B(_09927_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_1 _13431_ (.A(_09891_),
    .B(net3727),
    .Y(_09936_));
 sky130_fd_sc_hd__a22o_1 _13432_ (.A1(_09935_),
    .A2(_09195_),
    .B1(_09931_),
    .B2(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__inv_2 _13433_ (.A(_09937_),
    .Y(_01555_));
 sky130_fd_sc_hd__buf_4 _13434_ (.A(_09716_),
    .X(_09938_));
 sky130_fd_sc_hd__nand2_1 _13435_ (.A(_09938_),
    .B(net3210),
    .Y(_09939_));
 sky130_fd_sc_hd__a22o_1 _13436_ (.A1(_09935_),
    .A2(_09201_),
    .B1(_09931_),
    .B2(_09939_),
    .X(_09940_));
 sky130_fd_sc_hd__inv_2 _13437_ (.A(_09940_),
    .Y(_01556_));
 sky130_fd_sc_hd__and3_1 _13438_ (.A(_09926_),
    .B(_09395_),
    .C(_09833_),
    .X(_09941_));
 sky130_fd_sc_hd__a31o_1 _13439_ (.A1(_09930_),
    .A2(_09775_),
    .A3(net2017),
    .B1(_09941_),
    .X(_01557_));
 sky130_fd_sc_hd__nand2_1 _13440_ (.A(_09938_),
    .B(net3123),
    .Y(_09942_));
 sky130_fd_sc_hd__a22o_1 _13441_ (.A1(_09935_),
    .A2(_09398_),
    .B1(_09931_),
    .B2(_09942_),
    .X(_09943_));
 sky130_fd_sc_hd__inv_2 _13442_ (.A(_09943_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_1 _13443_ (.A(_09938_),
    .B(net4082),
    .Y(_09944_));
 sky130_fd_sc_hd__a22o_1 _13444_ (.A1(_09935_),
    .A2(_09212_),
    .B1(_09931_),
    .B2(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__inv_2 _13445_ (.A(_09945_),
    .Y(_01559_));
 sky130_fd_sc_hd__nor2_1 _13446_ (.A(_09216_),
    .B(_09931_),
    .Y(_09946_));
 sky130_fd_sc_hd__a31o_1 _13447_ (.A1(_09831_),
    .A2(net2312),
    .A3(_09930_),
    .B1(_09946_),
    .X(_01544_));
 sky130_fd_sc_hd__nand2_1 _13448_ (.A(_09938_),
    .B(net2931),
    .Y(_09947_));
 sky130_fd_sc_hd__a22o_1 _13449_ (.A1(_09935_),
    .A2(_09219_),
    .B1(_09931_),
    .B2(_09947_),
    .X(_09948_));
 sky130_fd_sc_hd__inv_2 _13450_ (.A(_09948_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_1 _13451_ (.A(_09938_),
    .B(net2918),
    .Y(_09949_));
 sky130_fd_sc_hd__a22o_1 _13452_ (.A1(_09935_),
    .A2(_09332_),
    .B1(_09931_),
    .B2(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__inv_2 _13453_ (.A(_09950_),
    .Y(_01546_));
 sky130_fd_sc_hd__nor2_1 _13454_ (.A(_09230_),
    .B(_09931_),
    .Y(_09951_));
 sky130_fd_sc_hd__a31o_1 _13455_ (.A1(_09831_),
    .A2(net1932),
    .A3(_09930_),
    .B1(_09951_),
    .X(_01547_));
 sky130_fd_sc_hd__nand2_1 _13456_ (.A(_09938_),
    .B(net3076),
    .Y(_09952_));
 sky130_fd_sc_hd__a22o_1 _13457_ (.A1(_09935_),
    .A2(_09593_),
    .B1(_09931_),
    .B2(_09952_),
    .X(_09953_));
 sky130_fd_sc_hd__inv_2 _13458_ (.A(_09953_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _13459_ (.A(_09236_),
    .B(_09931_),
    .Y(_09954_));
 sky130_fd_sc_hd__a31o_1 _13460_ (.A1(_09831_),
    .A2(net2127),
    .A3(_09930_),
    .B1(_09954_),
    .X(_01549_));
 sky130_fd_sc_hd__and3_1 _13461_ (.A(_09926_),
    .B(_09341_),
    .C(_09833_),
    .X(_09955_));
 sky130_fd_sc_hd__a31o_1 _13462_ (.A1(_09930_),
    .A2(_09775_),
    .A3(net1910),
    .B1(_09955_),
    .X(_01550_));
 sky130_fd_sc_hd__nor2_1 _13463_ (.A(_09243_),
    .B(_09931_),
    .Y(_09956_));
 sky130_fd_sc_hd__a31o_1 _13464_ (.A1(_09831_),
    .A2(net2182),
    .A3(_09930_),
    .B1(_09956_),
    .X(_01551_));
 sky130_fd_sc_hd__nand2_1 _13465_ (.A(_09938_),
    .B(net3096),
    .Y(_09957_));
 sky130_fd_sc_hd__a22o_1 _13466_ (.A1(_09935_),
    .A2(_09415_),
    .B1(_09929_),
    .B2(_09957_),
    .X(_09958_));
 sky130_fd_sc_hd__inv_2 _13467_ (.A(_09958_),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _13468_ (.A(_09938_),
    .B(net3666),
    .Y(_09959_));
 sky130_fd_sc_hd__a22o_1 _13469_ (.A1(_09935_),
    .A2(_09249_),
    .B1(_09929_),
    .B2(_09959_),
    .X(_09960_));
 sky130_fd_sc_hd__inv_2 _13470_ (.A(_09960_),
    .Y(_01537_));
 sky130_fd_sc_hd__nor2_1 _13471_ (.A(_09253_),
    .B(_09931_),
    .Y(_09961_));
 sky130_fd_sc_hd__a31o_1 _13472_ (.A1(_09831_),
    .A2(net2667),
    .A3(_09931_),
    .B1(_09961_),
    .X(_01538_));
 sky130_fd_sc_hd__and3_1 _13473_ (.A(_09926_),
    .B(_09351_),
    .C(_09833_),
    .X(_09962_));
 sky130_fd_sc_hd__a31o_1 _13474_ (.A1(_09930_),
    .A2(_09775_),
    .A3(net2580),
    .B1(_09962_),
    .X(_01539_));
 sky130_fd_sc_hd__nand2_1 _13475_ (.A(_09938_),
    .B(net2982),
    .Y(_09963_));
 sky130_fd_sc_hd__a22o_1 _13476_ (.A1(_09935_),
    .A2(_09354_),
    .B1(_09929_),
    .B2(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__inv_2 _13477_ (.A(_09964_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand2_1 _13478_ (.A(_09938_),
    .B(net3020),
    .Y(_09965_));
 sky130_fd_sc_hd__a22o_1 _13479_ (.A1(_09935_),
    .A2(_09263_),
    .B1(_09929_),
    .B2(_09965_),
    .X(_09966_));
 sky130_fd_sc_hd__inv_2 _13480_ (.A(_09966_),
    .Y(_01541_));
 sky130_fd_sc_hd__and3_1 _13481_ (.A(_09926_),
    .B(_09266_),
    .C(_09833_),
    .X(_09967_));
 sky130_fd_sc_hd__a31o_1 _13482_ (.A1(_09930_),
    .A2(_09775_),
    .A3(net2636),
    .B1(_09967_),
    .X(_01542_));
 sky130_fd_sc_hd__nand2_1 _13483_ (.A(_09938_),
    .B(net3455),
    .Y(_09968_));
 sky130_fd_sc_hd__a22o_1 _13484_ (.A1(_09935_),
    .A2(_09269_),
    .B1(_09929_),
    .B2(_09968_),
    .X(_09969_));
 sky130_fd_sc_hd__inv_2 _13485_ (.A(_09969_),
    .Y(_01543_));
 sky130_fd_sc_hd__and3_1 _13486_ (.A(_09926_),
    .B(_09274_),
    .C(_09833_),
    .X(_09970_));
 sky130_fd_sc_hd__a31o_1 _13487_ (.A1(_09930_),
    .A2(_09775_),
    .A3(net2613),
    .B1(_09970_),
    .X(_01528_));
 sky130_fd_sc_hd__nand2_1 _13488_ (.A(_09938_),
    .B(net3431),
    .Y(_09971_));
 sky130_fd_sc_hd__a22o_1 _13489_ (.A1(_09935_),
    .A2(_09366_),
    .B1(_09929_),
    .B2(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__inv_2 _13490_ (.A(_09972_),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_1 _13491_ (.A(_09938_),
    .B(net3594),
    .Y(_09973_));
 sky130_fd_sc_hd__a22o_1 _13492_ (.A1(_09935_),
    .A2(_09280_),
    .B1(_09929_),
    .B2(_09973_),
    .X(_09974_));
 sky130_fd_sc_hd__inv_2 _13493_ (.A(_09974_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand2_1 _13494_ (.A(_09938_),
    .B(net3539),
    .Y(_09975_));
 sky130_fd_sc_hd__a22o_1 _13495_ (.A1(_09935_),
    .A2(_09284_),
    .B1(_09929_),
    .B2(_09975_),
    .X(_09976_));
 sky130_fd_sc_hd__inv_2 _13496_ (.A(_09976_),
    .Y(_01531_));
 sky130_fd_sc_hd__buf_4 _13497_ (.A(_09223_),
    .X(_09977_));
 sky130_fd_sc_hd__and3_1 _13498_ (.A(_09926_),
    .B(_09373_),
    .C(_09833_),
    .X(_09978_));
 sky130_fd_sc_hd__a31o_1 _13499_ (.A1(_09930_),
    .A2(_09977_),
    .A3(net2624),
    .B1(_09978_),
    .X(_01532_));
 sky130_fd_sc_hd__and3_1 _13500_ (.A(_09926_),
    .B(_09730_),
    .C(_09833_),
    .X(_09979_));
 sky130_fd_sc_hd__a31o_1 _13501_ (.A1(_09930_),
    .A2(_09977_),
    .A3(net1986),
    .B1(_09979_),
    .X(_01533_));
 sky130_fd_sc_hd__nand2_1 _13502_ (.A(_09733_),
    .B(net3820),
    .Y(_09980_));
 sky130_fd_sc_hd__o2bb2a_1 _13503_ (.A1_N(_09980_),
    .A2_N(_09930_),
    .B1(_09298_),
    .B2(_09927_),
    .X(_01534_));
 sky130_fd_sc_hd__nand2_1 _13504_ (.A(_09733_),
    .B(net3678),
    .Y(_09981_));
 sky130_fd_sc_hd__o2bb2a_1 _13505_ (.A1_N(_09981_),
    .A2_N(_09930_),
    .B1(_09442_),
    .B2(_09927_),
    .X(_01535_));
 sky130_fd_sc_hd__nor2_8 _13506_ (.A(net2787),
    .B(net3791),
    .Y(_09982_));
 sky130_fd_sc_hd__nand2_1 _13507_ (.A(_09169_),
    .B(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__or2_2 _13508_ (.A(_09172_),
    .B(_09983_),
    .X(_09984_));
 sky130_fd_sc_hd__nor2_4 _13509_ (.A(_09444_),
    .B(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__inv_2 _13510_ (.A(_09985_),
    .Y(_09986_));
 sky130_fd_sc_hd__nor2_4 _13511_ (.A(_09190_),
    .B(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__nor2_1 _13512_ (.A(_09166_),
    .B(_09986_),
    .Y(_09988_));
 sky130_fd_sc_hd__inv_2 _13513_ (.A(_09988_),
    .Y(_09989_));
 sky130_fd_sc_hd__buf_4 _13514_ (.A(_09989_),
    .X(_09990_));
 sky130_fd_sc_hd__nand2_1 _13515_ (.A(_09938_),
    .B(net4330),
    .Y(_09991_));
 sky130_fd_sc_hd__a22o_1 _13516_ (.A1(_09987_),
    .A2(_09451_),
    .B1(_09990_),
    .B2(_09991_),
    .X(_09992_));
 sky130_fd_sc_hd__inv_2 _13517_ (.A(_09992_),
    .Y(_01520_));
 sky130_fd_sc_hd__buf_4 _13518_ (.A(_09989_),
    .X(_09993_));
 sky130_fd_sc_hd__nor2_1 _13519_ (.A(_09185_),
    .B(_09990_),
    .Y(_09994_));
 sky130_fd_sc_hd__a31o_1 _13520_ (.A1(_09831_),
    .A2(net2654),
    .A3(_09993_),
    .B1(_09994_),
    .X(_01521_));
 sky130_fd_sc_hd__nor2_1 _13521_ (.A(_09188_),
    .B(_09990_),
    .Y(_09995_));
 sky130_fd_sc_hd__a31o_1 _13522_ (.A1(_09831_),
    .A2(net2666),
    .A3(_09993_),
    .B1(_09995_),
    .X(_01522_));
 sky130_fd_sc_hd__and3_1 _13523_ (.A(_09985_),
    .B(_09463_),
    .C(_09833_),
    .X(_09996_));
 sky130_fd_sc_hd__a31o_1 _13524_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2642),
    .B1(_09996_),
    .X(_01523_));
 sky130_fd_sc_hd__and3_1 _13525_ (.A(_09985_),
    .B(_09321_),
    .C(_09833_),
    .X(_09997_));
 sky130_fd_sc_hd__a31o_1 _13526_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2657),
    .B1(_09997_),
    .X(_01524_));
 sky130_fd_sc_hd__and3_1 _13527_ (.A(_09985_),
    .B(_09395_),
    .C(_09833_),
    .X(_09998_));
 sky130_fd_sc_hd__a31o_1 _13528_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2694),
    .B1(_09998_),
    .X(_01525_));
 sky130_fd_sc_hd__nand2_1 _13529_ (.A(_09938_),
    .B(net4251),
    .Y(_09999_));
 sky130_fd_sc_hd__a22o_1 _13530_ (.A1(_09987_),
    .A2(_09398_),
    .B1(_09990_),
    .B2(_09999_),
    .X(_10000_));
 sky130_fd_sc_hd__inv_2 _13531_ (.A(_10000_),
    .Y(_01526_));
 sky130_fd_sc_hd__buf_4 _13532_ (.A(_09716_),
    .X(_10001_));
 sky130_fd_sc_hd__nand2_1 _13533_ (.A(_10001_),
    .B(net4308),
    .Y(_10002_));
 sky130_fd_sc_hd__a22o_1 _13534_ (.A1(_09987_),
    .A2(_09212_),
    .B1(_09990_),
    .B2(_10002_),
    .X(_10003_));
 sky130_fd_sc_hd__inv_2 _13535_ (.A(_10003_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _13536_ (.A(_09216_),
    .B(_09990_),
    .Y(_10004_));
 sky130_fd_sc_hd__a31o_1 _13537_ (.A1(_09831_),
    .A2(net2627),
    .A3(_09993_),
    .B1(_10004_),
    .X(_01512_));
 sky130_fd_sc_hd__nand2_1 _13538_ (.A(_10001_),
    .B(net3209),
    .Y(_10005_));
 sky130_fd_sc_hd__a22o_1 _13539_ (.A1(_09987_),
    .A2(_09219_),
    .B1(_09990_),
    .B2(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__inv_2 _13540_ (.A(_10006_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_1 _13541_ (.A(_10001_),
    .B(net2885),
    .Y(_10007_));
 sky130_fd_sc_hd__a22o_1 _13542_ (.A1(_09987_),
    .A2(_09332_),
    .B1(_09989_),
    .B2(_10007_),
    .X(_10008_));
 sky130_fd_sc_hd__inv_2 _13543_ (.A(_10008_),
    .Y(_01514_));
 sky130_fd_sc_hd__nor2_1 _13544_ (.A(_09230_),
    .B(_09990_),
    .Y(_10009_));
 sky130_fd_sc_hd__a31o_1 _13545_ (.A1(_09831_),
    .A2(net1735),
    .A3(_09993_),
    .B1(_10009_),
    .X(_01515_));
 sky130_fd_sc_hd__clkbuf_8 _13546_ (.A(_09302_),
    .X(_10010_));
 sky130_fd_sc_hd__nor2_1 _13547_ (.A(_09233_),
    .B(_09990_),
    .Y(_10011_));
 sky130_fd_sc_hd__a31o_1 _13548_ (.A1(_10010_),
    .A2(net1153),
    .A3(_09993_),
    .B1(_10011_),
    .X(_01516_));
 sky130_fd_sc_hd__nand2_1 _13549_ (.A(_10001_),
    .B(net3505),
    .Y(_10012_));
 sky130_fd_sc_hd__a22o_1 _13550_ (.A1(_09987_),
    .A2(_09338_),
    .B1(_09989_),
    .B2(_10012_),
    .X(_10013_));
 sky130_fd_sc_hd__inv_2 _13551_ (.A(_10013_),
    .Y(_01517_));
 sky130_fd_sc_hd__and3_1 _13552_ (.A(_09985_),
    .B(_09341_),
    .C(_09833_),
    .X(_10014_));
 sky130_fd_sc_hd__a31o_1 _13553_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2292),
    .B1(_10014_),
    .X(_01518_));
 sky130_fd_sc_hd__nand2_1 _13554_ (.A(_10001_),
    .B(net3191),
    .Y(_10015_));
 sky130_fd_sc_hd__a22o_1 _13555_ (.A1(_09987_),
    .A2(_09768_),
    .B1(_09989_),
    .B2(_10015_),
    .X(_10016_));
 sky130_fd_sc_hd__inv_2 _13556_ (.A(_10016_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _13557_ (.A(_10001_),
    .B(net3520),
    .Y(_10017_));
 sky130_fd_sc_hd__a22o_1 _13558_ (.A1(_09987_),
    .A2(_09415_),
    .B1(_09989_),
    .B2(_10017_),
    .X(_10018_));
 sky130_fd_sc_hd__inv_2 _13559_ (.A(_10018_),
    .Y(_01496_));
 sky130_fd_sc_hd__clkbuf_4 _13560_ (.A(_09359_),
    .X(_10019_));
 sky130_fd_sc_hd__and3_1 _13561_ (.A(_09985_),
    .B(_09345_),
    .C(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__a31o_1 _13562_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2499),
    .B1(_10020_),
    .X(_01497_));
 sky130_fd_sc_hd__nor2_1 _13563_ (.A(_09253_),
    .B(_09990_),
    .Y(_10021_));
 sky130_fd_sc_hd__a31o_1 _13564_ (.A1(_10010_),
    .A2(net2003),
    .A3(_09993_),
    .B1(_10021_),
    .X(_01498_));
 sky130_fd_sc_hd__nand2_1 _13565_ (.A(_10001_),
    .B(net2902),
    .Y(_10022_));
 sky130_fd_sc_hd__a22o_1 _13566_ (.A1(_09987_),
    .A2(_09256_),
    .B1(_09989_),
    .B2(_10022_),
    .X(_10023_));
 sky130_fd_sc_hd__inv_2 _13567_ (.A(_10023_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _13568_ (.A(_09260_),
    .B(_09990_),
    .Y(_10024_));
 sky130_fd_sc_hd__a31o_1 _13569_ (.A1(_10010_),
    .A2(net1349),
    .A3(_09990_),
    .B1(_10024_),
    .X(_01500_));
 sky130_fd_sc_hd__nand2_1 _13570_ (.A(_10001_),
    .B(net2876),
    .Y(_10025_));
 sky130_fd_sc_hd__a22o_1 _13571_ (.A1(_09987_),
    .A2(_09263_),
    .B1(_09989_),
    .B2(_10025_),
    .X(_10026_));
 sky130_fd_sc_hd__inv_2 _13572_ (.A(_10026_),
    .Y(_01501_));
 sky130_fd_sc_hd__nand2_1 _13573_ (.A(_10001_),
    .B(net3164),
    .Y(_10027_));
 sky130_fd_sc_hd__a22o_1 _13574_ (.A1(_09987_),
    .A2(_09425_),
    .B1(_09989_),
    .B2(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__inv_2 _13575_ (.A(_10028_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand2_1 _13576_ (.A(_10001_),
    .B(net3102),
    .Y(_10029_));
 sky130_fd_sc_hd__a22o_1 _13577_ (.A1(_09987_),
    .A2(_09269_),
    .B1(_09989_),
    .B2(_10029_),
    .X(_10030_));
 sky130_fd_sc_hd__inv_2 _13578_ (.A(_10030_),
    .Y(_01503_));
 sky130_fd_sc_hd__and3_1 _13579_ (.A(_09985_),
    .B(_09274_),
    .C(_10019_),
    .X(_10031_));
 sky130_fd_sc_hd__a31o_1 _13580_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2105),
    .B1(_10031_),
    .X(_01488_));
 sky130_fd_sc_hd__nor2_1 _13581_ (.A(_09277_),
    .B(_09990_),
    .Y(_10032_));
 sky130_fd_sc_hd__a31o_1 _13582_ (.A1(_10010_),
    .A2(net2480),
    .A3(_09990_),
    .B1(_10032_),
    .X(_01489_));
 sky130_fd_sc_hd__and3_1 _13583_ (.A(_09985_),
    .B(_09369_),
    .C(_10019_),
    .X(_10033_));
 sky130_fd_sc_hd__a31o_1 _13584_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2607),
    .B1(_10033_),
    .X(_01490_));
 sky130_fd_sc_hd__nand2_1 _13585_ (.A(_10001_),
    .B(net3904),
    .Y(_10034_));
 sky130_fd_sc_hd__a22o_1 _13586_ (.A1(_09987_),
    .A2(_09284_),
    .B1(_09989_),
    .B2(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__inv_2 _13587_ (.A(_10035_),
    .Y(_01491_));
 sky130_fd_sc_hd__and3_1 _13588_ (.A(_09985_),
    .B(_09373_),
    .C(_10019_),
    .X(_10036_));
 sky130_fd_sc_hd__a31o_1 _13589_ (.A1(_09993_),
    .A2(_09977_),
    .A3(net2382),
    .B1(_10036_),
    .X(_01492_));
 sky130_fd_sc_hd__nand2_1 _13590_ (.A(_09733_),
    .B(net3869),
    .Y(_10037_));
 sky130_fd_sc_hd__o2bb2a_1 _13591_ (.A1_N(_10037_),
    .A2_N(_09993_),
    .B1(_09294_),
    .B2(_09986_),
    .X(_01493_));
 sky130_fd_sc_hd__nand2_1 _13592_ (.A(_09733_),
    .B(net4008),
    .Y(_10038_));
 sky130_fd_sc_hd__o2bb2a_1 _13593_ (.A1_N(_10038_),
    .A2_N(_09993_),
    .B1(_09298_),
    .B2(_09986_),
    .X(_01494_));
 sky130_fd_sc_hd__nor2_1 _13594_ (.A(_09300_),
    .B(_09990_),
    .Y(_10039_));
 sky130_fd_sc_hd__a31o_1 _13595_ (.A1(_10010_),
    .A2(net1607),
    .A3(_09990_),
    .B1(_10039_),
    .X(_01495_));
 sky130_fd_sc_hd__inv_2 _13596_ (.A(_09305_),
    .Y(_10040_));
 sky130_fd_sc_hd__or2_2 _13597_ (.A(_10040_),
    .B(_09983_),
    .X(_10041_));
 sky130_fd_sc_hd__nor2_4 _13598_ (.A(_09444_),
    .B(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__inv_2 _13599_ (.A(_10042_),
    .Y(_10043_));
 sky130_fd_sc_hd__nor2_1 _13600_ (.A(_09304_),
    .B(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__clkinv_4 _13601_ (.A(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__buf_4 _13602_ (.A(_10045_),
    .X(_10046_));
 sky130_fd_sc_hd__buf_4 _13603_ (.A(_10045_),
    .X(_10047_));
 sky130_fd_sc_hd__nor2_1 _13604_ (.A(_09181_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__a31o_1 _13605_ (.A1(_10010_),
    .A2(net509),
    .A3(_10046_),
    .B1(_10048_),
    .X(_01480_));
 sky130_fd_sc_hd__nor2_1 _13606_ (.A(_09185_),
    .B(_10047_),
    .Y(_10049_));
 sky130_fd_sc_hd__a31o_1 _13607_ (.A1(_10010_),
    .A2(net931),
    .A3(_10046_),
    .B1(_10049_),
    .X(_01481_));
 sky130_fd_sc_hd__nor2_1 _13608_ (.A(_09188_),
    .B(_10047_),
    .Y(_10050_));
 sky130_fd_sc_hd__a31o_1 _13609_ (.A1(_10010_),
    .A2(net643),
    .A3(_10046_),
    .B1(_10050_),
    .X(_01482_));
 sky130_fd_sc_hd__and3_1 _13610_ (.A(_10042_),
    .B(_09463_),
    .C(_10019_),
    .X(_10051_));
 sky130_fd_sc_hd__a31o_1 _13611_ (.A1(_10046_),
    .A2(_09977_),
    .A3(net583),
    .B1(_10051_),
    .X(_01483_));
 sky130_fd_sc_hd__and3_1 _13612_ (.A(_10042_),
    .B(_09321_),
    .C(_10019_),
    .X(_10052_));
 sky130_fd_sc_hd__a31o_1 _13613_ (.A1(_10046_),
    .A2(_09977_),
    .A3(net1179),
    .B1(_10052_),
    .X(_01484_));
 sky130_fd_sc_hd__nor2_4 _13614_ (.A(_08795_),
    .B(_10043_),
    .Y(_10053_));
 sky130_fd_sc_hd__nand2_1 _13615_ (.A(_10001_),
    .B(net2866),
    .Y(_10054_));
 sky130_fd_sc_hd__a22o_1 _13616_ (.A1(_10053_),
    .A2(_09205_),
    .B1(_10047_),
    .B2(_10054_),
    .X(_10055_));
 sky130_fd_sc_hd__inv_2 _13617_ (.A(_10055_),
    .Y(_01485_));
 sky130_fd_sc_hd__nor2_1 _13618_ (.A(_09209_),
    .B(_10047_),
    .Y(_10056_));
 sky130_fd_sc_hd__a31o_1 _13619_ (.A1(_10010_),
    .A2(net557),
    .A3(_10046_),
    .B1(_10056_),
    .X(_01486_));
 sky130_fd_sc_hd__and3_1 _13620_ (.A(_10042_),
    .B(_09326_),
    .C(_10019_),
    .X(_10057_));
 sky130_fd_sc_hd__a31o_1 _13621_ (.A1(_10046_),
    .A2(_09977_),
    .A3(net1447),
    .B1(_10057_),
    .X(_01487_));
 sky130_fd_sc_hd__nand2_1 _13622_ (.A(_10001_),
    .B(net3168),
    .Y(_10058_));
 sky130_fd_sc_hd__a22o_1 _13623_ (.A1(_10053_),
    .A2(_09531_),
    .B1(_10047_),
    .B2(_10058_),
    .X(_10059_));
 sky130_fd_sc_hd__inv_2 _13624_ (.A(_10059_),
    .Y(_01472_));
 sky130_fd_sc_hd__nand2_1 _13625_ (.A(_10001_),
    .B(net3524),
    .Y(_10060_));
 sky130_fd_sc_hd__a22o_1 _13626_ (.A1(_10053_),
    .A2(_09219_),
    .B1(_10045_),
    .B2(_10060_),
    .X(_10061_));
 sky130_fd_sc_hd__inv_2 _13627_ (.A(_10061_),
    .Y(_01473_));
 sky130_fd_sc_hd__nand2_1 _13628_ (.A(_10001_),
    .B(net3731),
    .Y(_10062_));
 sky130_fd_sc_hd__a22o_1 _13629_ (.A1(_10053_),
    .A2(_09332_),
    .B1(_10045_),
    .B2(_10062_),
    .X(_10063_));
 sky130_fd_sc_hd__inv_2 _13630_ (.A(_10063_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor2_1 _13631_ (.A(_09230_),
    .B(_10047_),
    .Y(_10064_));
 sky130_fd_sc_hd__a31o_1 _13632_ (.A1(_10010_),
    .A2(net2132),
    .A3(_10046_),
    .B1(_10064_),
    .X(_01475_));
 sky130_fd_sc_hd__nor2_1 _13633_ (.A(_09233_),
    .B(_10047_),
    .Y(_10065_));
 sky130_fd_sc_hd__a31o_1 _13634_ (.A1(_10010_),
    .A2(net1417),
    .A3(_10046_),
    .B1(_10065_),
    .X(_01476_));
 sky130_fd_sc_hd__nor2_1 _13635_ (.A(_09236_),
    .B(_10047_),
    .Y(_10066_));
 sky130_fd_sc_hd__a31o_1 _13636_ (.A1(_10010_),
    .A2(net1129),
    .A3(_10047_),
    .B1(_10066_),
    .X(_01477_));
 sky130_fd_sc_hd__and3_1 _13637_ (.A(_10042_),
    .B(_09341_),
    .C(_10019_),
    .X(_10067_));
 sky130_fd_sc_hd__a31o_1 _13638_ (.A1(_10046_),
    .A2(_09977_),
    .A3(net1856),
    .B1(_10067_),
    .X(_01478_));
 sky130_fd_sc_hd__nor2_1 _13639_ (.A(_09243_),
    .B(_10047_),
    .Y(_10068_));
 sky130_fd_sc_hd__a31o_1 _13640_ (.A1(_10010_),
    .A2(net1331),
    .A3(_10047_),
    .B1(_10068_),
    .X(_01479_));
 sky130_fd_sc_hd__nor2_1 _13641_ (.A(_09246_),
    .B(_10047_),
    .Y(_10069_));
 sky130_fd_sc_hd__a31o_1 _13642_ (.A1(_10010_),
    .A2(net911),
    .A3(_10047_),
    .B1(_10069_),
    .X(_01464_));
 sky130_fd_sc_hd__and3_1 _13643_ (.A(_10042_),
    .B(_09345_),
    .C(_10019_),
    .X(_10070_));
 sky130_fd_sc_hd__a31o_1 _13644_ (.A1(_10046_),
    .A2(_09977_),
    .A3(net2025),
    .B1(_10070_),
    .X(_01465_));
 sky130_fd_sc_hd__nand2_1 _13645_ (.A(_10001_),
    .B(net2985),
    .Y(_10071_));
 sky130_fd_sc_hd__a22o_1 _13646_ (.A1(_10053_),
    .A2(_09348_),
    .B1(_10045_),
    .B2(_10071_),
    .X(_10072_));
 sky130_fd_sc_hd__inv_2 _13647_ (.A(_10072_),
    .Y(_01466_));
 sky130_fd_sc_hd__and3_1 _13648_ (.A(_10042_),
    .B(_09351_),
    .C(_10019_),
    .X(_10073_));
 sky130_fd_sc_hd__a31o_1 _13649_ (.A1(_10046_),
    .A2(_09977_),
    .A3(net2435),
    .B1(_10073_),
    .X(_01467_));
 sky130_fd_sc_hd__buf_4 _13650_ (.A(_09716_),
    .X(_10074_));
 sky130_fd_sc_hd__nand2_1 _13651_ (.A(_10074_),
    .B(net3676),
    .Y(_10075_));
 sky130_fd_sc_hd__a22o_1 _13652_ (.A1(_10053_),
    .A2(_09354_),
    .B1(_10045_),
    .B2(_10075_),
    .X(_10076_));
 sky130_fd_sc_hd__inv_2 _13653_ (.A(_10076_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _13654_ (.A(_10074_),
    .B(net3623),
    .Y(_10077_));
 sky130_fd_sc_hd__a22o_1 _13655_ (.A1(_10053_),
    .A2(_09263_),
    .B1(_10045_),
    .B2(_10077_),
    .X(_10078_));
 sky130_fd_sc_hd__inv_2 _13656_ (.A(_10078_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _13657_ (.A(_10074_),
    .B(net2914),
    .Y(_10079_));
 sky130_fd_sc_hd__a22o_1 _13658_ (.A1(_10053_),
    .A2(_09425_),
    .B1(_10045_),
    .B2(_10079_),
    .X(_10080_));
 sky130_fd_sc_hd__inv_2 _13659_ (.A(_10080_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _13660_ (.A(_10074_),
    .B(net3474),
    .Y(_10081_));
 sky130_fd_sc_hd__a22o_1 _13661_ (.A1(_10053_),
    .A2(_09269_),
    .B1(_10045_),
    .B2(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__inv_2 _13662_ (.A(_10082_),
    .Y(_01471_));
 sky130_fd_sc_hd__buf_4 _13663_ (.A(_09223_),
    .X(_10083_));
 sky130_fd_sc_hd__and3_1 _13664_ (.A(_10042_),
    .B(_09274_),
    .C(_10019_),
    .X(_10084_));
 sky130_fd_sc_hd__a31o_1 _13665_ (.A1(_10046_),
    .A2(_10083_),
    .A3(net2262),
    .B1(_10084_),
    .X(_01456_));
 sky130_fd_sc_hd__nand2_1 _13666_ (.A(_10074_),
    .B(net3939),
    .Y(_10085_));
 sky130_fd_sc_hd__a22o_1 _13667_ (.A1(_10053_),
    .A2(_09366_),
    .B1(_10045_),
    .B2(_10085_),
    .X(_10086_));
 sky130_fd_sc_hd__inv_2 _13668_ (.A(_10086_),
    .Y(_01457_));
 sky130_fd_sc_hd__and3_1 _13669_ (.A(_10042_),
    .B(_09369_),
    .C(_10019_),
    .X(_10087_));
 sky130_fd_sc_hd__a31o_1 _13670_ (.A1(_10046_),
    .A2(_10083_),
    .A3(net1287),
    .B1(_10087_),
    .X(_01458_));
 sky130_fd_sc_hd__nand2_1 _13671_ (.A(_10074_),
    .B(net3921),
    .Y(_10088_));
 sky130_fd_sc_hd__a22o_1 _13672_ (.A1(_10053_),
    .A2(_09284_),
    .B1(_10045_),
    .B2(_10088_),
    .X(_10089_));
 sky130_fd_sc_hd__inv_2 _13673_ (.A(_10089_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand2_1 _13674_ (.A(_10074_),
    .B(net3906),
    .Y(_10090_));
 sky130_fd_sc_hd__a22o_1 _13675_ (.A1(_10053_),
    .A2(_09288_),
    .B1(_10045_),
    .B2(_10090_),
    .X(_10091_));
 sky130_fd_sc_hd__inv_2 _13676_ (.A(_10091_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _13677_ (.A(_09733_),
    .B(net3782),
    .Y(_10092_));
 sky130_fd_sc_hd__o2bb2a_1 _13678_ (.A1_N(_10092_),
    .A2_N(_10046_),
    .B1(_09294_),
    .B2(_10043_),
    .X(_01461_));
 sky130_fd_sc_hd__nand2_1 _13679_ (.A(_09733_),
    .B(net3432),
    .Y(_10093_));
 sky130_fd_sc_hd__o2bb2a_1 _13680_ (.A1_N(_10093_),
    .A2_N(_10046_),
    .B1(_09298_),
    .B2(_10043_),
    .X(_01462_));
 sky130_fd_sc_hd__nor2_1 _13681_ (.A(_09300_),
    .B(_10047_),
    .Y(_10094_));
 sky130_fd_sc_hd__a31o_1 _13682_ (.A1(_10010_),
    .A2(net2618),
    .A3(_10047_),
    .B1(_10094_),
    .X(_01463_));
 sky130_fd_sc_hd__inv_2 _13683_ (.A(_09380_),
    .Y(_10095_));
 sky130_fd_sc_hd__or2_1 _13684_ (.A(_10095_),
    .B(_09983_),
    .X(_10096_));
 sky130_fd_sc_hd__nor2_2 _13685_ (.A(_09444_),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__inv_2 _13686_ (.A(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__nor2_4 _13687_ (.A(_08794_),
    .B(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__buf_4 _13688_ (.A(_10099_),
    .X(_10100_));
 sky130_fd_sc_hd__nor2_1 _13689_ (.A(_09625_),
    .B(_10098_),
    .Y(_10101_));
 sky130_fd_sc_hd__inv_2 _13690_ (.A(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__buf_4 _13691_ (.A(_10102_),
    .X(_10103_));
 sky130_fd_sc_hd__nand2_1 _13692_ (.A(_10074_),
    .B(net3026),
    .Y(_10104_));
 sky130_fd_sc_hd__a22o_1 _13693_ (.A1(_10100_),
    .A2(_09451_),
    .B1(_10103_),
    .B2(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__inv_2 _13694_ (.A(_10105_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _13695_ (.A(_10074_),
    .B(net3918),
    .Y(_10106_));
 sky130_fd_sc_hd__a22o_1 _13696_ (.A1(_10100_),
    .A2(_09315_),
    .B1(_10103_),
    .B2(_10106_),
    .X(_10107_));
 sky130_fd_sc_hd__inv_2 _13697_ (.A(_10107_),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_1 _13698_ (.A(_10074_),
    .B(net2898),
    .Y(_10108_));
 sky130_fd_sc_hd__a22o_1 _13699_ (.A1(_10100_),
    .A2(_09460_),
    .B1(_10103_),
    .B2(_10108_),
    .X(_10109_));
 sky130_fd_sc_hd__inv_2 _13700_ (.A(_10109_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand2_1 _13701_ (.A(_10074_),
    .B(net3894),
    .Y(_10110_));
 sky130_fd_sc_hd__a22o_1 _13702_ (.A1(_10100_),
    .A2(_09195_),
    .B1(_10103_),
    .B2(_10110_),
    .X(_10111_));
 sky130_fd_sc_hd__inv_2 _13703_ (.A(_10111_),
    .Y(_01451_));
 sky130_fd_sc_hd__nand2_1 _13704_ (.A(_10074_),
    .B(net3907),
    .Y(_10112_));
 sky130_fd_sc_hd__a22o_1 _13705_ (.A1(_10100_),
    .A2(_09201_),
    .B1(_10103_),
    .B2(_10112_),
    .X(_10113_));
 sky130_fd_sc_hd__inv_2 _13706_ (.A(_10113_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand2_1 _13707_ (.A(_10074_),
    .B(net2891),
    .Y(_10114_));
 sky130_fd_sc_hd__a22o_1 _13708_ (.A1(_10100_),
    .A2(_09205_),
    .B1(_10103_),
    .B2(_10114_),
    .X(_10115_));
 sky130_fd_sc_hd__inv_2 _13709_ (.A(_10115_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_1 _13710_ (.A(_10074_),
    .B(net2848),
    .Y(_10116_));
 sky130_fd_sc_hd__a22o_1 _13711_ (.A1(_10100_),
    .A2(_09398_),
    .B1(_10103_),
    .B2(_10116_),
    .X(_10117_));
 sky130_fd_sc_hd__inv_2 _13712_ (.A(_10117_),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_1 _13713_ (.A(_10074_),
    .B(net3893),
    .Y(_10118_));
 sky130_fd_sc_hd__a22o_1 _13714_ (.A1(_10100_),
    .A2(_09212_),
    .B1(_10103_),
    .B2(_10118_),
    .X(_10119_));
 sky130_fd_sc_hd__inv_2 _13715_ (.A(_10119_),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _13716_ (.A(_10074_),
    .B(net3097),
    .Y(_10120_));
 sky130_fd_sc_hd__a22o_1 _13717_ (.A1(_10100_),
    .A2(_09531_),
    .B1(_10103_),
    .B2(_10120_),
    .X(_10121_));
 sky130_fd_sc_hd__inv_2 _13718_ (.A(_10121_),
    .Y(_01440_));
 sky130_fd_sc_hd__buf_12 _13719_ (.A(net146),
    .X(_10122_));
 sky130_fd_sc_hd__buf_4 _13720_ (.A(_09716_),
    .X(_10123_));
 sky130_fd_sc_hd__nand2_1 _13721_ (.A(_10123_),
    .B(net3589),
    .Y(_10124_));
 sky130_fd_sc_hd__a22o_1 _13722_ (.A1(_10100_),
    .A2(_10122_),
    .B1(_10103_),
    .B2(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__inv_2 _13723_ (.A(_10125_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _13724_ (.A(_10123_),
    .B(net3027),
    .Y(_10126_));
 sky130_fd_sc_hd__a22o_1 _13725_ (.A1(_10100_),
    .A2(_09332_),
    .B1(_10103_),
    .B2(_10126_),
    .X(_10127_));
 sky130_fd_sc_hd__inv_2 _13726_ (.A(_10127_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _13727_ (.A(_10123_),
    .B(net3483),
    .Y(_10128_));
 sky130_fd_sc_hd__a22o_1 _13728_ (.A1(_10100_),
    .A2(_09589_),
    .B1(_10103_),
    .B2(_10128_),
    .X(_10129_));
 sky130_fd_sc_hd__inv_2 _13729_ (.A(_10129_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _13730_ (.A(_10123_),
    .B(net3030),
    .Y(_10130_));
 sky130_fd_sc_hd__a22o_1 _13731_ (.A1(_10100_),
    .A2(_09593_),
    .B1(_10103_),
    .B2(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__inv_2 _13732_ (.A(_10131_),
    .Y(_01444_));
 sky130_fd_sc_hd__buf_4 _13733_ (.A(_10102_),
    .X(_10132_));
 sky130_fd_sc_hd__nand2_1 _13734_ (.A(_10123_),
    .B(net3272),
    .Y(_10133_));
 sky130_fd_sc_hd__a22o_1 _13735_ (.A1(_10100_),
    .A2(_09338_),
    .B1(_10132_),
    .B2(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__inv_2 _13736_ (.A(_10134_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _13737_ (.A(_10123_),
    .B(net2963),
    .Y(_10135_));
 sky130_fd_sc_hd__a22o_1 _13738_ (.A1(_10100_),
    .A2(_09239_),
    .B1(_10132_),
    .B2(_10135_),
    .X(_10136_));
 sky130_fd_sc_hd__inv_2 _13739_ (.A(_10136_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand2_1 _13740_ (.A(_10123_),
    .B(net3095),
    .Y(_10137_));
 sky130_fd_sc_hd__a22o_1 _13741_ (.A1(_10100_),
    .A2(_09768_),
    .B1(_10132_),
    .B2(_10137_),
    .X(_10138_));
 sky130_fd_sc_hd__inv_2 _13742_ (.A(_10138_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _13743_ (.A(_10123_),
    .B(net3412),
    .Y(_10139_));
 sky130_fd_sc_hd__a22o_1 _13744_ (.A1(_10099_),
    .A2(_09415_),
    .B1(_10132_),
    .B2(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__inv_2 _13745_ (.A(_10140_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _13746_ (.A(_10123_),
    .B(net2944),
    .Y(_10141_));
 sky130_fd_sc_hd__a22o_1 _13747_ (.A1(_10099_),
    .A2(_09249_),
    .B1(_10132_),
    .B2(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__inv_2 _13748_ (.A(_10142_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _13749_ (.A(_10123_),
    .B(net3053),
    .Y(_10143_));
 sky130_fd_sc_hd__a22o_1 _13750_ (.A1(_10099_),
    .A2(_09348_),
    .B1(_10132_),
    .B2(_10143_),
    .X(_10144_));
 sky130_fd_sc_hd__inv_2 _13751_ (.A(_10144_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_1 _13752_ (.A(_10123_),
    .B(net3197),
    .Y(_10145_));
 sky130_fd_sc_hd__a22o_1 _13753_ (.A1(_10099_),
    .A2(_09256_),
    .B1(_10132_),
    .B2(_10145_),
    .X(_10146_));
 sky130_fd_sc_hd__inv_2 _13754_ (.A(_10146_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_1 _13755_ (.A(_10123_),
    .B(net3331),
    .Y(_10147_));
 sky130_fd_sc_hd__a22o_1 _13756_ (.A1(_10099_),
    .A2(_09354_),
    .B1(_10132_),
    .B2(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__inv_2 _13757_ (.A(_10148_),
    .Y(_01436_));
 sky130_fd_sc_hd__clkbuf_16 _13758_ (.A(net145),
    .X(_10149_));
 sky130_fd_sc_hd__nand2_1 _13759_ (.A(_10123_),
    .B(net3245),
    .Y(_10150_));
 sky130_fd_sc_hd__a22o_1 _13760_ (.A1(_10099_),
    .A2(_10149_),
    .B1(_10132_),
    .B2(_10150_),
    .X(_10151_));
 sky130_fd_sc_hd__inv_2 _13761_ (.A(_10151_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _13762_ (.A(_10123_),
    .B(net2875),
    .Y(_10152_));
 sky130_fd_sc_hd__a22o_1 _13763_ (.A1(_10099_),
    .A2(_09425_),
    .B1(_10132_),
    .B2(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__inv_2 _13764_ (.A(_10153_),
    .Y(_01438_));
 sky130_fd_sc_hd__clkbuf_16 _13765_ (.A(net144),
    .X(_10154_));
 sky130_fd_sc_hd__nand2_1 _13766_ (.A(_10123_),
    .B(net3124),
    .Y(_10155_));
 sky130_fd_sc_hd__a22o_1 _13767_ (.A1(_10099_),
    .A2(_10154_),
    .B1(_10132_),
    .B2(_10155_),
    .X(_10156_));
 sky130_fd_sc_hd__inv_2 _13768_ (.A(_10156_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_1 _13769_ (.A(_10123_),
    .B(net3485),
    .Y(_10157_));
 sky130_fd_sc_hd__a22o_1 _13770_ (.A1(_10099_),
    .A2(_09495_),
    .B1(_10132_),
    .B2(_10157_),
    .X(_10158_));
 sky130_fd_sc_hd__inv_2 _13771_ (.A(_10158_),
    .Y(_01424_));
 sky130_fd_sc_hd__buf_4 _13772_ (.A(_09716_),
    .X(_10159_));
 sky130_fd_sc_hd__nand2_1 _13773_ (.A(_10159_),
    .B(net2933),
    .Y(_10160_));
 sky130_fd_sc_hd__a22o_1 _13774_ (.A1(_10099_),
    .A2(_09366_),
    .B1(_10132_),
    .B2(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__inv_2 _13775_ (.A(_10161_),
    .Y(_01425_));
 sky130_fd_sc_hd__nand2_1 _13776_ (.A(_10159_),
    .B(net3137),
    .Y(_10162_));
 sky130_fd_sc_hd__a22o_1 _13777_ (.A1(_10099_),
    .A2(_09280_),
    .B1(_10132_),
    .B2(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__inv_2 _13778_ (.A(_10163_),
    .Y(_01426_));
 sky130_fd_sc_hd__clkbuf_16 _13779_ (.A(_09283_),
    .X(_10164_));
 sky130_fd_sc_hd__nand2_1 _13780_ (.A(_10159_),
    .B(net3624),
    .Y(_10165_));
 sky130_fd_sc_hd__a22o_1 _13781_ (.A1(_10099_),
    .A2(_10164_),
    .B1(_10132_),
    .B2(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__inv_2 _13782_ (.A(_10166_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _13783_ (.A(_10159_),
    .B(net2768),
    .Y(_10167_));
 sky130_fd_sc_hd__a22o_1 _13784_ (.A1(_10099_),
    .A2(_09288_),
    .B1(_10132_),
    .B2(_10167_),
    .X(_10168_));
 sky130_fd_sc_hd__inv_2 _13785_ (.A(_10168_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _13786_ (.A(_09733_),
    .B(net3062),
    .Y(_10169_));
 sky130_fd_sc_hd__o2bb2a_1 _13787_ (.A1_N(_10169_),
    .A2_N(_10103_),
    .B1(_09294_),
    .B2(_10098_),
    .X(_01429_));
 sky130_fd_sc_hd__nand2_1 _13788_ (.A(_09733_),
    .B(net3400),
    .Y(_10170_));
 sky130_fd_sc_hd__o2bb2a_1 _13789_ (.A1_N(_10170_),
    .A2_N(_10103_),
    .B1(_09298_),
    .B2(_10098_),
    .X(_01430_));
 sky130_fd_sc_hd__nand2_1 _13790_ (.A(_09733_),
    .B(net3358),
    .Y(_10171_));
 sky130_fd_sc_hd__o2bb2a_1 _13791_ (.A1_N(_10171_),
    .A2_N(_10103_),
    .B1(_09442_),
    .B2(_10098_),
    .X(_01431_));
 sky130_fd_sc_hd__inv_2 _13792_ (.A(_09445_),
    .Y(_10172_));
 sky130_fd_sc_hd__or2_2 _13793_ (.A(_10172_),
    .B(_09983_),
    .X(_10173_));
 sky130_fd_sc_hd__nor2_4 _13794_ (.A(_09444_),
    .B(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__inv_2 _13795_ (.A(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__nor2_1 _13796_ (.A(_09304_),
    .B(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__inv_2 _13797_ (.A(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__buf_4 _13798_ (.A(_10177_),
    .X(_10178_));
 sky130_fd_sc_hd__buf_4 _13799_ (.A(_10177_),
    .X(_10179_));
 sky130_fd_sc_hd__nor2_1 _13800_ (.A(_09181_),
    .B(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__a31o_1 _13801_ (.A1(_10010_),
    .A2(net901),
    .A3(_10178_),
    .B1(_10180_),
    .X(_01408_));
 sky130_fd_sc_hd__buf_4 _13802_ (.A(_09302_),
    .X(_10181_));
 sky130_fd_sc_hd__nor2_1 _13803_ (.A(_09185_),
    .B(_10179_),
    .Y(_10182_));
 sky130_fd_sc_hd__a31o_1 _13804_ (.A1(_10181_),
    .A2(net811),
    .A3(_10178_),
    .B1(_10182_),
    .X(_01409_));
 sky130_fd_sc_hd__nor2_4 _13805_ (.A(_09190_),
    .B(_10175_),
    .Y(_10183_));
 sky130_fd_sc_hd__nand2_1 _13806_ (.A(_10159_),
    .B(net2801),
    .Y(_10184_));
 sky130_fd_sc_hd__a22o_1 _13807_ (.A1(_10183_),
    .A2(_09460_),
    .B1(_10179_),
    .B2(_10184_),
    .X(_10185_));
 sky130_fd_sc_hd__inv_2 _13808_ (.A(_10185_),
    .Y(_01410_));
 sky130_fd_sc_hd__and3_1 _13809_ (.A(_10174_),
    .B(_09463_),
    .C(_10019_),
    .X(_10186_));
 sky130_fd_sc_hd__a31o_1 _13810_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net771),
    .B1(_10186_),
    .X(_01411_));
 sky130_fd_sc_hd__and3_1 _13811_ (.A(_10174_),
    .B(_09321_),
    .C(_10019_),
    .X(_10187_));
 sky130_fd_sc_hd__a31o_1 _13812_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net815),
    .B1(_10187_),
    .X(_01412_));
 sky130_fd_sc_hd__and3_1 _13813_ (.A(_10174_),
    .B(_09395_),
    .C(_10019_),
    .X(_10188_));
 sky130_fd_sc_hd__a31o_1 _13814_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net691),
    .B1(_10188_),
    .X(_01413_));
 sky130_fd_sc_hd__nor2_1 _13815_ (.A(_09209_),
    .B(_10179_),
    .Y(_10189_));
 sky130_fd_sc_hd__a31o_1 _13816_ (.A1(_10181_),
    .A2(net525),
    .A3(_10178_),
    .B1(_10189_),
    .X(_01414_));
 sky130_fd_sc_hd__nand2_1 _13817_ (.A(_10159_),
    .B(net2903),
    .Y(_10190_));
 sky130_fd_sc_hd__a22o_1 _13818_ (.A1(_10183_),
    .A2(_09212_),
    .B1(_10179_),
    .B2(_10190_),
    .X(_10191_));
 sky130_fd_sc_hd__inv_2 _13819_ (.A(_10191_),
    .Y(_01415_));
 sky130_fd_sc_hd__nor2_1 _13820_ (.A(_09216_),
    .B(_10179_),
    .Y(_10192_));
 sky130_fd_sc_hd__a31o_1 _13821_ (.A1(_10181_),
    .A2(net513),
    .A3(_10178_),
    .B1(_10192_),
    .X(_01400_));
 sky130_fd_sc_hd__nand2_1 _13822_ (.A(_10159_),
    .B(net2784),
    .Y(_10193_));
 sky130_fd_sc_hd__a22o_1 _13823_ (.A1(_10183_),
    .A2(_10122_),
    .B1(_10179_),
    .B2(_10193_),
    .X(_10194_));
 sky130_fd_sc_hd__inv_2 _13824_ (.A(_10194_),
    .Y(_01401_));
 sky130_fd_sc_hd__clkbuf_16 _13825_ (.A(_09331_),
    .X(_10195_));
 sky130_fd_sc_hd__nand2_1 _13826_ (.A(_10159_),
    .B(net3173),
    .Y(_10196_));
 sky130_fd_sc_hd__a22o_1 _13827_ (.A1(_10183_),
    .A2(_10195_),
    .B1(_10177_),
    .B2(_10196_),
    .X(_10197_));
 sky130_fd_sc_hd__inv_2 _13828_ (.A(_10197_),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_1 _13829_ (.A(_09230_),
    .B(_10179_),
    .Y(_10198_));
 sky130_fd_sc_hd__a31o_1 _13830_ (.A1(_10181_),
    .A2(net441),
    .A3(_10178_),
    .B1(_10198_),
    .X(_01403_));
 sky130_fd_sc_hd__nand2_1 _13831_ (.A(_10159_),
    .B(net2816),
    .Y(_10199_));
 sky130_fd_sc_hd__a22o_1 _13832_ (.A1(_10183_),
    .A2(_09593_),
    .B1(_10177_),
    .B2(_10199_),
    .X(_10200_));
 sky130_fd_sc_hd__inv_2 _13833_ (.A(_10200_),
    .Y(_01404_));
 sky130_fd_sc_hd__nor2_1 _13834_ (.A(_09236_),
    .B(_10179_),
    .Y(_10201_));
 sky130_fd_sc_hd__a31o_1 _13835_ (.A1(_10181_),
    .A2(net915),
    .A3(_10179_),
    .B1(_10201_),
    .X(_01405_));
 sky130_fd_sc_hd__buf_12 _13836_ (.A(_09238_),
    .X(_10202_));
 sky130_fd_sc_hd__nand2_1 _13837_ (.A(_10159_),
    .B(net3006),
    .Y(_10203_));
 sky130_fd_sc_hd__a22o_1 _13838_ (.A1(_10183_),
    .A2(_10202_),
    .B1(_10177_),
    .B2(_10203_),
    .X(_10204_));
 sky130_fd_sc_hd__inv_2 _13839_ (.A(_10204_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2_1 _13840_ (.A(_10159_),
    .B(net3349),
    .Y(_10205_));
 sky130_fd_sc_hd__a22o_1 _13841_ (.A1(_10183_),
    .A2(_09768_),
    .B1(_10177_),
    .B2(_10205_),
    .X(_10206_));
 sky130_fd_sc_hd__inv_2 _13842_ (.A(_10206_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _13843_ (.A(_09246_),
    .B(_10179_),
    .Y(_10207_));
 sky130_fd_sc_hd__a31o_1 _13844_ (.A1(_10181_),
    .A2(net1953),
    .A3(_10179_),
    .B1(_10207_),
    .X(_01392_));
 sky130_fd_sc_hd__and3_1 _13845_ (.A(_10174_),
    .B(_09345_),
    .C(_10019_),
    .X(_10208_));
 sky130_fd_sc_hd__a31o_1 _13846_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net1267),
    .B1(_10208_),
    .X(_01393_));
 sky130_fd_sc_hd__nor2_1 _13847_ (.A(_09253_),
    .B(_10179_),
    .Y(_10209_));
 sky130_fd_sc_hd__a31o_1 _13848_ (.A1(_10181_),
    .A2(net1830),
    .A3(_10179_),
    .B1(_10209_),
    .X(_01394_));
 sky130_fd_sc_hd__buf_4 _13849_ (.A(_09359_),
    .X(_10210_));
 sky130_fd_sc_hd__and3_1 _13850_ (.A(_10174_),
    .B(_09351_),
    .C(_10210_),
    .X(_10211_));
 sky130_fd_sc_hd__a31o_1 _13851_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net2390),
    .B1(_10211_),
    .X(_01395_));
 sky130_fd_sc_hd__nand2_1 _13852_ (.A(_10159_),
    .B(net3532),
    .Y(_10212_));
 sky130_fd_sc_hd__a22o_1 _13853_ (.A1(_10183_),
    .A2(_09354_),
    .B1(_10177_),
    .B2(_10212_),
    .X(_10213_));
 sky130_fd_sc_hd__inv_2 _13854_ (.A(_10213_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_1 _13855_ (.A(_10159_),
    .B(net3708),
    .Y(_10214_));
 sky130_fd_sc_hd__a22o_1 _13856_ (.A1(_10183_),
    .A2(_10149_),
    .B1(_10177_),
    .B2(_10214_),
    .X(_10215_));
 sky130_fd_sc_hd__inv_2 _13857_ (.A(_10215_),
    .Y(_01397_));
 sky130_fd_sc_hd__nand2_1 _13858_ (.A(_10159_),
    .B(net3023),
    .Y(_10216_));
 sky130_fd_sc_hd__a22o_1 _13859_ (.A1(_10183_),
    .A2(_09425_),
    .B1(_10177_),
    .B2(_10216_),
    .X(_10217_));
 sky130_fd_sc_hd__inv_2 _13860_ (.A(_10217_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand2_1 _13861_ (.A(_10159_),
    .B(net3324),
    .Y(_10218_));
 sky130_fd_sc_hd__a22o_1 _13862_ (.A1(_10183_),
    .A2(_10154_),
    .B1(_10177_),
    .B2(_10218_),
    .X(_10219_));
 sky130_fd_sc_hd__inv_2 _13863_ (.A(_10219_),
    .Y(_01399_));
 sky130_fd_sc_hd__and3_1 _13864_ (.A(_10174_),
    .B(_09274_),
    .C(_10210_),
    .X(_10220_));
 sky130_fd_sc_hd__a31o_1 _13865_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net1711),
    .B1(_10220_),
    .X(_01384_));
 sky130_fd_sc_hd__nor2_1 _13866_ (.A(_09277_),
    .B(_10179_),
    .Y(_10221_));
 sky130_fd_sc_hd__a31o_1 _13867_ (.A1(_10181_),
    .A2(net2465),
    .A3(_10179_),
    .B1(_10221_),
    .X(_01385_));
 sky130_fd_sc_hd__and3_1 _13868_ (.A(_10174_),
    .B(_09369_),
    .C(_10210_),
    .X(_10222_));
 sky130_fd_sc_hd__a31o_1 _13869_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net2420),
    .B1(_10222_),
    .X(_01386_));
 sky130_fd_sc_hd__nand2_1 _13870_ (.A(_10159_),
    .B(net4117),
    .Y(_10223_));
 sky130_fd_sc_hd__a22o_1 _13871_ (.A1(_10183_),
    .A2(_10164_),
    .B1(_10177_),
    .B2(_10223_),
    .X(_10224_));
 sky130_fd_sc_hd__inv_2 _13872_ (.A(_10224_),
    .Y(_01387_));
 sky130_fd_sc_hd__and3_1 _13873_ (.A(_10174_),
    .B(_09373_),
    .C(_10210_),
    .X(_10225_));
 sky130_fd_sc_hd__a31o_1 _13874_ (.A1(_10178_),
    .A2(_10083_),
    .A3(net1653),
    .B1(_10225_),
    .X(_01388_));
 sky130_fd_sc_hd__clkbuf_8 _13875_ (.A(_09375_),
    .X(_10226_));
 sky130_fd_sc_hd__nand2_1 _13876_ (.A(_10226_),
    .B(net3854),
    .Y(_10227_));
 sky130_fd_sc_hd__o2bb2a_1 _13877_ (.A1_N(_10227_),
    .A2_N(_10178_),
    .B1(_09294_),
    .B2(_10175_),
    .X(_01389_));
 sky130_fd_sc_hd__nand2_1 _13878_ (.A(_10226_),
    .B(net4119),
    .Y(_10228_));
 sky130_fd_sc_hd__o2bb2a_1 _13879_ (.A1_N(_10228_),
    .A2_N(_10178_),
    .B1(_09298_),
    .B2(_10175_),
    .X(_01390_));
 sky130_fd_sc_hd__nand2_1 _13880_ (.A(_10226_),
    .B(net4112),
    .Y(_10229_));
 sky130_fd_sc_hd__o2bb2a_1 _13881_ (.A1_N(_10229_),
    .A2_N(_10178_),
    .B1(_09442_),
    .B2(_10175_),
    .X(_01391_));
 sky130_fd_sc_hd__nand2_1 _13882_ (.A(_10226_),
    .B(net4293),
    .Y(_10230_));
 sky130_fd_sc_hd__nand2_1 _13883_ (.A(net2927),
    .B(net3899),
    .Y(_10231_));
 sky130_fd_sc_hd__nor2_1 _13884_ (.A(_09167_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__clkinv_4 _13885_ (.A(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__nor2_1 _13886_ (.A(_09172_),
    .B(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__nand2_2 _13887_ (.A(_10234_),
    .B(_09444_),
    .Y(_10235_));
 sky130_fd_sc_hd__or2_1 _13888_ (.A(_08727_),
    .B(_10235_),
    .X(_10236_));
 sky130_fd_sc_hd__clkbuf_4 _13889_ (.A(_10236_),
    .X(_10237_));
 sky130_fd_sc_hd__buf_4 _13890_ (.A(_10237_),
    .X(_10238_));
 sky130_fd_sc_hd__buf_12 _13891_ (.A(_09450_),
    .X(_10239_));
 sky130_fd_sc_hd__inv_2 _13892_ (.A(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__or2_1 _13893_ (.A(_08794_),
    .B(_10235_),
    .X(_10241_));
 sky130_fd_sc_hd__clkbuf_4 _13894_ (.A(_10241_),
    .X(_10242_));
 sky130_fd_sc_hd__o2bb2a_1 _13895_ (.A1_N(_10230_),
    .A2_N(_10238_),
    .B1(_10240_),
    .B2(_10242_),
    .X(_01376_));
 sky130_fd_sc_hd__buf_4 _13896_ (.A(_10237_),
    .X(_10243_));
 sky130_fd_sc_hd__nor2_1 _13897_ (.A(_09185_),
    .B(_10237_),
    .Y(_10244_));
 sky130_fd_sc_hd__a31o_1 _13898_ (.A1(_10181_),
    .A2(net2746),
    .A3(_10243_),
    .B1(_10244_),
    .X(_01377_));
 sky130_fd_sc_hd__nand2_1 _13899_ (.A(_09196_),
    .B(net2767),
    .Y(_10245_));
 sky130_fd_sc_hd__nand2_1 _13900_ (.A(_10238_),
    .B(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__o31a_1 _13901_ (.A1(_09193_),
    .A2(net68),
    .A3(_10242_),
    .B1(_10246_),
    .X(_01378_));
 sky130_fd_sc_hd__nor2_2 _13902_ (.A(_08728_),
    .B(_10235_),
    .Y(_10247_));
 sky130_fd_sc_hd__and2_1 _13903_ (.A(_10247_),
    .B(_09463_),
    .X(_10248_));
 sky130_fd_sc_hd__a31o_1 _13904_ (.A1(_10238_),
    .A2(_10083_),
    .A3(net2723),
    .B1(_10248_),
    .X(_01379_));
 sky130_fd_sc_hd__and2_1 _13905_ (.A(_10247_),
    .B(_09321_),
    .X(_10249_));
 sky130_fd_sc_hd__a31o_1 _13906_ (.A1(_10238_),
    .A2(_10083_),
    .A3(net2747),
    .B1(_10249_),
    .X(_01380_));
 sky130_fd_sc_hd__nand2_1 _13907_ (.A(_10226_),
    .B(net4309),
    .Y(_10250_));
 sky130_fd_sc_hd__inv_2 _13908_ (.A(_09204_),
    .Y(_10251_));
 sky130_fd_sc_hd__o2bb2a_1 _13909_ (.A1_N(_10250_),
    .A2_N(_10238_),
    .B1(_10251_),
    .B2(_10242_),
    .X(_01381_));
 sky130_fd_sc_hd__nand2_1 _13910_ (.A(_09196_),
    .B(net3928),
    .Y(_10252_));
 sky130_fd_sc_hd__nand2_1 _13911_ (.A(_10238_),
    .B(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__o31a_1 _13912_ (.A1(_09193_),
    .A2(net73),
    .A3(_10242_),
    .B1(_10253_),
    .X(_01382_));
 sky130_fd_sc_hd__and2_1 _13913_ (.A(_10247_),
    .B(_09326_),
    .X(_10254_));
 sky130_fd_sc_hd__a31o_1 _13914_ (.A1(_10243_),
    .A2(_10083_),
    .A3(net2736),
    .B1(_10254_),
    .X(_01383_));
 sky130_fd_sc_hd__nor2_1 _13915_ (.A(_09216_),
    .B(_10237_),
    .Y(_10255_));
 sky130_fd_sc_hd__a31o_1 _13916_ (.A1(_10181_),
    .A2(net665),
    .A3(_10243_),
    .B1(_10255_),
    .X(_01368_));
 sky130_fd_sc_hd__nand2_1 _13917_ (.A(_10226_),
    .B(net3649),
    .Y(_10256_));
 sky130_fd_sc_hd__inv_2 _13918_ (.A(net146),
    .Y(_10257_));
 sky130_fd_sc_hd__o2bb2a_1 _13919_ (.A1_N(_10256_),
    .A2_N(_10238_),
    .B1(_10257_),
    .B2(_10242_),
    .X(_01369_));
 sky130_fd_sc_hd__nand2_1 _13920_ (.A(_10226_),
    .B(net3707),
    .Y(_10258_));
 sky130_fd_sc_hd__inv_2 _13921_ (.A(_09331_),
    .Y(_10259_));
 sky130_fd_sc_hd__o2bb2a_1 _13922_ (.A1_N(_10258_),
    .A2_N(_10238_),
    .B1(_10259_),
    .B2(_10242_),
    .X(_01370_));
 sky130_fd_sc_hd__nor2_1 _13923_ (.A(_09230_),
    .B(_10237_),
    .Y(_10260_));
 sky130_fd_sc_hd__a31o_1 _13924_ (.A1(_10181_),
    .A2(net2550),
    .A3(_10243_),
    .B1(_10260_),
    .X(_01371_));
 sky130_fd_sc_hd__nor2_1 _13925_ (.A(_09233_),
    .B(_10237_),
    .Y(_10261_));
 sky130_fd_sc_hd__a31o_1 _13926_ (.A1(_10181_),
    .A2(net1755),
    .A3(_10243_),
    .B1(_10261_),
    .X(_01372_));
 sky130_fd_sc_hd__nor2_1 _13927_ (.A(_09236_),
    .B(_10237_),
    .Y(_10262_));
 sky130_fd_sc_hd__a31o_1 _13928_ (.A1(_10181_),
    .A2(net1023),
    .A3(_10243_),
    .B1(_10262_),
    .X(_01373_));
 sky130_fd_sc_hd__and2_1 _13929_ (.A(_10247_),
    .B(_09341_),
    .X(_10263_));
 sky130_fd_sc_hd__a31o_1 _13930_ (.A1(_10243_),
    .A2(_10083_),
    .A3(net2134),
    .B1(_10263_),
    .X(_01374_));
 sky130_fd_sc_hd__nor2_1 _13931_ (.A(_09243_),
    .B(_10237_),
    .Y(_10264_));
 sky130_fd_sc_hd__a31o_1 _13932_ (.A1(_10181_),
    .A2(net1993),
    .A3(_10243_),
    .B1(_10264_),
    .X(_01375_));
 sky130_fd_sc_hd__nor2_1 _13933_ (.A(_09246_),
    .B(_10237_),
    .Y(_10265_));
 sky130_fd_sc_hd__a31o_1 _13934_ (.A1(_10181_),
    .A2(net1225),
    .A3(_10243_),
    .B1(_10265_),
    .X(_01360_));
 sky130_fd_sc_hd__and2_1 _13935_ (.A(_10247_),
    .B(_09345_),
    .X(_10266_));
 sky130_fd_sc_hd__a31o_1 _13936_ (.A1(_10243_),
    .A2(_10083_),
    .A3(net2566),
    .B1(_10266_),
    .X(_01361_));
 sky130_fd_sc_hd__nand2_1 _13937_ (.A(_09196_),
    .B(net2740),
    .Y(_10267_));
 sky130_fd_sc_hd__nand2_1 _13938_ (.A(_10238_),
    .B(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__o31a_1 _13939_ (.A1(_09193_),
    .A2(net51),
    .A3(_10242_),
    .B1(_10268_),
    .X(_01362_));
 sky130_fd_sc_hd__nand2_1 _13940_ (.A(_09196_),
    .B(net2725),
    .Y(_10269_));
 sky130_fd_sc_hd__nand2_1 _13941_ (.A(_10238_),
    .B(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__o31a_1 _13942_ (.A1(_09193_),
    .A2(_09351_),
    .A3(_10242_),
    .B1(_10270_),
    .X(_01363_));
 sky130_fd_sc_hd__nor2_1 _13943_ (.A(_09260_),
    .B(_10237_),
    .Y(_10271_));
 sky130_fd_sc_hd__a31o_1 _13944_ (.A1(_10181_),
    .A2(net2468),
    .A3(_10243_),
    .B1(_10271_),
    .X(_01364_));
 sky130_fd_sc_hd__nand2_1 _13945_ (.A(_10226_),
    .B(net3615),
    .Y(_10272_));
 sky130_fd_sc_hd__inv_2 _13946_ (.A(net145),
    .Y(_10273_));
 sky130_fd_sc_hd__o2bb2a_1 _13947_ (.A1_N(_10272_),
    .A2_N(_10238_),
    .B1(_10273_),
    .B2(_10242_),
    .X(_01365_));
 sky130_fd_sc_hd__and2_1 _13948_ (.A(_10247_),
    .B(_09266_),
    .X(_10274_));
 sky130_fd_sc_hd__a31o_1 _13949_ (.A1(_10243_),
    .A2(_10083_),
    .A3(net2476),
    .B1(_10274_),
    .X(_01366_));
 sky130_fd_sc_hd__nand2_1 _13950_ (.A(_10226_),
    .B(net3681),
    .Y(_10275_));
 sky130_fd_sc_hd__inv_2 _13951_ (.A(net144),
    .Y(_10276_));
 sky130_fd_sc_hd__o2bb2a_1 _13952_ (.A1_N(_10275_),
    .A2_N(_10238_),
    .B1(_10276_),
    .B2(_10242_),
    .X(_01367_));
 sky130_fd_sc_hd__clkbuf_8 _13953_ (.A(_09223_),
    .X(_10277_));
 sky130_fd_sc_hd__and2_1 _13954_ (.A(_10247_),
    .B(_09274_),
    .X(_10278_));
 sky130_fd_sc_hd__a31o_1 _13955_ (.A1(_10243_),
    .A2(_10277_),
    .A3(net2546),
    .B1(_10278_),
    .X(_01352_));
 sky130_fd_sc_hd__buf_4 _13956_ (.A(_08776_),
    .X(_10279_));
 sky130_fd_sc_hd__clkbuf_8 _13957_ (.A(_10279_),
    .X(_10280_));
 sky130_fd_sc_hd__nor2_1 _13958_ (.A(_09277_),
    .B(_10237_),
    .Y(_10281_));
 sky130_fd_sc_hd__a31o_1 _13959_ (.A1(_10280_),
    .A2(net605),
    .A3(_10243_),
    .B1(_10281_),
    .X(_01353_));
 sky130_fd_sc_hd__nand2_1 _13960_ (.A(_09196_),
    .B(net2722),
    .Y(_10282_));
 sky130_fd_sc_hd__nand2_1 _13961_ (.A(_10238_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__o31a_1 _13962_ (.A1(_09193_),
    .A2(_09369_),
    .A3(_10242_),
    .B1(_10283_),
    .X(_01354_));
 sky130_fd_sc_hd__nand2_1 _13963_ (.A(_10226_),
    .B(net3647),
    .Y(_10284_));
 sky130_fd_sc_hd__inv_2 _13964_ (.A(_09283_),
    .Y(_10285_));
 sky130_fd_sc_hd__o2bb2a_1 _13965_ (.A1_N(_10284_),
    .A2_N(_10238_),
    .B1(_10285_),
    .B2(_10242_),
    .X(_01355_));
 sky130_fd_sc_hd__and2_1 _13966_ (.A(_10247_),
    .B(_09373_),
    .X(_10286_));
 sky130_fd_sc_hd__a31o_1 _13967_ (.A1(_10243_),
    .A2(_10277_),
    .A3(net2629),
    .B1(_10286_),
    .X(_01356_));
 sky130_fd_sc_hd__and2_1 _13968_ (.A(_10247_),
    .B(_09730_),
    .X(_10287_));
 sky130_fd_sc_hd__a31o_1 _13969_ (.A1(_10243_),
    .A2(_10277_),
    .A3(net2498),
    .B1(_10287_),
    .X(_01357_));
 sky130_fd_sc_hd__nand2_1 _13970_ (.A(_10226_),
    .B(net3957),
    .Y(_10288_));
 sky130_fd_sc_hd__buf_8 _13971_ (.A(_09297_),
    .X(_10289_));
 sky130_fd_sc_hd__o2bb2a_1 _13972_ (.A1_N(_10288_),
    .A2_N(_10238_),
    .B1(_10289_),
    .B2(_10235_),
    .X(_01358_));
 sky130_fd_sc_hd__nor2_1 _13973_ (.A(_09300_),
    .B(_10237_),
    .Y(_10290_));
 sky130_fd_sc_hd__a31o_1 _13974_ (.A1(_10280_),
    .A2(net2514),
    .A3(_10237_),
    .B1(_10290_),
    .X(_01359_));
 sky130_fd_sc_hd__nor2_8 _13975_ (.A(\line_cache_idx[8] ),
    .B(_10040_),
    .Y(_10291_));
 sky130_fd_sc_hd__clkinv_16 _13976_ (.A(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__nor2_4 _13977_ (.A(_10233_),
    .B(_10292_),
    .Y(_10293_));
 sky130_fd_sc_hd__nand2_4 _13978_ (.A(_10293_),
    .B(_09226_),
    .Y(_10294_));
 sky130_fd_sc_hd__nand2_1 _13979_ (.A(_08777_),
    .B(net4305),
    .Y(_10295_));
 sky130_fd_sc_hd__nand2_1 _13980_ (.A(_10293_),
    .B(_08778_),
    .Y(_10296_));
 sky130_fd_sc_hd__inv_2 _13981_ (.A(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__a22o_1 _13982_ (.A1(_10294_),
    .A2(_10295_),
    .B1(_10297_),
    .B2(_09451_),
    .X(_10298_));
 sky130_fd_sc_hd__inv_2 _13983_ (.A(_10298_),
    .Y(_01344_));
 sky130_fd_sc_hd__buf_4 _13984_ (.A(_10294_),
    .X(_10299_));
 sky130_fd_sc_hd__buf_4 _13985_ (.A(_10294_),
    .X(_10300_));
 sky130_fd_sc_hd__nor2_1 _13986_ (.A(_09185_),
    .B(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__a31o_1 _13987_ (.A1(_10280_),
    .A2(net1375),
    .A3(_10299_),
    .B1(_10301_),
    .X(_01345_));
 sky130_fd_sc_hd__nor2_1 _13988_ (.A(_09188_),
    .B(_10300_),
    .Y(_10302_));
 sky130_fd_sc_hd__a31o_1 _13989_ (.A1(_10280_),
    .A2(net2524),
    .A3(_10299_),
    .B1(_10302_),
    .X(_01346_));
 sky130_fd_sc_hd__and3_1 _13990_ (.A(_10293_),
    .B(_09463_),
    .C(_10210_),
    .X(_10303_));
 sky130_fd_sc_hd__a31o_1 _13991_ (.A1(_10280_),
    .A2(net2118),
    .A3(_10299_),
    .B1(_10303_),
    .X(_01347_));
 sky130_fd_sc_hd__and3_1 _13992_ (.A(_10293_),
    .B(_09321_),
    .C(_10210_),
    .X(_10304_));
 sky130_fd_sc_hd__a31o_1 _13993_ (.A1(_10280_),
    .A2(net2585),
    .A3(_10299_),
    .B1(_10304_),
    .X(_01348_));
 sky130_fd_sc_hd__and3_1 _13994_ (.A(_10293_),
    .B(_09395_),
    .C(_10210_),
    .X(_10305_));
 sky130_fd_sc_hd__a31o_1 _13995_ (.A1(_10280_),
    .A2(net2665),
    .A3(_10299_),
    .B1(_10305_),
    .X(_01349_));
 sky130_fd_sc_hd__nor2_1 _13996_ (.A(_09209_),
    .B(_10300_),
    .Y(_10306_));
 sky130_fd_sc_hd__a31o_1 _13997_ (.A1(_10280_),
    .A2(net2423),
    .A3(_10299_),
    .B1(_10306_),
    .X(_01350_));
 sky130_fd_sc_hd__and3_1 _13998_ (.A(_10293_),
    .B(_09326_),
    .C(_10210_),
    .X(_10307_));
 sky130_fd_sc_hd__a31o_1 _13999_ (.A1(_10280_),
    .A2(net1798),
    .A3(_10299_),
    .B1(_10307_),
    .X(_01351_));
 sky130_fd_sc_hd__nand2_1 _14000_ (.A(_08777_),
    .B(net4154),
    .Y(_10308_));
 sky130_fd_sc_hd__a22o_1 _14001_ (.A1(_10294_),
    .A2(_10308_),
    .B1(_10297_),
    .B2(_09531_),
    .X(_10309_));
 sky130_fd_sc_hd__inv_2 _14002_ (.A(_10309_),
    .Y(_01336_));
 sky130_fd_sc_hd__buf_8 _14003_ (.A(_08775_),
    .X(_10310_));
 sky130_fd_sc_hd__buf_4 _14004_ (.A(_10310_),
    .X(_10311_));
 sky130_fd_sc_hd__nand2_1 _14005_ (.A(_10311_),
    .B(net4218),
    .Y(_10312_));
 sky130_fd_sc_hd__buf_12 _14006_ (.A(net146),
    .X(_10313_));
 sky130_fd_sc_hd__a22o_1 _14007_ (.A1(_10294_),
    .A2(_10312_),
    .B1(_10297_),
    .B2(_10313_),
    .X(_10314_));
 sky130_fd_sc_hd__inv_2 _14008_ (.A(_10314_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _14009_ (.A(_10311_),
    .B(net4127),
    .Y(_10315_));
 sky130_fd_sc_hd__buf_12 _14010_ (.A(_09331_),
    .X(_10316_));
 sky130_fd_sc_hd__a22o_1 _14011_ (.A1(_10294_),
    .A2(_10315_),
    .B1(_10297_),
    .B2(_10316_),
    .X(_10317_));
 sky130_fd_sc_hd__inv_2 _14012_ (.A(_10317_),
    .Y(_01338_));
 sky130_fd_sc_hd__nor2_1 _14013_ (.A(_09230_),
    .B(_10300_),
    .Y(_10318_));
 sky130_fd_sc_hd__a31o_1 _14014_ (.A1(_10280_),
    .A2(net2345),
    .A3(_10299_),
    .B1(_10318_),
    .X(_01339_));
 sky130_fd_sc_hd__nor2_1 _14015_ (.A(_09233_),
    .B(_10300_),
    .Y(_10319_));
 sky130_fd_sc_hd__a31o_1 _14016_ (.A1(_10280_),
    .A2(net1866),
    .A3(_10299_),
    .B1(_10319_),
    .X(_01340_));
 sky130_fd_sc_hd__nor2_1 _14017_ (.A(_09236_),
    .B(_10300_),
    .Y(_10320_));
 sky130_fd_sc_hd__a31o_1 _14018_ (.A1(_10280_),
    .A2(net2022),
    .A3(_10299_),
    .B1(_10320_),
    .X(_01341_));
 sky130_fd_sc_hd__nand2_1 _14019_ (.A(_10311_),
    .B(net4238),
    .Y(_10321_));
 sky130_fd_sc_hd__a22o_1 _14020_ (.A1(_10294_),
    .A2(_10321_),
    .B1(_10297_),
    .B2(_09239_),
    .X(_10322_));
 sky130_fd_sc_hd__inv_2 _14021_ (.A(_10322_),
    .Y(_01342_));
 sky130_fd_sc_hd__nor2_1 _14022_ (.A(_09243_),
    .B(_10300_),
    .Y(_10323_));
 sky130_fd_sc_hd__a31o_1 _14023_ (.A1(_10280_),
    .A2(net1527),
    .A3(_10299_),
    .B1(_10323_),
    .X(_01343_));
 sky130_fd_sc_hd__nor2_1 _14024_ (.A(_09246_),
    .B(_10300_),
    .Y(_10324_));
 sky130_fd_sc_hd__a31o_1 _14025_ (.A1(_10280_),
    .A2(net2093),
    .A3(_10299_),
    .B1(_10324_),
    .X(_01320_));
 sky130_fd_sc_hd__and3_1 _14026_ (.A(_10293_),
    .B(_09345_),
    .C(_10210_),
    .X(_10325_));
 sky130_fd_sc_hd__a31o_1 _14027_ (.A1(_10280_),
    .A2(net1698),
    .A3(_10299_),
    .B1(_10325_),
    .X(_01321_));
 sky130_fd_sc_hd__nor2_1 _14028_ (.A(_09253_),
    .B(_10300_),
    .Y(_10326_));
 sky130_fd_sc_hd__a31o_1 _14029_ (.A1(_10280_),
    .A2(net1898),
    .A3(_10299_),
    .B1(_10326_),
    .X(_01322_));
 sky130_fd_sc_hd__buf_4 _14030_ (.A(_10279_),
    .X(_10327_));
 sky130_fd_sc_hd__and3_1 _14031_ (.A(_10293_),
    .B(_09351_),
    .C(_10210_),
    .X(_10328_));
 sky130_fd_sc_hd__a31o_1 _14032_ (.A1(_10327_),
    .A2(net1661),
    .A3(_10299_),
    .B1(_10328_),
    .X(_01323_));
 sky130_fd_sc_hd__nor2_1 _14033_ (.A(_09260_),
    .B(_10300_),
    .Y(_10329_));
 sky130_fd_sc_hd__a31o_1 _14034_ (.A1(_10327_),
    .A2(net1055),
    .A3(_10299_),
    .B1(_10329_),
    .X(_01324_));
 sky130_fd_sc_hd__nand2_1 _14035_ (.A(_10311_),
    .B(net4129),
    .Y(_10330_));
 sky130_fd_sc_hd__buf_12 _14036_ (.A(net145),
    .X(_10331_));
 sky130_fd_sc_hd__a22o_1 _14037_ (.A1(_10294_),
    .A2(_10330_),
    .B1(_10297_),
    .B2(_10331_),
    .X(_10332_));
 sky130_fd_sc_hd__inv_2 _14038_ (.A(_10332_),
    .Y(_01325_));
 sky130_fd_sc_hd__and3_1 _14039_ (.A(_10293_),
    .B(_09266_),
    .C(_10210_),
    .X(_10333_));
 sky130_fd_sc_hd__a31o_1 _14040_ (.A1(_10327_),
    .A2(net1441),
    .A3(_10300_),
    .B1(_10333_),
    .X(_01326_));
 sky130_fd_sc_hd__nand2_1 _14041_ (.A(_10311_),
    .B(net4232),
    .Y(_10334_));
 sky130_fd_sc_hd__buf_12 _14042_ (.A(net144),
    .X(_10335_));
 sky130_fd_sc_hd__a22o_1 _14043_ (.A1(_10294_),
    .A2(_10334_),
    .B1(_10297_),
    .B2(_10335_),
    .X(_10336_));
 sky130_fd_sc_hd__inv_2 _14044_ (.A(_10336_),
    .Y(_01327_));
 sky130_fd_sc_hd__nand2_1 _14045_ (.A(_10311_),
    .B(net4132),
    .Y(_10337_));
 sky130_fd_sc_hd__a22o_1 _14046_ (.A1(_10294_),
    .A2(_10337_),
    .B1(_10297_),
    .B2(_09495_),
    .X(_10338_));
 sky130_fd_sc_hd__inv_2 _14047_ (.A(_10338_),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _14048_ (.A(_09277_),
    .B(_10300_),
    .Y(_10339_));
 sky130_fd_sc_hd__a31o_1 _14049_ (.A1(_10327_),
    .A2(net2101),
    .A3(_10300_),
    .B1(_10339_),
    .X(_01313_));
 sky130_fd_sc_hd__and3_1 _14050_ (.A(_10293_),
    .B(_09369_),
    .C(_10210_),
    .X(_10340_));
 sky130_fd_sc_hd__a31o_1 _14051_ (.A1(_10327_),
    .A2(net2466),
    .A3(_10300_),
    .B1(_10340_),
    .X(_01314_));
 sky130_fd_sc_hd__nand2_1 _14052_ (.A(_10311_),
    .B(net4239),
    .Y(_10341_));
 sky130_fd_sc_hd__buf_12 _14053_ (.A(_09283_),
    .X(_10342_));
 sky130_fd_sc_hd__a22o_1 _14054_ (.A1(_10294_),
    .A2(_10341_),
    .B1(_10297_),
    .B2(_10342_),
    .X(_10343_));
 sky130_fd_sc_hd__inv_2 _14055_ (.A(_10343_),
    .Y(_01315_));
 sky130_fd_sc_hd__nand2_1 _14056_ (.A(_10311_),
    .B(net4143),
    .Y(_10344_));
 sky130_fd_sc_hd__a22o_1 _14057_ (.A1(_10294_),
    .A2(_10344_),
    .B1(_10297_),
    .B2(_09288_),
    .X(_10345_));
 sky130_fd_sc_hd__inv_2 _14058_ (.A(_10345_),
    .Y(_01316_));
 sky130_fd_sc_hd__nand2_1 _14059_ (.A(_10311_),
    .B(net3965),
    .Y(_10346_));
 sky130_fd_sc_hd__a22o_1 _14060_ (.A1(_10294_),
    .A2(_10346_),
    .B1(_10297_),
    .B2(net136),
    .X(_10347_));
 sky130_fd_sc_hd__inv_2 _14061_ (.A(_10347_),
    .Y(_01317_));
 sky130_fd_sc_hd__buf_12 _14062_ (.A(_09296_),
    .X(_10348_));
 sky130_fd_sc_hd__buf_4 _14063_ (.A(_08775_),
    .X(_10349_));
 sky130_fd_sc_hd__clkbuf_8 _14064_ (.A(_10349_),
    .X(_10350_));
 sky130_fd_sc_hd__nand2_1 _14065_ (.A(_10350_),
    .B(net3121),
    .Y(_10351_));
 sky130_fd_sc_hd__a22o_1 _14066_ (.A1(_10348_),
    .A2(_10293_),
    .B1(_10300_),
    .B2(_10351_),
    .X(_10352_));
 sky130_fd_sc_hd__inv_2 _14067_ (.A(_10352_),
    .Y(_01318_));
 sky130_fd_sc_hd__nand2_1 _14068_ (.A(_10350_),
    .B(net3021),
    .Y(_10353_));
 sky130_fd_sc_hd__a22o_1 _14069_ (.A1(net142),
    .A2(_10293_),
    .B1(_10300_),
    .B2(_10353_),
    .X(_10354_));
 sky130_fd_sc_hd__inv_2 _14070_ (.A(_10354_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_8 _14071_ (.A(\line_cache_idx[8] ),
    .B(_10095_),
    .Y(_10355_));
 sky130_fd_sc_hd__inv_16 _14072_ (.A(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__nor2_4 _14073_ (.A(_10233_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_4 _14074_ (.A(_10357_),
    .B(_09226_),
    .Y(_10358_));
 sky130_fd_sc_hd__buf_4 _14075_ (.A(_10358_),
    .X(_10359_));
 sky130_fd_sc_hd__buf_4 _14076_ (.A(_10358_),
    .X(_10360_));
 sky130_fd_sc_hd__nor2_1 _14077_ (.A(_09181_),
    .B(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__a31o_1 _14078_ (.A1(_10327_),
    .A2(net1401),
    .A3(_10359_),
    .B1(_10361_),
    .X(_01304_));
 sky130_fd_sc_hd__nor2_1 _14079_ (.A(_09185_),
    .B(_10360_),
    .Y(_10362_));
 sky130_fd_sc_hd__a31o_1 _14080_ (.A1(_10327_),
    .A2(net1449),
    .A3(_10359_),
    .B1(_10362_),
    .X(_01305_));
 sky130_fd_sc_hd__nor2_1 _14081_ (.A(_09188_),
    .B(_10360_),
    .Y(_10363_));
 sky130_fd_sc_hd__a31o_1 _14082_ (.A1(_10327_),
    .A2(net1926),
    .A3(_10359_),
    .B1(_10363_),
    .X(_01306_));
 sky130_fd_sc_hd__and3_1 _14083_ (.A(_10357_),
    .B(_09463_),
    .C(_10210_),
    .X(_10364_));
 sky130_fd_sc_hd__a31o_1 _14084_ (.A1(_10327_),
    .A2(net1700),
    .A3(_10359_),
    .B1(_10364_),
    .X(_01307_));
 sky130_fd_sc_hd__and3_1 _14085_ (.A(_10357_),
    .B(_09321_),
    .C(_10210_),
    .X(_10365_));
 sky130_fd_sc_hd__a31o_1 _14086_ (.A1(_10327_),
    .A2(net2377),
    .A3(_10359_),
    .B1(_10365_),
    .X(_01308_));
 sky130_fd_sc_hd__nand2_1 _14087_ (.A(_10311_),
    .B(net4109),
    .Y(_10366_));
 sky130_fd_sc_hd__nand2_1 _14088_ (.A(_10357_),
    .B(_08778_),
    .Y(_10367_));
 sky130_fd_sc_hd__inv_2 _14089_ (.A(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__a22o_1 _14090_ (.A1(_10358_),
    .A2(_10366_),
    .B1(_10368_),
    .B2(_09205_),
    .X(_10369_));
 sky130_fd_sc_hd__inv_2 _14091_ (.A(_10369_),
    .Y(_01309_));
 sky130_fd_sc_hd__nor2_1 _14092_ (.A(_09209_),
    .B(_10360_),
    .Y(_10370_));
 sky130_fd_sc_hd__a31o_1 _14093_ (.A1(_10327_),
    .A2(net797),
    .A3(_10359_),
    .B1(_10370_),
    .X(_01310_));
 sky130_fd_sc_hd__nand2_1 _14094_ (.A(_10311_),
    .B(net3950),
    .Y(_10371_));
 sky130_fd_sc_hd__a22o_1 _14095_ (.A1(_10358_),
    .A2(_10371_),
    .B1(_10368_),
    .B2(_09212_),
    .X(_10372_));
 sky130_fd_sc_hd__inv_2 _14096_ (.A(_10372_),
    .Y(_01311_));
 sky130_fd_sc_hd__nor2_1 _14097_ (.A(_09216_),
    .B(_10360_),
    .Y(_10373_));
 sky130_fd_sc_hd__a31o_1 _14098_ (.A1(_10327_),
    .A2(net935),
    .A3(_10359_),
    .B1(_10373_),
    .X(_01296_));
 sky130_fd_sc_hd__nand2_1 _14099_ (.A(_10311_),
    .B(net4199),
    .Y(_10374_));
 sky130_fd_sc_hd__a22o_1 _14100_ (.A1(_10358_),
    .A2(_10374_),
    .B1(_10368_),
    .B2(_10313_),
    .X(_10375_));
 sky130_fd_sc_hd__inv_2 _14101_ (.A(_10375_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _14102_ (.A(_10311_),
    .B(net4279),
    .Y(_10376_));
 sky130_fd_sc_hd__a22o_1 _14103_ (.A1(_10358_),
    .A2(_10376_),
    .B1(_10368_),
    .B2(_10316_),
    .X(_10377_));
 sky130_fd_sc_hd__inv_2 _14104_ (.A(_10377_),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _14105_ (.A(_10311_),
    .B(net4226),
    .Y(_10378_));
 sky130_fd_sc_hd__a22o_1 _14106_ (.A1(_10358_),
    .A2(_10378_),
    .B1(_10368_),
    .B2(_09589_),
    .X(_10379_));
 sky130_fd_sc_hd__inv_2 _14107_ (.A(_10379_),
    .Y(_01299_));
 sky130_fd_sc_hd__nor2_1 _14108_ (.A(_09233_),
    .B(_10360_),
    .Y(_10380_));
 sky130_fd_sc_hd__a31o_1 _14109_ (.A1(_10327_),
    .A2(net1239),
    .A3(_10359_),
    .B1(_10380_),
    .X(_01300_));
 sky130_fd_sc_hd__nor2_1 _14110_ (.A(_09236_),
    .B(_10360_),
    .Y(_10381_));
 sky130_fd_sc_hd__a31o_1 _14111_ (.A1(_10327_),
    .A2(net1011),
    .A3(_10359_),
    .B1(_10381_),
    .X(_01301_));
 sky130_fd_sc_hd__and3_1 _14112_ (.A(_10357_),
    .B(_09341_),
    .C(_10210_),
    .X(_10382_));
 sky130_fd_sc_hd__a31o_1 _14113_ (.A1(_10327_),
    .A2(net1195),
    .A3(_10359_),
    .B1(_10382_),
    .X(_01302_));
 sky130_fd_sc_hd__nor2_1 _14114_ (.A(_09243_),
    .B(_10360_),
    .Y(_10383_));
 sky130_fd_sc_hd__a31o_1 _14115_ (.A1(_10327_),
    .A2(net885),
    .A3(_10359_),
    .B1(_10383_),
    .X(_01303_));
 sky130_fd_sc_hd__nand2_1 _14116_ (.A(_10311_),
    .B(net3992),
    .Y(_10384_));
 sky130_fd_sc_hd__a22o_1 _14117_ (.A1(_10358_),
    .A2(_10384_),
    .B1(_10368_),
    .B2(_09415_),
    .X(_10385_));
 sky130_fd_sc_hd__inv_2 _14118_ (.A(_10385_),
    .Y(_01288_));
 sky130_fd_sc_hd__buf_4 _14119_ (.A(_10279_),
    .X(_10386_));
 sky130_fd_sc_hd__and3_1 _14120_ (.A(_10357_),
    .B(_09345_),
    .C(_10210_),
    .X(_10387_));
 sky130_fd_sc_hd__a31o_1 _14121_ (.A1(_10386_),
    .A2(net2173),
    .A3(_10359_),
    .B1(_10387_),
    .X(_01289_));
 sky130_fd_sc_hd__nor2_1 _14122_ (.A(_09253_),
    .B(_10360_),
    .Y(_10388_));
 sky130_fd_sc_hd__a31o_1 _14123_ (.A1(_10386_),
    .A2(net1113),
    .A3(_10359_),
    .B1(_10388_),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_4 _14124_ (.A(_09359_),
    .X(_10389_));
 sky130_fd_sc_hd__and3_1 _14125_ (.A(_10357_),
    .B(_09351_),
    .C(_10389_),
    .X(_10390_));
 sky130_fd_sc_hd__a31o_1 _14126_ (.A1(_10386_),
    .A2(net825),
    .A3(_10359_),
    .B1(_10390_),
    .X(_01291_));
 sky130_fd_sc_hd__nor2_1 _14127_ (.A(_09260_),
    .B(_10360_),
    .Y(_10391_));
 sky130_fd_sc_hd__a31o_1 _14128_ (.A1(_10386_),
    .A2(net1145),
    .A3(_10359_),
    .B1(_10391_),
    .X(_01292_));
 sky130_fd_sc_hd__nand2_1 _14129_ (.A(_10311_),
    .B(net4231),
    .Y(_10392_));
 sky130_fd_sc_hd__a22o_1 _14130_ (.A1(_10358_),
    .A2(_10392_),
    .B1(_10368_),
    .B2(_10331_),
    .X(_10393_));
 sky130_fd_sc_hd__inv_2 _14131_ (.A(_10393_),
    .Y(_01293_));
 sky130_fd_sc_hd__and3_1 _14132_ (.A(_10357_),
    .B(_09266_),
    .C(_10389_),
    .X(_10394_));
 sky130_fd_sc_hd__a31o_1 _14133_ (.A1(_10386_),
    .A2(net1353),
    .A3(_10359_),
    .B1(_10394_),
    .X(_01294_));
 sky130_fd_sc_hd__clkbuf_8 _14134_ (.A(_10310_),
    .X(_10395_));
 sky130_fd_sc_hd__nand2_1 _14135_ (.A(_10395_),
    .B(net4240),
    .Y(_10396_));
 sky130_fd_sc_hd__a22o_1 _14136_ (.A1(_10358_),
    .A2(_10396_),
    .B1(_10368_),
    .B2(_10335_),
    .X(_10397_));
 sky130_fd_sc_hd__inv_2 _14137_ (.A(_10397_),
    .Y(_01295_));
 sky130_fd_sc_hd__and3_1 _14138_ (.A(_10357_),
    .B(_09274_),
    .C(_10389_),
    .X(_10398_));
 sky130_fd_sc_hd__a31o_1 _14139_ (.A1(_10386_),
    .A2(net705),
    .A3(_10360_),
    .B1(_10398_),
    .X(_01280_));
 sky130_fd_sc_hd__nand2_1 _14140_ (.A(_10395_),
    .B(net3913),
    .Y(_10399_));
 sky130_fd_sc_hd__a22o_1 _14141_ (.A1(_10358_),
    .A2(_10399_),
    .B1(_10368_),
    .B2(_09366_),
    .X(_10400_));
 sky130_fd_sc_hd__inv_2 _14142_ (.A(_10400_),
    .Y(_01281_));
 sky130_fd_sc_hd__and3_1 _14143_ (.A(_10357_),
    .B(_09369_),
    .C(_10389_),
    .X(_10401_));
 sky130_fd_sc_hd__a31o_1 _14144_ (.A1(_10386_),
    .A2(net1051),
    .A3(_10360_),
    .B1(_10401_),
    .X(_01282_));
 sky130_fd_sc_hd__nand2_1 _14145_ (.A(_10395_),
    .B(net4131),
    .Y(_10402_));
 sky130_fd_sc_hd__a22o_1 _14146_ (.A1(_10358_),
    .A2(_10402_),
    .B1(_10368_),
    .B2(_10342_),
    .X(_10403_));
 sky130_fd_sc_hd__inv_2 _14147_ (.A(_10403_),
    .Y(_01283_));
 sky130_fd_sc_hd__and3_1 _14148_ (.A(_10357_),
    .B(_09373_),
    .C(_10389_),
    .X(_10404_));
 sky130_fd_sc_hd__a31o_1 _14149_ (.A1(_10386_),
    .A2(net733),
    .A3(_10360_),
    .B1(_10404_),
    .X(_01284_));
 sky130_fd_sc_hd__and3_1 _14150_ (.A(_10357_),
    .B(_09730_),
    .C(_10389_),
    .X(_10405_));
 sky130_fd_sc_hd__a31o_1 _14151_ (.A1(_10386_),
    .A2(net681),
    .A3(_10360_),
    .B1(_10405_),
    .X(_01285_));
 sky130_fd_sc_hd__nand2_1 _14152_ (.A(_10350_),
    .B(net3148),
    .Y(_10406_));
 sky130_fd_sc_hd__a22o_1 _14153_ (.A1(_10348_),
    .A2(_10357_),
    .B1(_10360_),
    .B2(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__inv_2 _14154_ (.A(_10407_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _14155_ (.A(_10350_),
    .B(net2947),
    .Y(_10408_));
 sky130_fd_sc_hd__a22o_1 _14156_ (.A1(net142),
    .A2(_10357_),
    .B1(_10360_),
    .B2(_10408_),
    .X(_10409_));
 sky130_fd_sc_hd__inv_2 _14157_ (.A(_10409_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_4 _14158_ (.A(\line_cache_idx[8] ),
    .B(_10172_),
    .Y(_10410_));
 sky130_fd_sc_hd__clkinv_16 _14159_ (.A(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__nor2_4 _14160_ (.A(_10233_),
    .B(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__buf_12 _14161_ (.A(_09225_),
    .X(_10413_));
 sky130_fd_sc_hd__nand2_4 _14162_ (.A(_10412_),
    .B(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__buf_4 _14163_ (.A(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__nand2_1 _14164_ (.A(_10395_),
    .B(net3979),
    .Y(_10416_));
 sky130_fd_sc_hd__nand2_1 _14165_ (.A(_10412_),
    .B(_08778_),
    .Y(_10417_));
 sky130_fd_sc_hd__inv_2 _14166_ (.A(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__a22o_1 _14167_ (.A1(_10415_),
    .A2(_10416_),
    .B1(_10418_),
    .B2(_09451_),
    .X(_10419_));
 sky130_fd_sc_hd__inv_2 _14168_ (.A(_10419_),
    .Y(_01272_));
 sky130_fd_sc_hd__buf_4 _14169_ (.A(_10414_),
    .X(_10420_));
 sky130_fd_sc_hd__nor2_1 _14170_ (.A(_09185_),
    .B(_10415_),
    .Y(_10421_));
 sky130_fd_sc_hd__a31o_1 _14171_ (.A1(_10386_),
    .A2(net469),
    .A3(_10420_),
    .B1(_10421_),
    .X(_01273_));
 sky130_fd_sc_hd__nor2_1 _14172_ (.A(_09188_),
    .B(_10415_),
    .Y(_10422_));
 sky130_fd_sc_hd__a31o_1 _14173_ (.A1(_10386_),
    .A2(net417),
    .A3(_10420_),
    .B1(_10422_),
    .X(_01274_));
 sky130_fd_sc_hd__nand2_1 _14174_ (.A(_10395_),
    .B(net3963),
    .Y(_10423_));
 sky130_fd_sc_hd__a22o_1 _14175_ (.A1(_10415_),
    .A2(_10423_),
    .B1(_10418_),
    .B2(_09195_),
    .X(_10424_));
 sky130_fd_sc_hd__inv_2 _14176_ (.A(_10424_),
    .Y(_01275_));
 sky130_fd_sc_hd__and3_1 _14177_ (.A(_10412_),
    .B(_09321_),
    .C(_10389_),
    .X(_10425_));
 sky130_fd_sc_hd__a31o_1 _14178_ (.A1(_10386_),
    .A2(net501),
    .A3(_10420_),
    .B1(_10425_),
    .X(_01276_));
 sky130_fd_sc_hd__and3_1 _14179_ (.A(_10412_),
    .B(_09395_),
    .C(_10389_),
    .X(_10426_));
 sky130_fd_sc_hd__a31o_1 _14180_ (.A1(_10386_),
    .A2(net427),
    .A3(_10420_),
    .B1(_10426_),
    .X(_01277_));
 sky130_fd_sc_hd__nor2_1 _14181_ (.A(_09209_),
    .B(_10415_),
    .Y(_10427_));
 sky130_fd_sc_hd__a31o_1 _14182_ (.A1(_10386_),
    .A2(net457),
    .A3(_10420_),
    .B1(_10427_),
    .X(_01278_));
 sky130_fd_sc_hd__and3_1 _14183_ (.A(_10412_),
    .B(_09326_),
    .C(_10389_),
    .X(_10428_));
 sky130_fd_sc_hd__a31o_1 _14184_ (.A1(_10386_),
    .A2(net527),
    .A3(_10420_),
    .B1(_10428_),
    .X(_01279_));
 sky130_fd_sc_hd__nor2_1 _14185_ (.A(_09216_),
    .B(_10415_),
    .Y(_10429_));
 sky130_fd_sc_hd__a31o_1 _14186_ (.A1(_10386_),
    .A2(net549),
    .A3(_10420_),
    .B1(_10429_),
    .X(_01264_));
 sky130_fd_sc_hd__nand2_1 _14187_ (.A(_10395_),
    .B(net3953),
    .Y(_10430_));
 sky130_fd_sc_hd__a22o_1 _14188_ (.A1(_10414_),
    .A2(_10430_),
    .B1(_10418_),
    .B2(_10313_),
    .X(_10431_));
 sky130_fd_sc_hd__inv_2 _14189_ (.A(_10431_),
    .Y(_01265_));
 sky130_fd_sc_hd__nand2_1 _14190_ (.A(_10395_),
    .B(net4032),
    .Y(_10432_));
 sky130_fd_sc_hd__a22o_1 _14191_ (.A1(_10414_),
    .A2(_10432_),
    .B1(_10418_),
    .B2(_10316_),
    .X(_10433_));
 sky130_fd_sc_hd__inv_2 _14192_ (.A(_10433_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _14193_ (.A(_10395_),
    .B(net4028),
    .Y(_10434_));
 sky130_fd_sc_hd__a22o_1 _14194_ (.A1(_10414_),
    .A2(_10434_),
    .B1(_10418_),
    .B2(_09589_),
    .X(_10435_));
 sky130_fd_sc_hd__inv_2 _14195_ (.A(_10435_),
    .Y(_01267_));
 sky130_fd_sc_hd__buf_4 _14196_ (.A(_10279_),
    .X(_10436_));
 sky130_fd_sc_hd__nor2_1 _14197_ (.A(_09233_),
    .B(_10415_),
    .Y(_10437_));
 sky130_fd_sc_hd__a31o_1 _14198_ (.A1(_10436_),
    .A2(net453),
    .A3(_10420_),
    .B1(_10437_),
    .X(_01268_));
 sky130_fd_sc_hd__nor2_1 _14199_ (.A(_09236_),
    .B(_10415_),
    .Y(_10438_));
 sky130_fd_sc_hd__a31o_1 _14200_ (.A1(_10436_),
    .A2(net535),
    .A3(_10420_),
    .B1(_10438_),
    .X(_01269_));
 sky130_fd_sc_hd__nand2_1 _14201_ (.A(_10395_),
    .B(net3991),
    .Y(_10439_));
 sky130_fd_sc_hd__a22o_1 _14202_ (.A1(_10414_),
    .A2(_10439_),
    .B1(_10418_),
    .B2(_09239_),
    .X(_10440_));
 sky130_fd_sc_hd__inv_2 _14203_ (.A(_10440_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _14204_ (.A(_09243_),
    .B(_10415_),
    .Y(_10441_));
 sky130_fd_sc_hd__a31o_1 _14205_ (.A1(_10436_),
    .A2(net447),
    .A3(_10420_),
    .B1(_10441_),
    .X(_01271_));
 sky130_fd_sc_hd__nor2_1 _14206_ (.A(_09246_),
    .B(_10415_),
    .Y(_10442_));
 sky130_fd_sc_hd__a31o_1 _14207_ (.A1(_10436_),
    .A2(net523),
    .A3(_10420_),
    .B1(_10442_),
    .X(_01256_));
 sky130_fd_sc_hd__and3_1 _14208_ (.A(_10412_),
    .B(_09345_),
    .C(_10389_),
    .X(_10443_));
 sky130_fd_sc_hd__a31o_1 _14209_ (.A1(_10436_),
    .A2(net541),
    .A3(_10420_),
    .B1(_10443_),
    .X(_01257_));
 sky130_fd_sc_hd__nand2_1 _14210_ (.A(_10395_),
    .B(net4153),
    .Y(_10444_));
 sky130_fd_sc_hd__a22o_1 _14211_ (.A1(_10414_),
    .A2(_10444_),
    .B1(_10418_),
    .B2(_09348_),
    .X(_10445_));
 sky130_fd_sc_hd__inv_2 _14212_ (.A(_10445_),
    .Y(_01258_));
 sky130_fd_sc_hd__and3_1 _14213_ (.A(_10412_),
    .B(_09351_),
    .C(_10389_),
    .X(_10446_));
 sky130_fd_sc_hd__a31o_1 _14214_ (.A1(_10436_),
    .A2(net591),
    .A3(_10420_),
    .B1(_10446_),
    .X(_01259_));
 sky130_fd_sc_hd__nand2_1 _14215_ (.A(_10395_),
    .B(net4201),
    .Y(_10447_));
 sky130_fd_sc_hd__a22o_1 _14216_ (.A1(_10414_),
    .A2(_10447_),
    .B1(_10418_),
    .B2(_09354_),
    .X(_10448_));
 sky130_fd_sc_hd__inv_2 _14217_ (.A(_10448_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_1 _14218_ (.A(_10395_),
    .B(net4142),
    .Y(_10449_));
 sky130_fd_sc_hd__a22o_1 _14219_ (.A1(_10414_),
    .A2(_10449_),
    .B1(_10418_),
    .B2(_10331_),
    .X(_10450_));
 sky130_fd_sc_hd__inv_2 _14220_ (.A(_10450_),
    .Y(_01261_));
 sky130_fd_sc_hd__and3_1 _14221_ (.A(_10412_),
    .B(_09266_),
    .C(_10389_),
    .X(_10451_));
 sky130_fd_sc_hd__a31o_1 _14222_ (.A1(_10436_),
    .A2(net479),
    .A3(_10420_),
    .B1(_10451_),
    .X(_01262_));
 sky130_fd_sc_hd__nand2_1 _14223_ (.A(_10395_),
    .B(net3930),
    .Y(_10452_));
 sky130_fd_sc_hd__a22o_1 _14224_ (.A1(_10414_),
    .A2(_10452_),
    .B1(_10418_),
    .B2(_10335_),
    .X(_10453_));
 sky130_fd_sc_hd__inv_2 _14225_ (.A(_10453_),
    .Y(_01263_));
 sky130_fd_sc_hd__and3_1 _14226_ (.A(_10412_),
    .B(_09274_),
    .C(_10389_),
    .X(_10454_));
 sky130_fd_sc_hd__a31o_1 _14227_ (.A1(_10436_),
    .A2(net1706),
    .A3(_10420_),
    .B1(_10454_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_1 _14228_ (.A(_09277_),
    .B(_10415_),
    .Y(_10455_));
 sky130_fd_sc_hd__a31o_1 _14229_ (.A1(_10436_),
    .A2(net1945),
    .A3(_10420_),
    .B1(_10455_),
    .X(_01249_));
 sky130_fd_sc_hd__and3_1 _14230_ (.A(_10412_),
    .B(_09369_),
    .C(_10389_),
    .X(_10456_));
 sky130_fd_sc_hd__a31o_1 _14231_ (.A1(_10436_),
    .A2(net1523),
    .A3(_10415_),
    .B1(_10456_),
    .X(_01250_));
 sky130_fd_sc_hd__nand2_1 _14232_ (.A(_10395_),
    .B(net4025),
    .Y(_10457_));
 sky130_fd_sc_hd__a22o_1 _14233_ (.A1(_10414_),
    .A2(_10457_),
    .B1(_10418_),
    .B2(_10342_),
    .X(_10458_));
 sky130_fd_sc_hd__inv_2 _14234_ (.A(_10458_),
    .Y(_01251_));
 sky130_fd_sc_hd__and3_1 _14235_ (.A(_10412_),
    .B(_09373_),
    .C(_10389_),
    .X(_10459_));
 sky130_fd_sc_hd__a31o_1 _14236_ (.A1(_10436_),
    .A2(net659),
    .A3(_10415_),
    .B1(_10459_),
    .X(_01252_));
 sky130_fd_sc_hd__and3_1 _14237_ (.A(_10412_),
    .B(_09730_),
    .C(_10389_),
    .X(_10460_));
 sky130_fd_sc_hd__a31o_1 _14238_ (.A1(_10436_),
    .A2(net837),
    .A3(_10415_),
    .B1(_10460_),
    .X(_01253_));
 sky130_fd_sc_hd__nand2_1 _14239_ (.A(_10350_),
    .B(net2941),
    .Y(_10461_));
 sky130_fd_sc_hd__a22o_1 _14240_ (.A1(_10348_),
    .A2(_10412_),
    .B1(_10415_),
    .B2(_10461_),
    .X(_10462_));
 sky130_fd_sc_hd__inv_2 _14241_ (.A(_10462_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand2_1 _14242_ (.A(_10350_),
    .B(net3000),
    .Y(_10463_));
 sky130_fd_sc_hd__a22o_1 _14243_ (.A1(net142),
    .A2(_10412_),
    .B1(_10415_),
    .B2(_10463_),
    .X(_10464_));
 sky130_fd_sc_hd__inv_2 _14244_ (.A(_10464_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2_1 _14245_ (.A(_10226_),
    .B(net3656),
    .Y(_10465_));
 sky130_fd_sc_hd__inv_4 _14246_ (.A(_10231_),
    .Y(_10466_));
 sky130_fd_sc_hd__nand2_4 _14247_ (.A(_09509_),
    .B(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__nor2_4 _14248_ (.A(\line_cache_idx[8] ),
    .B(_09172_),
    .Y(_10468_));
 sky130_fd_sc_hd__inv_16 _14249_ (.A(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__nor2_4 _14250_ (.A(_10467_),
    .B(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__nand2_4 _14251_ (.A(_10470_),
    .B(_09226_),
    .Y(_10471_));
 sky130_fd_sc_hd__clkbuf_4 _14252_ (.A(_10471_),
    .X(_10472_));
 sky130_fd_sc_hd__nand2_4 _14253_ (.A(_10470_),
    .B(_08778_),
    .Y(_10473_));
 sky130_fd_sc_hd__o2bb2a_1 _14254_ (.A1_N(_10465_),
    .A2_N(_10472_),
    .B1(_10240_),
    .B2(_10473_),
    .X(_01232_));
 sky130_fd_sc_hd__nand2_1 _14255_ (.A(_10226_),
    .B(net3618),
    .Y(_10474_));
 sky130_fd_sc_hd__inv_2 _14256_ (.A(_09314_),
    .Y(_10475_));
 sky130_fd_sc_hd__o2bb2a_1 _14257_ (.A1_N(_10474_),
    .A2_N(_10472_),
    .B1(_10475_),
    .B2(_10473_),
    .X(_01233_));
 sky130_fd_sc_hd__buf_4 _14258_ (.A(_10471_),
    .X(_10476_));
 sky130_fd_sc_hd__nor2_1 _14259_ (.A(_09188_),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__a31o_1 _14260_ (.A1(_10436_),
    .A2(net569),
    .A3(_10472_),
    .B1(_10477_),
    .X(_01234_));
 sky130_fd_sc_hd__nand2_1 _14261_ (.A(_10226_),
    .B(net3408),
    .Y(_10478_));
 sky130_fd_sc_hd__inv_2 _14262_ (.A(_09194_),
    .Y(_10479_));
 sky130_fd_sc_hd__o2bb2a_1 _14263_ (.A1_N(_10478_),
    .A2_N(_10472_),
    .B1(_10479_),
    .B2(_10473_),
    .X(_01235_));
 sky130_fd_sc_hd__buf_4 _14264_ (.A(_09359_),
    .X(_10480_));
 sky130_fd_sc_hd__and3_1 _14265_ (.A(_10470_),
    .B(_09321_),
    .C(_10480_),
    .X(_10481_));
 sky130_fd_sc_hd__a31o_1 _14266_ (.A1(_10436_),
    .A2(net543),
    .A3(_10472_),
    .B1(_10481_),
    .X(_01236_));
 sky130_fd_sc_hd__nand2_1 _14267_ (.A(_10226_),
    .B(net3214),
    .Y(_10482_));
 sky130_fd_sc_hd__o2bb2a_1 _14268_ (.A1_N(_10482_),
    .A2_N(_10472_),
    .B1(_10251_),
    .B2(_10473_),
    .X(_01237_));
 sky130_fd_sc_hd__nor2_1 _14269_ (.A(_09209_),
    .B(_10476_),
    .Y(_10483_));
 sky130_fd_sc_hd__a31o_1 _14270_ (.A1(_10436_),
    .A2(net537),
    .A3(_10472_),
    .B1(_10483_),
    .X(_01238_));
 sky130_fd_sc_hd__and3_1 _14271_ (.A(_10470_),
    .B(_09326_),
    .C(_10480_),
    .X(_10484_));
 sky130_fd_sc_hd__a31o_1 _14272_ (.A1(_10436_),
    .A2(net987),
    .A3(_10472_),
    .B1(_10484_),
    .X(_01239_));
 sky130_fd_sc_hd__buf_4 _14273_ (.A(_10279_),
    .X(_10485_));
 sky130_fd_sc_hd__nor2_1 _14274_ (.A(_09216_),
    .B(_10471_),
    .Y(_10486_));
 sky130_fd_sc_hd__a31o_1 _14275_ (.A1(_10485_),
    .A2(net1311),
    .A3(_10476_),
    .B1(_10486_),
    .X(_01224_));
 sky130_fd_sc_hd__nand2_1 _14276_ (.A(_10226_),
    .B(net3862),
    .Y(_10487_));
 sky130_fd_sc_hd__o2bb2a_1 _14277_ (.A1_N(_10487_),
    .A2_N(_10472_),
    .B1(_10257_),
    .B2(_10473_),
    .X(_01225_));
 sky130_fd_sc_hd__clkbuf_8 _14278_ (.A(_09375_),
    .X(_10488_));
 sky130_fd_sc_hd__nand2_1 _14279_ (.A(_10488_),
    .B(net3721),
    .Y(_10489_));
 sky130_fd_sc_hd__o2bb2a_1 _14280_ (.A1_N(_10489_),
    .A2_N(_10472_),
    .B1(_10259_),
    .B2(_10473_),
    .X(_01226_));
 sky130_fd_sc_hd__nor2_1 _14281_ (.A(_09230_),
    .B(_10471_),
    .Y(_10490_));
 sky130_fd_sc_hd__a31o_1 _14282_ (.A1(_10485_),
    .A2(net1579),
    .A3(_10476_),
    .B1(_10490_),
    .X(_01227_));
 sky130_fd_sc_hd__nor2_1 _14283_ (.A(_09233_),
    .B(_10471_),
    .Y(_10491_));
 sky130_fd_sc_hd__a31o_1 _14284_ (.A1(_10485_),
    .A2(net2106),
    .A3(_10476_),
    .B1(_10491_),
    .X(_01228_));
 sky130_fd_sc_hd__nand2_1 _14285_ (.A(_10488_),
    .B(net3853),
    .Y(_10492_));
 sky130_fd_sc_hd__inv_2 _14286_ (.A(_09337_),
    .Y(_10493_));
 sky130_fd_sc_hd__o2bb2a_1 _14287_ (.A1_N(_10492_),
    .A2_N(_10472_),
    .B1(_10493_),
    .B2(_10473_),
    .X(_01229_));
 sky130_fd_sc_hd__and3_1 _14288_ (.A(_10470_),
    .B(_09341_),
    .C(_10480_),
    .X(_10494_));
 sky130_fd_sc_hd__a31o_1 _14289_ (.A1(_10485_),
    .A2(net1451),
    .A3(_10476_),
    .B1(_10494_),
    .X(_01230_));
 sky130_fd_sc_hd__nor2_1 _14290_ (.A(_09243_),
    .B(_10471_),
    .Y(_10495_));
 sky130_fd_sc_hd__a31o_1 _14291_ (.A1(_10485_),
    .A2(net1013),
    .A3(_10476_),
    .B1(_10495_),
    .X(_01231_));
 sky130_fd_sc_hd__nor2_1 _14292_ (.A(_09246_),
    .B(_10471_),
    .Y(_10496_));
 sky130_fd_sc_hd__a31o_1 _14293_ (.A1(_10485_),
    .A2(net1503),
    .A3(_10476_),
    .B1(_10496_),
    .X(_01216_));
 sky130_fd_sc_hd__nand2_1 _14294_ (.A(_10488_),
    .B(net3878),
    .Y(_10497_));
 sky130_fd_sc_hd__inv_2 _14295_ (.A(_09248_),
    .Y(_10498_));
 sky130_fd_sc_hd__o2bb2a_1 _14296_ (.A1_N(_10497_),
    .A2_N(_10472_),
    .B1(_10498_),
    .B2(_10473_),
    .X(_01217_));
 sky130_fd_sc_hd__nor2_1 _14297_ (.A(_09253_),
    .B(_10471_),
    .Y(_10499_));
 sky130_fd_sc_hd__a31o_1 _14298_ (.A1(_10485_),
    .A2(net1717),
    .A3(_10476_),
    .B1(_10499_),
    .X(_01218_));
 sky130_fd_sc_hd__clkbuf_16 _14299_ (.A(net52),
    .X(_10500_));
 sky130_fd_sc_hd__and3_1 _14300_ (.A(_10470_),
    .B(_10500_),
    .C(_10480_),
    .X(_10501_));
 sky130_fd_sc_hd__a31o_1 _14301_ (.A1(_10485_),
    .A2(net1975),
    .A3(_10476_),
    .B1(_10501_),
    .X(_01219_));
 sky130_fd_sc_hd__nand2_1 _14302_ (.A(_10488_),
    .B(net3944),
    .Y(_10502_));
 sky130_fd_sc_hd__inv_2 _14303_ (.A(_09353_),
    .Y(_10503_));
 sky130_fd_sc_hd__o2bb2a_1 _14304_ (.A1_N(_10502_),
    .A2_N(_10472_),
    .B1(_10503_),
    .B2(_10473_),
    .X(_01220_));
 sky130_fd_sc_hd__nand2_1 _14305_ (.A(_10488_),
    .B(net3750),
    .Y(_10504_));
 sky130_fd_sc_hd__o2bb2a_1 _14306_ (.A1_N(_10504_),
    .A2_N(_10472_),
    .B1(_10273_),
    .B2(_10473_),
    .X(_01221_));
 sky130_fd_sc_hd__and3_1 _14307_ (.A(_10470_),
    .B(_09266_),
    .C(_10480_),
    .X(_10505_));
 sky130_fd_sc_hd__a31o_1 _14308_ (.A1(_10485_),
    .A2(net2224),
    .A3(_10476_),
    .B1(_10505_),
    .X(_01222_));
 sky130_fd_sc_hd__nand2_1 _14309_ (.A(_10488_),
    .B(net3873),
    .Y(_10506_));
 sky130_fd_sc_hd__o2bb2a_1 _14310_ (.A1_N(_10506_),
    .A2_N(_10472_),
    .B1(_10276_),
    .B2(_10473_),
    .X(_01223_));
 sky130_fd_sc_hd__and3_1 _14311_ (.A(_10470_),
    .B(_09274_),
    .C(_10480_),
    .X(_10507_));
 sky130_fd_sc_hd__a31o_1 _14312_ (.A1(_10485_),
    .A2(net2154),
    .A3(_10476_),
    .B1(_10507_),
    .X(_01208_));
 sky130_fd_sc_hd__nor2_1 _14313_ (.A(_09277_),
    .B(_10471_),
    .Y(_10508_));
 sky130_fd_sc_hd__a31o_1 _14314_ (.A1(_10485_),
    .A2(net1628),
    .A3(_10476_),
    .B1(_10508_),
    .X(_01209_));
 sky130_fd_sc_hd__and3_1 _14315_ (.A(_10470_),
    .B(_09369_),
    .C(_10480_),
    .X(_10509_));
 sky130_fd_sc_hd__a31o_1 _14316_ (.A1(_10485_),
    .A2(net1413),
    .A3(_10476_),
    .B1(_10509_),
    .X(_01210_));
 sky130_fd_sc_hd__nand2_1 _14317_ (.A(_10488_),
    .B(net4116),
    .Y(_10510_));
 sky130_fd_sc_hd__o2bb2a_1 _14318_ (.A1_N(_10510_),
    .A2_N(_10472_),
    .B1(_10285_),
    .B2(_10473_),
    .X(_01211_));
 sky130_fd_sc_hd__and3_1 _14319_ (.A(_10470_),
    .B(_09373_),
    .C(_10480_),
    .X(_10511_));
 sky130_fd_sc_hd__a31o_1 _14320_ (.A1(_10485_),
    .A2(net2373),
    .A3(_10476_),
    .B1(_10511_),
    .X(_01212_));
 sky130_fd_sc_hd__and3_1 _14321_ (.A(_10470_),
    .B(_09730_),
    .C(_10480_),
    .X(_10512_));
 sky130_fd_sc_hd__a31o_1 _14322_ (.A1(_10485_),
    .A2(net1819),
    .A3(_10476_),
    .B1(_10512_),
    .X(_01213_));
 sky130_fd_sc_hd__nand2_1 _14323_ (.A(_10350_),
    .B(net3699),
    .Y(_10513_));
 sky130_fd_sc_hd__a22o_1 _14324_ (.A1(_10348_),
    .A2(_10470_),
    .B1(_10471_),
    .B2(_10513_),
    .X(_10514_));
 sky130_fd_sc_hd__inv_2 _14325_ (.A(net3700),
    .Y(_01214_));
 sky130_fd_sc_hd__nand2_1 _14326_ (.A(_10350_),
    .B(net3077),
    .Y(_10515_));
 sky130_fd_sc_hd__a22o_1 _14327_ (.A1(net142),
    .A2(_10470_),
    .B1(_10471_),
    .B2(_10515_),
    .X(_10516_));
 sky130_fd_sc_hd__inv_2 _14328_ (.A(net3078),
    .Y(_01215_));
 sky130_fd_sc_hd__nor2_2 _14329_ (.A(_10467_),
    .B(_10292_),
    .Y(_10517_));
 sky130_fd_sc_hd__inv_2 _14330_ (.A(_10517_),
    .Y(_10518_));
 sky130_fd_sc_hd__nor2_1 _14331_ (.A(_08727_),
    .B(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__clkinv_4 _14332_ (.A(_10519_),
    .Y(_10520_));
 sky130_fd_sc_hd__buf_4 _14333_ (.A(_10520_),
    .X(_10521_));
 sky130_fd_sc_hd__buf_4 _14334_ (.A(_10520_),
    .X(_10522_));
 sky130_fd_sc_hd__nor2_1 _14335_ (.A(_09181_),
    .B(_10522_),
    .Y(_10523_));
 sky130_fd_sc_hd__a31o_1 _14336_ (.A1(_10485_),
    .A2(net909),
    .A3(_10521_),
    .B1(_10523_),
    .X(_01200_));
 sky130_fd_sc_hd__nor2_8 _14337_ (.A(_08794_),
    .B(_10518_),
    .Y(_10524_));
 sky130_fd_sc_hd__nand2_1 _14338_ (.A(_10350_),
    .B(net3903),
    .Y(_10525_));
 sky130_fd_sc_hd__a22o_1 _14339_ (.A1(_10524_),
    .A2(_09315_),
    .B1(_10522_),
    .B2(_10525_),
    .X(_10526_));
 sky130_fd_sc_hd__inv_2 _14340_ (.A(_10526_),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _14341_ (.A(_09188_),
    .B(_10522_),
    .Y(_10527_));
 sky130_fd_sc_hd__a31o_1 _14342_ (.A1(_10485_),
    .A2(net2188),
    .A3(_10521_),
    .B1(_10527_),
    .X(_01202_));
 sky130_fd_sc_hd__and3_1 _14343_ (.A(_10517_),
    .B(_09463_),
    .C(_10480_),
    .X(_10528_));
 sky130_fd_sc_hd__a31o_1 _14344_ (.A1(_10521_),
    .A2(_10277_),
    .A3(net2578),
    .B1(_10528_),
    .X(_01203_));
 sky130_fd_sc_hd__nand2_1 _14345_ (.A(_10350_),
    .B(net3434),
    .Y(_10529_));
 sky130_fd_sc_hd__a22o_1 _14346_ (.A1(_10524_),
    .A2(_09201_),
    .B1(_10522_),
    .B2(_10529_),
    .X(_10530_));
 sky130_fd_sc_hd__inv_2 _14347_ (.A(_10530_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _14348_ (.A(_10350_),
    .B(net3533),
    .Y(_10531_));
 sky130_fd_sc_hd__a22o_1 _14349_ (.A1(_10524_),
    .A2(_09205_),
    .B1(_10522_),
    .B2(_10531_),
    .X(_10532_));
 sky130_fd_sc_hd__inv_2 _14350_ (.A(_10532_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _14351_ (.A(_10350_),
    .B(net3850),
    .Y(_10533_));
 sky130_fd_sc_hd__a22o_1 _14352_ (.A1(_10524_),
    .A2(_09398_),
    .B1(_10522_),
    .B2(_10533_),
    .X(_10534_));
 sky130_fd_sc_hd__inv_2 _14353_ (.A(_10534_),
    .Y(_01206_));
 sky130_fd_sc_hd__and3_1 _14354_ (.A(_10517_),
    .B(_09326_),
    .C(_10480_),
    .X(_10535_));
 sky130_fd_sc_hd__a31o_1 _14355_ (.A1(_10521_),
    .A2(_10277_),
    .A3(net2456),
    .B1(_10535_),
    .X(_01207_));
 sky130_fd_sc_hd__nand2_1 _14356_ (.A(_10350_),
    .B(net3616),
    .Y(_10536_));
 sky130_fd_sc_hd__a22o_1 _14357_ (.A1(_10524_),
    .A2(_09531_),
    .B1(_10522_),
    .B2(_10536_),
    .X(_10537_));
 sky130_fd_sc_hd__inv_2 _14358_ (.A(_10537_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _14359_ (.A(_10350_),
    .B(net2791),
    .Y(_10538_));
 sky130_fd_sc_hd__a22o_1 _14360_ (.A1(_10524_),
    .A2(_10122_),
    .B1(_10522_),
    .B2(_10538_),
    .X(_10539_));
 sky130_fd_sc_hd__inv_2 _14361_ (.A(_10539_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_1 _14362_ (.A(_10350_),
    .B(net2904),
    .Y(_10540_));
 sky130_fd_sc_hd__a22o_1 _14363_ (.A1(_10524_),
    .A2(_10195_),
    .B1(_10520_),
    .B2(_10540_),
    .X(_10541_));
 sky130_fd_sc_hd__inv_2 _14364_ (.A(_10541_),
    .Y(_01194_));
 sky130_fd_sc_hd__buf_4 _14365_ (.A(_10279_),
    .X(_10542_));
 sky130_fd_sc_hd__nor2_1 _14366_ (.A(_09230_),
    .B(_10522_),
    .Y(_10543_));
 sky130_fd_sc_hd__a31o_1 _14367_ (.A1(_10542_),
    .A2(net1691),
    .A3(_10521_),
    .B1(_10543_),
    .X(_01195_));
 sky130_fd_sc_hd__nor2_1 _14368_ (.A(_09233_),
    .B(_10522_),
    .Y(_10544_));
 sky130_fd_sc_hd__a31o_1 _14369_ (.A1(_10542_),
    .A2(net1029),
    .A3(_10521_),
    .B1(_10544_),
    .X(_01196_));
 sky130_fd_sc_hd__nor2_1 _14370_ (.A(_09236_),
    .B(_10522_),
    .Y(_10545_));
 sky130_fd_sc_hd__a31o_1 _14371_ (.A1(_10542_),
    .A2(net955),
    .A3(_10521_),
    .B1(_10545_),
    .X(_01197_));
 sky130_fd_sc_hd__nand2_1 _14372_ (.A(_10350_),
    .B(net3374),
    .Y(_10546_));
 sky130_fd_sc_hd__a22o_1 _14373_ (.A1(_10524_),
    .A2(_10202_),
    .B1(_10520_),
    .B2(_10546_),
    .X(_10547_));
 sky130_fd_sc_hd__inv_2 _14374_ (.A(_10547_),
    .Y(_01198_));
 sky130_fd_sc_hd__nor2_1 _14375_ (.A(_09243_),
    .B(_10522_),
    .Y(_10548_));
 sky130_fd_sc_hd__a31o_1 _14376_ (.A1(_10542_),
    .A2(net2125),
    .A3(_10521_),
    .B1(_10548_),
    .X(_01199_));
 sky130_fd_sc_hd__nor2_1 _14377_ (.A(_09246_),
    .B(_10522_),
    .Y(_10549_));
 sky130_fd_sc_hd__a31o_1 _14378_ (.A1(_10542_),
    .A2(net635),
    .A3(_10521_),
    .B1(_10549_),
    .X(_01184_));
 sky130_fd_sc_hd__and3_1 _14379_ (.A(_10517_),
    .B(_09345_),
    .C(_10480_),
    .X(_10550_));
 sky130_fd_sc_hd__a31o_1 _14380_ (.A1(_10521_),
    .A2(_10277_),
    .A3(net2071),
    .B1(_10550_),
    .X(_01185_));
 sky130_fd_sc_hd__nor2_1 _14381_ (.A(_09253_),
    .B(_10522_),
    .Y(_10551_));
 sky130_fd_sc_hd__a31o_1 _14382_ (.A1(_10542_),
    .A2(net2388),
    .A3(_10521_),
    .B1(_10551_),
    .X(_01186_));
 sky130_fd_sc_hd__and3_1 _14383_ (.A(_10517_),
    .B(_10500_),
    .C(_10480_),
    .X(_10552_));
 sky130_fd_sc_hd__a31o_1 _14384_ (.A1(_10521_),
    .A2(_10277_),
    .A3(net2441),
    .B1(_10552_),
    .X(_01187_));
 sky130_fd_sc_hd__nor2_1 _14385_ (.A(_09260_),
    .B(_10522_),
    .Y(_10553_));
 sky130_fd_sc_hd__a31o_1 _14386_ (.A1(_10542_),
    .A2(net1803),
    .A3(_10521_),
    .B1(_10553_),
    .X(_01188_));
 sky130_fd_sc_hd__buf_4 _14387_ (.A(_10349_),
    .X(_10554_));
 sky130_fd_sc_hd__nand2_1 _14388_ (.A(_10554_),
    .B(net3645),
    .Y(_10555_));
 sky130_fd_sc_hd__a22o_1 _14389_ (.A1(_10524_),
    .A2(_10149_),
    .B1(_10520_),
    .B2(_10555_),
    .X(_10556_));
 sky130_fd_sc_hd__inv_2 _14390_ (.A(_10556_),
    .Y(_01189_));
 sky130_fd_sc_hd__and3_1 _14391_ (.A(_10517_),
    .B(_09266_),
    .C(_10480_),
    .X(_10557_));
 sky130_fd_sc_hd__a31o_1 _14392_ (.A1(_10521_),
    .A2(_10277_),
    .A3(net2272),
    .B1(_10557_),
    .X(_01190_));
 sky130_fd_sc_hd__nand2_1 _14393_ (.A(_10554_),
    .B(net3172),
    .Y(_10558_));
 sky130_fd_sc_hd__a22o_1 _14394_ (.A1(_10524_),
    .A2(_10154_),
    .B1(_10520_),
    .B2(_10558_),
    .X(_10559_));
 sky130_fd_sc_hd__inv_2 _14395_ (.A(_10559_),
    .Y(_01191_));
 sky130_fd_sc_hd__nand2_1 _14396_ (.A(_10554_),
    .B(net4051),
    .Y(_10560_));
 sky130_fd_sc_hd__a22o_1 _14397_ (.A1(_10524_),
    .A2(_09495_),
    .B1(_10520_),
    .B2(_10560_),
    .X(_10561_));
 sky130_fd_sc_hd__inv_2 _14398_ (.A(_10561_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_1 _14399_ (.A(_10554_),
    .B(net3858),
    .Y(_10562_));
 sky130_fd_sc_hd__a22o_1 _14400_ (.A1(_10524_),
    .A2(_09366_),
    .B1(_10520_),
    .B2(_10562_),
    .X(_10563_));
 sky130_fd_sc_hd__inv_2 _14401_ (.A(_10563_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_1 _14402_ (.A(_10554_),
    .B(net3825),
    .Y(_10564_));
 sky130_fd_sc_hd__a22o_1 _14403_ (.A1(_10524_),
    .A2(_09280_),
    .B1(_10520_),
    .B2(_10564_),
    .X(_10565_));
 sky130_fd_sc_hd__inv_2 _14404_ (.A(_10565_),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_1 _14405_ (.A(_10554_),
    .B(net3468),
    .Y(_10566_));
 sky130_fd_sc_hd__a22o_1 _14406_ (.A1(_10524_),
    .A2(_10164_),
    .B1(_10520_),
    .B2(_10566_),
    .X(_10567_));
 sky130_fd_sc_hd__inv_2 _14407_ (.A(_10567_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand2_1 _14408_ (.A(_10554_),
    .B(net3476),
    .Y(_10568_));
 sky130_fd_sc_hd__a22o_1 _14409_ (.A1(_10524_),
    .A2(_09288_),
    .B1(_10520_),
    .B2(_10568_),
    .X(_10569_));
 sky130_fd_sc_hd__inv_2 _14410_ (.A(_10569_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _14411_ (.A(_10554_),
    .B(net3762),
    .Y(_10570_));
 sky130_fd_sc_hd__a22o_1 _14412_ (.A1(_10524_),
    .A2(_09504_),
    .B1(_10520_),
    .B2(_10570_),
    .X(_10571_));
 sky130_fd_sc_hd__inv_2 _14413_ (.A(_10571_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand2_1 _14414_ (.A(_10488_),
    .B(net4023),
    .Y(_10572_));
 sky130_fd_sc_hd__o2bb2a_1 _14415_ (.A1_N(_10572_),
    .A2_N(_10521_),
    .B1(_10289_),
    .B2(_10518_),
    .X(_01182_));
 sky130_fd_sc_hd__nor2_1 _14416_ (.A(_09300_),
    .B(_10522_),
    .Y(_10573_));
 sky130_fd_sc_hd__a31o_1 _14417_ (.A1(_10542_),
    .A2(net2089),
    .A3(_10521_),
    .B1(_10573_),
    .X(_01183_));
 sky130_fd_sc_hd__nor2_2 _14418_ (.A(_10467_),
    .B(_10356_),
    .Y(_10574_));
 sky130_fd_sc_hd__inv_2 _14419_ (.A(_10574_),
    .Y(_10575_));
 sky130_fd_sc_hd__nor2_1 _14420_ (.A(_09166_),
    .B(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__inv_2 _14421_ (.A(_10576_),
    .Y(_10577_));
 sky130_fd_sc_hd__buf_4 _14422_ (.A(_10577_),
    .X(_10578_));
 sky130_fd_sc_hd__buf_4 _14423_ (.A(_10577_),
    .X(_10579_));
 sky130_fd_sc_hd__nor2_1 _14424_ (.A(_09181_),
    .B(_10579_),
    .Y(_10580_));
 sky130_fd_sc_hd__a31o_1 _14425_ (.A1(_10542_),
    .A2(net669),
    .A3(_10578_),
    .B1(_10580_),
    .X(_01168_));
 sky130_fd_sc_hd__nor2_1 _14426_ (.A(_09185_),
    .B(_10579_),
    .Y(_10581_));
 sky130_fd_sc_hd__a31o_1 _14427_ (.A1(_10542_),
    .A2(net2308),
    .A3(_10578_),
    .B1(_10581_),
    .X(_01169_));
 sky130_fd_sc_hd__nor2_1 _14428_ (.A(_09188_),
    .B(_10579_),
    .Y(_10582_));
 sky130_fd_sc_hd__a31o_1 _14429_ (.A1(_10542_),
    .A2(net667),
    .A3(_10578_),
    .B1(_10582_),
    .X(_01170_));
 sky130_fd_sc_hd__nor2_4 _14430_ (.A(_08795_),
    .B(_10575_),
    .Y(_10583_));
 sky130_fd_sc_hd__nand2_1 _14431_ (.A(_10554_),
    .B(net3646),
    .Y(_10584_));
 sky130_fd_sc_hd__a22o_1 _14432_ (.A1(_10583_),
    .A2(_09195_),
    .B1(_10577_),
    .B2(_10584_),
    .X(_10585_));
 sky130_fd_sc_hd__inv_2 _14433_ (.A(_10585_),
    .Y(_01171_));
 sky130_fd_sc_hd__buf_12 _14434_ (.A(net70),
    .X(_10586_));
 sky130_fd_sc_hd__buf_8 _14435_ (.A(_10586_),
    .X(_10587_));
 sky130_fd_sc_hd__and3_1 _14436_ (.A(_10574_),
    .B(_10587_),
    .C(_10480_),
    .X(_10588_));
 sky130_fd_sc_hd__a31o_1 _14437_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net1548),
    .B1(_10588_),
    .X(_01172_));
 sky130_fd_sc_hd__and3_1 _14438_ (.A(_10574_),
    .B(_09395_),
    .C(_10480_),
    .X(_10589_));
 sky130_fd_sc_hd__a31o_1 _14439_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net1595),
    .B1(_10589_),
    .X(_01173_));
 sky130_fd_sc_hd__nor2_1 _14440_ (.A(_09209_),
    .B(_10579_),
    .Y(_10590_));
 sky130_fd_sc_hd__a31o_1 _14441_ (.A1(_10542_),
    .A2(net1217),
    .A3(_10578_),
    .B1(_10590_),
    .X(_01174_));
 sky130_fd_sc_hd__buf_12 _14442_ (.A(_09211_),
    .X(_10591_));
 sky130_fd_sc_hd__nand2_1 _14443_ (.A(_10554_),
    .B(net4047),
    .Y(_10592_));
 sky130_fd_sc_hd__a22o_1 _14444_ (.A1(_10583_),
    .A2(_10591_),
    .B1(_10577_),
    .B2(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__inv_2 _14445_ (.A(_10593_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor2_1 _14446_ (.A(_09216_),
    .B(_10579_),
    .Y(_10594_));
 sky130_fd_sc_hd__a31o_1 _14447_ (.A1(_10542_),
    .A2(net493),
    .A3(_10578_),
    .B1(_10594_),
    .X(_01160_));
 sky130_fd_sc_hd__nand2_1 _14448_ (.A(_10554_),
    .B(net3882),
    .Y(_10595_));
 sky130_fd_sc_hd__a22o_1 _14449_ (.A1(_10583_),
    .A2(_10122_),
    .B1(_10577_),
    .B2(_10595_),
    .X(_10596_));
 sky130_fd_sc_hd__inv_2 _14450_ (.A(_10596_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2_1 _14451_ (.A(_10554_),
    .B(net3651),
    .Y(_10597_));
 sky130_fd_sc_hd__a22o_1 _14452_ (.A1(_10583_),
    .A2(_10195_),
    .B1(_10577_),
    .B2(_10597_),
    .X(_10598_));
 sky130_fd_sc_hd__inv_2 _14453_ (.A(_10598_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2_1 _14454_ (.A(_10554_),
    .B(net3883),
    .Y(_10599_));
 sky130_fd_sc_hd__a22o_1 _14455_ (.A1(_10583_),
    .A2(_09589_),
    .B1(_10577_),
    .B2(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__inv_2 _14456_ (.A(_10600_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_1 _14457_ (.A(_09233_),
    .B(_10579_),
    .Y(_10601_));
 sky130_fd_sc_hd__a31o_1 _14458_ (.A1(_10542_),
    .A2(net1083),
    .A3(_10578_),
    .B1(_10601_),
    .X(_01164_));
 sky130_fd_sc_hd__buf_12 _14459_ (.A(_09235_),
    .X(_10602_));
 sky130_fd_sc_hd__nor2_1 _14460_ (.A(_10602_),
    .B(_10579_),
    .Y(_10603_));
 sky130_fd_sc_hd__a31o_1 _14461_ (.A1(_10542_),
    .A2(net775),
    .A3(_10579_),
    .B1(_10603_),
    .X(_01165_));
 sky130_fd_sc_hd__nand2_1 _14462_ (.A(_10554_),
    .B(net3499),
    .Y(_10604_));
 sky130_fd_sc_hd__a22o_1 _14463_ (.A1(_10583_),
    .A2(_10202_),
    .B1(_10577_),
    .B2(_10604_),
    .X(_10605_));
 sky130_fd_sc_hd__inv_2 _14464_ (.A(_10605_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand2_1 _14465_ (.A(_10554_),
    .B(net3970),
    .Y(_10606_));
 sky130_fd_sc_hd__a22o_1 _14466_ (.A1(_10583_),
    .A2(_09768_),
    .B1(_10577_),
    .B2(_10606_),
    .X(_10607_));
 sky130_fd_sc_hd__inv_2 _14467_ (.A(_10607_),
    .Y(_01167_));
 sky130_fd_sc_hd__nor2_1 _14468_ (.A(_09246_),
    .B(_10579_),
    .Y(_10608_));
 sky130_fd_sc_hd__a31o_1 _14469_ (.A1(_10542_),
    .A2(net481),
    .A3(_10579_),
    .B1(_10608_),
    .X(_01144_));
 sky130_fd_sc_hd__clkbuf_4 _14470_ (.A(_09359_),
    .X(_10609_));
 sky130_fd_sc_hd__and3_1 _14471_ (.A(_10574_),
    .B(_09345_),
    .C(_10609_),
    .X(_10610_));
 sky130_fd_sc_hd__a31o_1 _14472_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net707),
    .B1(_10610_),
    .X(_01145_));
 sky130_fd_sc_hd__buf_4 _14473_ (.A(_10279_),
    .X(_10611_));
 sky130_fd_sc_hd__nor2_1 _14474_ (.A(_09253_),
    .B(_10579_),
    .Y(_10612_));
 sky130_fd_sc_hd__a31o_1 _14475_ (.A1(_10611_),
    .A2(net425),
    .A3(_10579_),
    .B1(_10612_),
    .X(_01146_));
 sky130_fd_sc_hd__and3_1 _14476_ (.A(_10574_),
    .B(_10500_),
    .C(_10609_),
    .X(_10613_));
 sky130_fd_sc_hd__a31o_1 _14477_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net619),
    .B1(_10613_),
    .X(_01147_));
 sky130_fd_sc_hd__nor2_1 _14478_ (.A(_09260_),
    .B(_10579_),
    .Y(_10614_));
 sky130_fd_sc_hd__a31o_1 _14479_ (.A1(_10611_),
    .A2(net519),
    .A3(_10579_),
    .B1(_10614_),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_1 _14480_ (.A(_10554_),
    .B(net3879),
    .Y(_10615_));
 sky130_fd_sc_hd__a22o_1 _14481_ (.A1(_10583_),
    .A2(_10149_),
    .B1(_10577_),
    .B2(_10615_),
    .X(_10616_));
 sky130_fd_sc_hd__inv_2 _14482_ (.A(_10616_),
    .Y(_01149_));
 sky130_fd_sc_hd__buf_8 _14483_ (.A(net55),
    .X(_10617_));
 sky130_fd_sc_hd__and3_1 _14484_ (.A(_10574_),
    .B(_10617_),
    .C(_10609_),
    .X(_10618_));
 sky130_fd_sc_hd__a31o_1 _14485_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net645),
    .B1(_10618_),
    .X(_01150_));
 sky130_fd_sc_hd__buf_4 _14486_ (.A(_10349_),
    .X(_10619_));
 sky130_fd_sc_hd__nand2_1 _14487_ (.A(_10619_),
    .B(net2874),
    .Y(_10620_));
 sky130_fd_sc_hd__a22o_1 _14488_ (.A1(_10583_),
    .A2(_10154_),
    .B1(_10577_),
    .B2(_10620_),
    .X(_10621_));
 sky130_fd_sc_hd__inv_2 _14489_ (.A(_10621_),
    .Y(_01151_));
 sky130_fd_sc_hd__and3_1 _14490_ (.A(_10574_),
    .B(_09274_),
    .C(_10609_),
    .X(_10622_));
 sky130_fd_sc_hd__a31o_1 _14491_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net1245),
    .B1(_10622_),
    .X(_01136_));
 sky130_fd_sc_hd__nor2_1 _14492_ (.A(_09277_),
    .B(_10579_),
    .Y(_10623_));
 sky130_fd_sc_hd__a31o_1 _14493_ (.A1(_10611_),
    .A2(net439),
    .A3(_10579_),
    .B1(_10623_),
    .X(_01137_));
 sky130_fd_sc_hd__buf_12 _14494_ (.A(_09279_),
    .X(_10624_));
 sky130_fd_sc_hd__nand2_1 _14495_ (.A(_10619_),
    .B(net3008),
    .Y(_10625_));
 sky130_fd_sc_hd__a22o_1 _14496_ (.A1(_10583_),
    .A2(_10624_),
    .B1(_10577_),
    .B2(_10625_),
    .X(_10626_));
 sky130_fd_sc_hd__inv_2 _14497_ (.A(_10626_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand2_1 _14498_ (.A(_10619_),
    .B(net3713),
    .Y(_10627_));
 sky130_fd_sc_hd__a22o_1 _14499_ (.A1(_10583_),
    .A2(_10164_),
    .B1(_10577_),
    .B2(_10627_),
    .X(_10628_));
 sky130_fd_sc_hd__inv_2 _14500_ (.A(_10628_),
    .Y(_01139_));
 sky130_fd_sc_hd__and3_1 _14501_ (.A(_10574_),
    .B(_09373_),
    .C(_10609_),
    .X(_10629_));
 sky130_fd_sc_hd__a31o_1 _14502_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net587),
    .B1(_10629_),
    .X(_01140_));
 sky130_fd_sc_hd__and3_1 _14503_ (.A(_10574_),
    .B(_09730_),
    .C(_10609_),
    .X(_10630_));
 sky130_fd_sc_hd__a31o_1 _14504_ (.A1(_10578_),
    .A2(_10277_),
    .A3(net595),
    .B1(_10630_),
    .X(_01141_));
 sky130_fd_sc_hd__nand2_1 _14505_ (.A(_10488_),
    .B(net3663),
    .Y(_10631_));
 sky130_fd_sc_hd__o2bb2a_1 _14506_ (.A1_N(_10631_),
    .A2_N(_10578_),
    .B1(_10289_),
    .B2(_10575_),
    .X(_01142_));
 sky130_fd_sc_hd__nand2_1 _14507_ (.A(_10488_),
    .B(net3392),
    .Y(_10632_));
 sky130_fd_sc_hd__o2bb2a_1 _14508_ (.A1_N(_10632_),
    .A2_N(_10578_),
    .B1(_09442_),
    .B2(_10575_),
    .X(_01143_));
 sky130_fd_sc_hd__nor2_4 _14509_ (.A(_10467_),
    .B(_10411_),
    .Y(_10633_));
 sky130_fd_sc_hd__inv_2 _14510_ (.A(_10633_),
    .Y(_10634_));
 sky130_fd_sc_hd__nor2_1 _14511_ (.A(_09304_),
    .B(_10634_),
    .Y(_10635_));
 sky130_fd_sc_hd__inv_2 _14512_ (.A(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__buf_4 _14513_ (.A(_10636_),
    .X(_10637_));
 sky130_fd_sc_hd__buf_4 _14514_ (.A(_10636_),
    .X(_10638_));
 sky130_fd_sc_hd__nor2_1 _14515_ (.A(_09181_),
    .B(_10638_),
    .Y(_10639_));
 sky130_fd_sc_hd__a31o_1 _14516_ (.A1(_10611_),
    .A2(net565),
    .A3(_10637_),
    .B1(_10639_),
    .X(_01128_));
 sky130_fd_sc_hd__nor2_4 _14517_ (.A(_08795_),
    .B(_10634_),
    .Y(_10640_));
 sky130_fd_sc_hd__nand2_1 _14518_ (.A(_10619_),
    .B(net2803),
    .Y(_10641_));
 sky130_fd_sc_hd__a22o_1 _14519_ (.A1(_10640_),
    .A2(_09315_),
    .B1(_10638_),
    .B2(_10641_),
    .X(_10642_));
 sky130_fd_sc_hd__inv_2 _14520_ (.A(_10642_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_1 _14521_ (.A(_10619_),
    .B(net3226),
    .Y(_10643_));
 sky130_fd_sc_hd__a22o_1 _14522_ (.A1(_10640_),
    .A2(_09460_),
    .B1(_10636_),
    .B2(_10643_),
    .X(_10644_));
 sky130_fd_sc_hd__inv_2 _14523_ (.A(_10644_),
    .Y(_01130_));
 sky130_fd_sc_hd__buf_6 _14524_ (.A(_09222_),
    .X(_10645_));
 sky130_fd_sc_hd__clkbuf_8 _14525_ (.A(_10645_),
    .X(_10646_));
 sky130_fd_sc_hd__and3_1 _14526_ (.A(_10633_),
    .B(_09463_),
    .C(_10609_),
    .X(_10647_));
 sky130_fd_sc_hd__a31o_1 _14527_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net603),
    .B1(_10647_),
    .X(_01131_));
 sky130_fd_sc_hd__and3_1 _14528_ (.A(_10633_),
    .B(_10587_),
    .C(_10609_),
    .X(_10648_));
 sky130_fd_sc_hd__a31o_1 _14529_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net737),
    .B1(_10648_),
    .X(_01132_));
 sky130_fd_sc_hd__and3_1 _14530_ (.A(_10633_),
    .B(_09395_),
    .C(_10609_),
    .X(_10649_));
 sky130_fd_sc_hd__a31o_1 _14531_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net673),
    .B1(_10649_),
    .X(_01133_));
 sky130_fd_sc_hd__nor2_1 _14532_ (.A(_09209_),
    .B(_10638_),
    .Y(_10650_));
 sky130_fd_sc_hd__a31o_1 _14533_ (.A1(_10611_),
    .A2(net1558),
    .A3(_10637_),
    .B1(_10650_),
    .X(_01134_));
 sky130_fd_sc_hd__and3_1 _14534_ (.A(_10633_),
    .B(_09326_),
    .C(_10609_),
    .X(_10651_));
 sky130_fd_sc_hd__a31o_1 _14535_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net685),
    .B1(_10651_),
    .X(_01135_));
 sky130_fd_sc_hd__nor2_1 _14536_ (.A(_09216_),
    .B(_10638_),
    .Y(_10652_));
 sky130_fd_sc_hd__a31o_1 _14537_ (.A1(_10611_),
    .A2(net511),
    .A3(_10637_),
    .B1(_10652_),
    .X(_01120_));
 sky130_fd_sc_hd__nand2_1 _14538_ (.A(_10619_),
    .B(net2819),
    .Y(_10653_));
 sky130_fd_sc_hd__a22o_1 _14539_ (.A1(_10640_),
    .A2(_10122_),
    .B1(_10636_),
    .B2(_10653_),
    .X(_10654_));
 sky130_fd_sc_hd__inv_2 _14540_ (.A(_10654_),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_1 _14541_ (.A(_10619_),
    .B(net2912),
    .Y(_10655_));
 sky130_fd_sc_hd__a22o_1 _14542_ (.A1(_10640_),
    .A2(_10195_),
    .B1(_10636_),
    .B2(_10655_),
    .X(_10656_));
 sky130_fd_sc_hd__inv_2 _14543_ (.A(_10656_),
    .Y(_01122_));
 sky130_fd_sc_hd__buf_12 _14544_ (.A(_09229_),
    .X(_10657_));
 sky130_fd_sc_hd__nor2_1 _14545_ (.A(_10657_),
    .B(_10638_),
    .Y(_10658_));
 sky130_fd_sc_hd__a31o_1 _14546_ (.A1(_10611_),
    .A2(net429),
    .A3(_10638_),
    .B1(_10658_),
    .X(_01123_));
 sky130_fd_sc_hd__nor2_1 _14547_ (.A(_09233_),
    .B(_10638_),
    .Y(_10659_));
 sky130_fd_sc_hd__a31o_1 _14548_ (.A1(_10611_),
    .A2(net699),
    .A3(_10638_),
    .B1(_10659_),
    .X(_01124_));
 sky130_fd_sc_hd__nor2_1 _14549_ (.A(_10602_),
    .B(_10638_),
    .Y(_10660_));
 sky130_fd_sc_hd__a31o_1 _14550_ (.A1(_10611_),
    .A2(net487),
    .A3(_10638_),
    .B1(_10660_),
    .X(_01125_));
 sky130_fd_sc_hd__nand2_1 _14551_ (.A(_10619_),
    .B(net2813),
    .Y(_10661_));
 sky130_fd_sc_hd__a22o_1 _14552_ (.A1(_10640_),
    .A2(_10202_),
    .B1(_10636_),
    .B2(_10661_),
    .X(_10662_));
 sky130_fd_sc_hd__inv_2 _14553_ (.A(_10662_),
    .Y(_01126_));
 sky130_fd_sc_hd__buf_12 _14554_ (.A(_09242_),
    .X(_10663_));
 sky130_fd_sc_hd__nor2_1 _14555_ (.A(_10663_),
    .B(_10638_),
    .Y(_10664_));
 sky130_fd_sc_hd__a31o_1 _14556_ (.A1(_10611_),
    .A2(net423),
    .A3(_10638_),
    .B1(_10664_),
    .X(_01127_));
 sky130_fd_sc_hd__nand2_1 _14557_ (.A(_10619_),
    .B(net2780),
    .Y(_10665_));
 sky130_fd_sc_hd__a22o_1 _14558_ (.A1(_10640_),
    .A2(_09415_),
    .B1(_10636_),
    .B2(_10665_),
    .X(_10666_));
 sky130_fd_sc_hd__inv_2 _14559_ (.A(_10666_),
    .Y(_01112_));
 sky130_fd_sc_hd__buf_8 _14560_ (.A(net82),
    .X(_10667_));
 sky130_fd_sc_hd__and3_1 _14561_ (.A(_10633_),
    .B(_10667_),
    .C(_10609_),
    .X(_10668_));
 sky130_fd_sc_hd__a31o_1 _14562_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net2393),
    .B1(_10668_),
    .X(_01113_));
 sky130_fd_sc_hd__buf_12 _14563_ (.A(_09252_),
    .X(_10669_));
 sky130_fd_sc_hd__nor2_1 _14564_ (.A(_10669_),
    .B(_10638_),
    .Y(_10670_));
 sky130_fd_sc_hd__a31o_1 _14565_ (.A1(_10611_),
    .A2(net545),
    .A3(_10638_),
    .B1(_10670_),
    .X(_01114_));
 sky130_fd_sc_hd__and3_1 _14566_ (.A(_10633_),
    .B(_10500_),
    .C(_10609_),
    .X(_10671_));
 sky130_fd_sc_hd__a31o_1 _14567_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net1603),
    .B1(_10671_),
    .X(_01115_));
 sky130_fd_sc_hd__nand2_1 _14568_ (.A(_10619_),
    .B(net2825),
    .Y(_10672_));
 sky130_fd_sc_hd__a22o_1 _14569_ (.A1(_10640_),
    .A2(_09354_),
    .B1(_10636_),
    .B2(_10672_),
    .X(_10673_));
 sky130_fd_sc_hd__inv_2 _14570_ (.A(_10673_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _14571_ (.A(_10619_),
    .B(net2952),
    .Y(_10674_));
 sky130_fd_sc_hd__a22o_1 _14572_ (.A1(_10640_),
    .A2(_10149_),
    .B1(_10636_),
    .B2(_10674_),
    .X(_10675_));
 sky130_fd_sc_hd__inv_2 _14573_ (.A(_10675_),
    .Y(_01117_));
 sky130_fd_sc_hd__and3_1 _14574_ (.A(_10633_),
    .B(_10617_),
    .C(_10609_),
    .X(_10676_));
 sky130_fd_sc_hd__a31o_1 _14575_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net567),
    .B1(_10676_),
    .X(_01118_));
 sky130_fd_sc_hd__nand2_1 _14576_ (.A(_10619_),
    .B(net2776),
    .Y(_10677_));
 sky130_fd_sc_hd__a22o_1 _14577_ (.A1(_10640_),
    .A2(_10154_),
    .B1(_10636_),
    .B2(_10677_),
    .X(_10678_));
 sky130_fd_sc_hd__inv_2 _14578_ (.A(_10678_),
    .Y(_01119_));
 sky130_fd_sc_hd__clkbuf_16 _14579_ (.A(net50),
    .X(_10679_));
 sky130_fd_sc_hd__and3_1 _14580_ (.A(_10633_),
    .B(_10679_),
    .C(_10609_),
    .X(_10680_));
 sky130_fd_sc_hd__a31o_1 _14581_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net593),
    .B1(_10680_),
    .X(_01104_));
 sky130_fd_sc_hd__buf_12 _14582_ (.A(_09276_),
    .X(_10681_));
 sky130_fd_sc_hd__nor2_1 _14583_ (.A(_10681_),
    .B(_10638_),
    .Y(_10682_));
 sky130_fd_sc_hd__a31o_1 _14584_ (.A1(_10611_),
    .A2(net521),
    .A3(_10638_),
    .B1(_10682_),
    .X(_01105_));
 sky130_fd_sc_hd__and3_1 _14585_ (.A(_10633_),
    .B(_09369_),
    .C(_10609_),
    .X(_10683_));
 sky130_fd_sc_hd__a31o_1 _14586_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net961),
    .B1(_10683_),
    .X(_01106_));
 sky130_fd_sc_hd__nand2_1 _14587_ (.A(_10619_),
    .B(net2922),
    .Y(_10684_));
 sky130_fd_sc_hd__a22o_1 _14588_ (.A1(_10640_),
    .A2(_10164_),
    .B1(_10636_),
    .B2(_10684_),
    .X(_10685_));
 sky130_fd_sc_hd__inv_2 _14589_ (.A(_10685_),
    .Y(_01107_));
 sky130_fd_sc_hd__and3_1 _14590_ (.A(_10633_),
    .B(_09373_),
    .C(_10609_),
    .X(_10686_));
 sky130_fd_sc_hd__a31o_1 _14591_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net551),
    .B1(_10686_),
    .X(_01108_));
 sky130_fd_sc_hd__buf_4 _14592_ (.A(_09359_),
    .X(_10687_));
 sky130_fd_sc_hd__and3_1 _14593_ (.A(_10633_),
    .B(_09730_),
    .C(_10687_),
    .X(_10688_));
 sky130_fd_sc_hd__a31o_1 _14594_ (.A1(_10637_),
    .A2(_10646_),
    .A3(net637),
    .B1(_10688_),
    .X(_01109_));
 sky130_fd_sc_hd__nand2_1 _14595_ (.A(_10488_),
    .B(net3246),
    .Y(_10689_));
 sky130_fd_sc_hd__o2bb2a_1 _14596_ (.A1_N(_10689_),
    .A2_N(_10637_),
    .B1(_10289_),
    .B2(_10634_),
    .X(_01110_));
 sky130_fd_sc_hd__nand2_1 _14597_ (.A(_10488_),
    .B(net3301),
    .Y(_10690_));
 sky130_fd_sc_hd__o2bb2a_1 _14598_ (.A1_N(_10690_),
    .A2_N(_10637_),
    .B1(_09442_),
    .B2(_10634_),
    .X(_01111_));
 sky130_fd_sc_hd__nand2_8 _14599_ (.A(_09735_),
    .B(_10466_),
    .Y(_10691_));
 sky130_fd_sc_hd__nor2_8 _14600_ (.A(_10691_),
    .B(_10469_),
    .Y(_10692_));
 sky130_fd_sc_hd__nand2_2 _14601_ (.A(_10692_),
    .B(_10413_),
    .Y(_10693_));
 sky130_fd_sc_hd__buf_4 _14602_ (.A(_10693_),
    .X(_10694_));
 sky130_fd_sc_hd__buf_4 _14603_ (.A(_10693_),
    .X(_10695_));
 sky130_fd_sc_hd__nor2_1 _14604_ (.A(_09181_),
    .B(_10695_),
    .Y(_10696_));
 sky130_fd_sc_hd__a31o_1 _14605_ (.A1(_10611_),
    .A2(net2140),
    .A3(_10694_),
    .B1(_10696_),
    .X(_01096_));
 sky130_fd_sc_hd__nor2_1 _14606_ (.A(_09185_),
    .B(_10695_),
    .Y(_10697_));
 sky130_fd_sc_hd__a31o_1 _14607_ (.A1(_10611_),
    .A2(net1573),
    .A3(_10694_),
    .B1(_10697_),
    .X(_01097_));
 sky130_fd_sc_hd__buf_12 _14608_ (.A(_09187_),
    .X(_10698_));
 sky130_fd_sc_hd__nor2_1 _14609_ (.A(_10698_),
    .B(_10695_),
    .Y(_10699_));
 sky130_fd_sc_hd__a31o_1 _14610_ (.A1(_10611_),
    .A2(net2458),
    .A3(_10694_),
    .B1(_10699_),
    .X(_01098_));
 sky130_fd_sc_hd__nand2_1 _14611_ (.A(_10488_),
    .B(net4004),
    .Y(_10700_));
 sky130_fd_sc_hd__nand2_4 _14612_ (.A(_10692_),
    .B(_08778_),
    .Y(_10701_));
 sky130_fd_sc_hd__o2bb2a_1 _14613_ (.A1_N(_10700_),
    .A2_N(_10694_),
    .B1(_10479_),
    .B2(_10701_),
    .X(_01099_));
 sky130_fd_sc_hd__and3_1 _14614_ (.A(_10692_),
    .B(_10587_),
    .C(_10687_),
    .X(_10702_));
 sky130_fd_sc_hd__a31o_1 _14615_ (.A1(_10611_),
    .A2(net2621),
    .A3(_10694_),
    .B1(_10702_),
    .X(_01100_));
 sky130_fd_sc_hd__buf_4 _14616_ (.A(_10279_),
    .X(_10703_));
 sky130_fd_sc_hd__and3_1 _14617_ (.A(_10692_),
    .B(_09395_),
    .C(_10687_),
    .X(_10704_));
 sky130_fd_sc_hd__a31o_1 _14618_ (.A1(_10703_),
    .A2(net2121),
    .A3(_10694_),
    .B1(_10704_),
    .X(_01101_));
 sky130_fd_sc_hd__nor2_1 _14619_ (.A(_09209_),
    .B(_10695_),
    .Y(_10705_));
 sky130_fd_sc_hd__a31o_1 _14620_ (.A1(_10703_),
    .A2(net1365),
    .A3(_10694_),
    .B1(_10705_),
    .X(_01102_));
 sky130_fd_sc_hd__and3_1 _14621_ (.A(_10692_),
    .B(_09326_),
    .C(_10687_),
    .X(_10706_));
 sky130_fd_sc_hd__a31o_1 _14622_ (.A1(_10703_),
    .A2(net2477),
    .A3(_10694_),
    .B1(_10706_),
    .X(_01103_));
 sky130_fd_sc_hd__clkbuf_8 _14623_ (.A(_10310_),
    .X(_10707_));
 sky130_fd_sc_hd__a22o_1 _14624_ (.A1(_10707_),
    .A2(net2758),
    .B1(_10692_),
    .B2(_09227_),
    .X(_10708_));
 sky130_fd_sc_hd__o31a_1 _14625_ (.A1(_09193_),
    .A2(net57),
    .A3(_10701_),
    .B1(net2759),
    .X(_01088_));
 sky130_fd_sc_hd__nand2_1 _14626_ (.A(_10488_),
    .B(net3827),
    .Y(_10709_));
 sky130_fd_sc_hd__o2bb2a_1 _14627_ (.A1_N(_10709_),
    .A2_N(_10694_),
    .B1(_10257_),
    .B2(_10701_),
    .X(_01089_));
 sky130_fd_sc_hd__nand2_1 _14628_ (.A(_10488_),
    .B(net4195),
    .Y(_10710_));
 sky130_fd_sc_hd__o2bb2a_1 _14629_ (.A1_N(_10710_),
    .A2_N(_10694_),
    .B1(_10259_),
    .B2(_10701_),
    .X(_01090_));
 sky130_fd_sc_hd__nor2_1 _14630_ (.A(_10657_),
    .B(_10695_),
    .Y(_10711_));
 sky130_fd_sc_hd__a31o_1 _14631_ (.A1(_10703_),
    .A2(net2050),
    .A3(_10694_),
    .B1(_10711_),
    .X(_01091_));
 sky130_fd_sc_hd__a22o_1 _14632_ (.A1(_10707_),
    .A2(net3889),
    .B1(_10692_),
    .B2(_09227_),
    .X(_10712_));
 sky130_fd_sc_hd__o31a_1 _14633_ (.A1(_09193_),
    .A2(net62),
    .A3(_10701_),
    .B1(_10712_),
    .X(_01092_));
 sky130_fd_sc_hd__nor2_1 _14634_ (.A(_10602_),
    .B(_10695_),
    .Y(_10713_));
 sky130_fd_sc_hd__a31o_1 _14635_ (.A1(_10703_),
    .A2(net1727),
    .A3(_10695_),
    .B1(_10713_),
    .X(_01093_));
 sky130_fd_sc_hd__a22o_1 _14636_ (.A1(_10707_),
    .A2(net2834),
    .B1(_10692_),
    .B2(_09227_),
    .X(_10714_));
 sky130_fd_sc_hd__o31a_1 _14637_ (.A1(_09193_),
    .A2(_09341_),
    .A3(_10701_),
    .B1(_10714_),
    .X(_01094_));
 sky130_fd_sc_hd__nor2_1 _14638_ (.A(_10663_),
    .B(_10693_),
    .Y(_10715_));
 sky130_fd_sc_hd__a31o_1 _14639_ (.A1(_10703_),
    .A2(net2042),
    .A3(_10695_),
    .B1(_10715_),
    .X(_01095_));
 sky130_fd_sc_hd__a22o_1 _14640_ (.A1(_10707_),
    .A2(net2821),
    .B1(_10692_),
    .B2(_09227_),
    .X(_10716_));
 sky130_fd_sc_hd__o31a_1 _14641_ (.A1(_09193_),
    .A2(net81),
    .A3(_10701_),
    .B1(_10716_),
    .X(_01080_));
 sky130_fd_sc_hd__nand2_1 _14642_ (.A(_10488_),
    .B(net3764),
    .Y(_10717_));
 sky130_fd_sc_hd__o2bb2a_1 _14643_ (.A1_N(_10717_),
    .A2_N(_10694_),
    .B1(_10498_),
    .B2(_10701_),
    .X(_01081_));
 sky130_fd_sc_hd__nor2_1 _14644_ (.A(_10669_),
    .B(_10693_),
    .Y(_10718_));
 sky130_fd_sc_hd__a31o_1 _14645_ (.A1(_10703_),
    .A2(net1824),
    .A3(_10695_),
    .B1(_10718_),
    .X(_01082_));
 sky130_fd_sc_hd__and3_1 _14646_ (.A(_10692_),
    .B(_10500_),
    .C(_10687_),
    .X(_10719_));
 sky130_fd_sc_hd__a31o_1 _14647_ (.A1(_10703_),
    .A2(net2226),
    .A3(_10695_),
    .B1(_10719_),
    .X(_01083_));
 sky130_fd_sc_hd__nor2_1 _14648_ (.A(_09260_),
    .B(_10693_),
    .Y(_10720_));
 sky130_fd_sc_hd__a31o_1 _14649_ (.A1(_10703_),
    .A2(net1381),
    .A3(_10695_),
    .B1(_10720_),
    .X(_01084_));
 sky130_fd_sc_hd__buf_6 _14650_ (.A(_09375_),
    .X(_10721_));
 sky130_fd_sc_hd__nand2_1 _14651_ (.A(_10721_),
    .B(net4245),
    .Y(_10722_));
 sky130_fd_sc_hd__o2bb2a_1 _14652_ (.A1_N(_10722_),
    .A2_N(_10694_),
    .B1(_10273_),
    .B2(_10701_),
    .X(_01085_));
 sky130_fd_sc_hd__and3_1 _14653_ (.A(_10692_),
    .B(_10617_),
    .C(_10687_),
    .X(_10723_));
 sky130_fd_sc_hd__a31o_1 _14654_ (.A1(_10703_),
    .A2(net1678),
    .A3(_10695_),
    .B1(_10723_),
    .X(_01086_));
 sky130_fd_sc_hd__nand2_1 _14655_ (.A(_10721_),
    .B(net3872),
    .Y(_10724_));
 sky130_fd_sc_hd__o2bb2a_1 _14656_ (.A1_N(_10724_),
    .A2_N(_10694_),
    .B1(_10276_),
    .B2(_10701_),
    .X(_01087_));
 sky130_fd_sc_hd__and3_1 _14657_ (.A(_10692_),
    .B(_10679_),
    .C(_10687_),
    .X(_10725_));
 sky130_fd_sc_hd__a31o_1 _14658_ (.A1(_10703_),
    .A2(net1025),
    .A3(_10695_),
    .B1(_10725_),
    .X(_01072_));
 sky130_fd_sc_hd__nand2_1 _14659_ (.A(_10721_),
    .B(net3876),
    .Y(_10726_));
 sky130_fd_sc_hd__inv_2 _14660_ (.A(_09365_),
    .Y(_10727_));
 sky130_fd_sc_hd__o2bb2a_1 _14661_ (.A1_N(_10726_),
    .A2_N(_10694_),
    .B1(_10727_),
    .B2(_10701_),
    .X(_01073_));
 sky130_fd_sc_hd__buf_8 _14662_ (.A(net72),
    .X(_10728_));
 sky130_fd_sc_hd__and3_1 _14663_ (.A(_10692_),
    .B(_10728_),
    .C(_10687_),
    .X(_10729_));
 sky130_fd_sc_hd__a31o_1 _14664_ (.A1(_10703_),
    .A2(net925),
    .A3(_10695_),
    .B1(_10729_),
    .X(_01074_));
 sky130_fd_sc_hd__nand2_1 _14665_ (.A(_10721_),
    .B(net3988),
    .Y(_10730_));
 sky130_fd_sc_hd__o2bb2a_1 _14666_ (.A1_N(_10730_),
    .A2_N(_10694_),
    .B1(_10285_),
    .B2(_10701_),
    .X(_01075_));
 sky130_fd_sc_hd__a22o_1 _14667_ (.A1(_09302_),
    .A2(net3296),
    .B1(_10692_),
    .B2(_09227_),
    .X(_10731_));
 sky130_fd_sc_hd__o31a_1 _14668_ (.A1(_09193_),
    .A2(_09373_),
    .A3(_10701_),
    .B1(_10731_),
    .X(_01076_));
 sky130_fd_sc_hd__and3_1 _14669_ (.A(_10692_),
    .B(_09730_),
    .C(_10687_),
    .X(_10732_));
 sky130_fd_sc_hd__a31o_1 _14670_ (.A1(_10703_),
    .A2(net1804),
    .A3(_10695_),
    .B1(_10732_),
    .X(_01077_));
 sky130_fd_sc_hd__nand2_1 _14671_ (.A(_10619_),
    .B(net3068),
    .Y(_10733_));
 sky130_fd_sc_hd__a22o_1 _14672_ (.A1(_10348_),
    .A2(_10692_),
    .B1(_10693_),
    .B2(_10733_),
    .X(_10734_));
 sky130_fd_sc_hd__inv_2 _14673_ (.A(_10734_),
    .Y(_01078_));
 sky130_fd_sc_hd__nor2_1 _14674_ (.A(_09300_),
    .B(_10693_),
    .Y(_10735_));
 sky130_fd_sc_hd__a31o_1 _14675_ (.A1(_10703_),
    .A2(net2046),
    .A3(_10695_),
    .B1(_10735_),
    .X(_01079_));
 sky130_fd_sc_hd__nor2_2 _14676_ (.A(_10691_),
    .B(_10292_),
    .Y(_10736_));
 sky130_fd_sc_hd__inv_2 _14677_ (.A(_10736_),
    .Y(_10737_));
 sky130_fd_sc_hd__nor2_1 _14678_ (.A(_08797_),
    .B(_10737_),
    .Y(_10738_));
 sky130_fd_sc_hd__buf_4 _14679_ (.A(_10738_),
    .X(_10739_));
 sky130_fd_sc_hd__nor2_1 _14680_ (.A(_09625_),
    .B(_10737_),
    .Y(_10740_));
 sky130_fd_sc_hd__inv_2 _14681_ (.A(_10740_),
    .Y(_10741_));
 sky130_fd_sc_hd__buf_4 _14682_ (.A(_10741_),
    .X(_10742_));
 sky130_fd_sc_hd__nand2_1 _14683_ (.A(_10619_),
    .B(net3870),
    .Y(_10743_));
 sky130_fd_sc_hd__a22o_1 _14684_ (.A1(_10739_),
    .A2(_09451_),
    .B1(_10742_),
    .B2(_10743_),
    .X(_10744_));
 sky130_fd_sc_hd__inv_2 _14685_ (.A(_10744_),
    .Y(_01056_));
 sky130_fd_sc_hd__buf_4 _14686_ (.A(_10741_),
    .X(_10745_));
 sky130_fd_sc_hd__buf_12 _14687_ (.A(_09184_),
    .X(_10746_));
 sky130_fd_sc_hd__nor2_1 _14688_ (.A(_10746_),
    .B(_10745_),
    .Y(_10747_));
 sky130_fd_sc_hd__a31o_1 _14689_ (.A1(_10703_),
    .A2(net761),
    .A3(_10745_),
    .B1(_10747_),
    .X(_01057_));
 sky130_fd_sc_hd__nand2_1 _14690_ (.A(_10619_),
    .B(net3702),
    .Y(_10748_));
 sky130_fd_sc_hd__a22o_1 _14691_ (.A1(_10739_),
    .A2(_09460_),
    .B1(_10742_),
    .B2(_10748_),
    .X(_10749_));
 sky130_fd_sc_hd__inv_2 _14692_ (.A(_10749_),
    .Y(_01058_));
 sky130_fd_sc_hd__buf_4 _14693_ (.A(_10349_),
    .X(_10750_));
 sky130_fd_sc_hd__nand2_1 _14694_ (.A(_10750_),
    .B(net3033),
    .Y(_10751_));
 sky130_fd_sc_hd__a22o_1 _14695_ (.A1(_10739_),
    .A2(_09195_),
    .B1(_10742_),
    .B2(_10751_),
    .X(_10752_));
 sky130_fd_sc_hd__inv_2 _14696_ (.A(_10752_),
    .Y(_01059_));
 sky130_fd_sc_hd__nand2_1 _14697_ (.A(_10750_),
    .B(net3779),
    .Y(_10753_));
 sky130_fd_sc_hd__a22o_1 _14698_ (.A1(_10739_),
    .A2(_09201_),
    .B1(_10742_),
    .B2(_10753_),
    .X(_10754_));
 sky130_fd_sc_hd__inv_2 _14699_ (.A(_10754_),
    .Y(_01060_));
 sky130_fd_sc_hd__nand2_1 _14700_ (.A(_10750_),
    .B(net3571),
    .Y(_10755_));
 sky130_fd_sc_hd__a22o_1 _14701_ (.A1(_10739_),
    .A2(_09205_),
    .B1(_10742_),
    .B2(_10755_),
    .X(_10756_));
 sky130_fd_sc_hd__inv_2 _14702_ (.A(_10756_),
    .Y(_01061_));
 sky130_fd_sc_hd__nor2_1 _14703_ (.A(_09209_),
    .B(_10742_),
    .Y(_10757_));
 sky130_fd_sc_hd__a31o_1 _14704_ (.A1(_10703_),
    .A2(net2181),
    .A3(_10745_),
    .B1(_10757_),
    .X(_01062_));
 sky130_fd_sc_hd__and3_1 _14705_ (.A(_10736_),
    .B(_09326_),
    .C(_10687_),
    .X(_10758_));
 sky130_fd_sc_hd__a31o_1 _14706_ (.A1(_10745_),
    .A2(_10646_),
    .A3(net2520),
    .B1(_10758_),
    .X(_01063_));
 sky130_fd_sc_hd__buf_4 _14707_ (.A(_10279_),
    .X(_10759_));
 sky130_fd_sc_hd__clkbuf_16 _14708_ (.A(_09215_),
    .X(_10760_));
 sky130_fd_sc_hd__nor2_1 _14709_ (.A(_10760_),
    .B(_10742_),
    .Y(_10761_));
 sky130_fd_sc_hd__a31o_1 _14710_ (.A1(_10759_),
    .A2(net713),
    .A3(_10745_),
    .B1(_10761_),
    .X(_01048_));
 sky130_fd_sc_hd__nand2_1 _14711_ (.A(_10750_),
    .B(net3118),
    .Y(_10762_));
 sky130_fd_sc_hd__a22o_1 _14712_ (.A1(_10739_),
    .A2(_10122_),
    .B1(_10742_),
    .B2(_10762_),
    .X(_10763_));
 sky130_fd_sc_hd__inv_2 _14713_ (.A(_10763_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand2_1 _14714_ (.A(_10750_),
    .B(net2886),
    .Y(_10764_));
 sky130_fd_sc_hd__a22o_1 _14715_ (.A1(_10739_),
    .A2(_10195_),
    .B1(_10742_),
    .B2(_10764_),
    .X(_10765_));
 sky130_fd_sc_hd__inv_2 _14716_ (.A(_10765_),
    .Y(_01050_));
 sky130_fd_sc_hd__nor2_1 _14717_ (.A(_10657_),
    .B(_10742_),
    .Y(_10766_));
 sky130_fd_sc_hd__a31o_1 _14718_ (.A1(_10759_),
    .A2(net851),
    .A3(_10745_),
    .B1(_10766_),
    .X(_01051_));
 sky130_fd_sc_hd__clkbuf_16 _14719_ (.A(_09232_),
    .X(_10767_));
 sky130_fd_sc_hd__nor2_1 _14720_ (.A(_10767_),
    .B(_10742_),
    .Y(_10768_));
 sky130_fd_sc_hd__a31o_1 _14721_ (.A1(_10759_),
    .A2(net2092),
    .A3(_10745_),
    .B1(_10768_),
    .X(_01052_));
 sky130_fd_sc_hd__nor2_1 _14722_ (.A(_10602_),
    .B(_10742_),
    .Y(_10769_));
 sky130_fd_sc_hd__a31o_1 _14723_ (.A1(_10759_),
    .A2(net1813),
    .A3(_10745_),
    .B1(_10769_),
    .X(_01053_));
 sky130_fd_sc_hd__nand2_1 _14724_ (.A(_10750_),
    .B(net3361),
    .Y(_10770_));
 sky130_fd_sc_hd__a22o_1 _14725_ (.A1(_10739_),
    .A2(_10202_),
    .B1(_10742_),
    .B2(_10770_),
    .X(_10771_));
 sky130_fd_sc_hd__inv_2 _14726_ (.A(_10771_),
    .Y(_01054_));
 sky130_fd_sc_hd__nor2_1 _14727_ (.A(_10663_),
    .B(_10742_),
    .Y(_10772_));
 sky130_fd_sc_hd__a31o_1 _14728_ (.A1(_10759_),
    .A2(net963),
    .A3(_10745_),
    .B1(_10772_),
    .X(_01055_));
 sky130_fd_sc_hd__nand2_1 _14729_ (.A(_10750_),
    .B(net3387),
    .Y(_10773_));
 sky130_fd_sc_hd__a22o_1 _14730_ (.A1(_10739_),
    .A2(_09415_),
    .B1(_10741_),
    .B2(_10773_),
    .X(_10774_));
 sky130_fd_sc_hd__inv_2 _14731_ (.A(_10774_),
    .Y(_01040_));
 sky130_fd_sc_hd__and3_1 _14732_ (.A(_10736_),
    .B(_10667_),
    .C(_10687_),
    .X(_10775_));
 sky130_fd_sc_hd__a31o_1 _14733_ (.A1(_10745_),
    .A2(_10646_),
    .A3(net1981),
    .B1(_10775_),
    .X(_01041_));
 sky130_fd_sc_hd__nand2_1 _14734_ (.A(_10750_),
    .B(net3149),
    .Y(_10776_));
 sky130_fd_sc_hd__a22o_1 _14735_ (.A1(_10739_),
    .A2(_09348_),
    .B1(_10741_),
    .B2(_10776_),
    .X(_10777_));
 sky130_fd_sc_hd__inv_2 _14736_ (.A(_10777_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2_1 _14737_ (.A(_10750_),
    .B(net3471),
    .Y(_10778_));
 sky130_fd_sc_hd__a22o_1 _14738_ (.A1(_10739_),
    .A2(_09256_),
    .B1(_10741_),
    .B2(_10778_),
    .X(_10779_));
 sky130_fd_sc_hd__inv_2 _14739_ (.A(_10779_),
    .Y(_01043_));
 sky130_fd_sc_hd__nor2_1 _14740_ (.A(_09260_),
    .B(_10742_),
    .Y(_10780_));
 sky130_fd_sc_hd__a31o_1 _14741_ (.A1(_10759_),
    .A2(net2503),
    .A3(_10745_),
    .B1(_10780_),
    .X(_01044_));
 sky130_fd_sc_hd__nand2_1 _14742_ (.A(_10750_),
    .B(net2984),
    .Y(_10781_));
 sky130_fd_sc_hd__a22o_1 _14743_ (.A1(_10739_),
    .A2(_10149_),
    .B1(_10741_),
    .B2(_10781_),
    .X(_10782_));
 sky130_fd_sc_hd__inv_2 _14744_ (.A(_10782_),
    .Y(_01045_));
 sky130_fd_sc_hd__and3_1 _14745_ (.A(_10736_),
    .B(_10617_),
    .C(_10687_),
    .X(_10783_));
 sky130_fd_sc_hd__a31o_1 _14746_ (.A1(_10745_),
    .A2(_10646_),
    .A3(net2197),
    .B1(_10783_),
    .X(_01046_));
 sky130_fd_sc_hd__nand2_1 _14747_ (.A(_10750_),
    .B(net2925),
    .Y(_10784_));
 sky130_fd_sc_hd__a22o_1 _14748_ (.A1(_10739_),
    .A2(_10154_),
    .B1(_10741_),
    .B2(_10784_),
    .X(_10785_));
 sky130_fd_sc_hd__inv_2 _14749_ (.A(_10785_),
    .Y(_01047_));
 sky130_fd_sc_hd__nand2_1 _14750_ (.A(_10750_),
    .B(net3109),
    .Y(_10786_));
 sky130_fd_sc_hd__a22o_1 _14751_ (.A1(_10739_),
    .A2(_09495_),
    .B1(_10741_),
    .B2(_10786_),
    .X(_10787_));
 sky130_fd_sc_hd__inv_2 _14752_ (.A(_10787_),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_1 _14753_ (.A(_10750_),
    .B(net3452),
    .Y(_10788_));
 sky130_fd_sc_hd__a22o_1 _14754_ (.A1(_10739_),
    .A2(_09366_),
    .B1(_10741_),
    .B2(_10788_),
    .X(_10789_));
 sky130_fd_sc_hd__inv_2 _14755_ (.A(_10789_),
    .Y(_01033_));
 sky130_fd_sc_hd__and3_1 _14756_ (.A(_10736_),
    .B(_10728_),
    .C(_10687_),
    .X(_10790_));
 sky130_fd_sc_hd__a31o_1 _14757_ (.A1(_10745_),
    .A2(_10646_),
    .A3(net2060),
    .B1(_10790_),
    .X(_01034_));
 sky130_fd_sc_hd__nand2_1 _14758_ (.A(_10750_),
    .B(net3423),
    .Y(_10791_));
 sky130_fd_sc_hd__a22o_1 _14759_ (.A1(_10739_),
    .A2(_10164_),
    .B1(_10741_),
    .B2(_10791_),
    .X(_10792_));
 sky130_fd_sc_hd__inv_2 _14760_ (.A(_10792_),
    .Y(_01035_));
 sky130_fd_sc_hd__nand2_1 _14761_ (.A(_10750_),
    .B(net3575),
    .Y(_10793_));
 sky130_fd_sc_hd__a22o_1 _14762_ (.A1(_10738_),
    .A2(net139),
    .B1(_10741_),
    .B2(_10793_),
    .X(_10794_));
 sky130_fd_sc_hd__inv_2 _14763_ (.A(_10794_),
    .Y(_01036_));
 sky130_fd_sc_hd__and3_1 _14764_ (.A(_10736_),
    .B(_09730_),
    .C(_10687_),
    .X(_10795_));
 sky130_fd_sc_hd__a31o_1 _14765_ (.A1(_10745_),
    .A2(_10646_),
    .A3(net2162),
    .B1(_10795_),
    .X(_01037_));
 sky130_fd_sc_hd__nand2_1 _14766_ (.A(_10721_),
    .B(net3658),
    .Y(_10796_));
 sky130_fd_sc_hd__o2bb2a_1 _14767_ (.A1_N(_10796_),
    .A2_N(_10745_),
    .B1(_10289_),
    .B2(_10737_),
    .X(_01038_));
 sky130_fd_sc_hd__nor2_1 _14768_ (.A(_09300_),
    .B(_10742_),
    .Y(_10797_));
 sky130_fd_sc_hd__a31o_1 _14769_ (.A1(_10759_),
    .A2(net2405),
    .A3(_10745_),
    .B1(_10797_),
    .X(_01039_));
 sky130_fd_sc_hd__nor2_4 _14770_ (.A(_10691_),
    .B(_10356_),
    .Y(_10798_));
 sky130_fd_sc_hd__inv_2 _14771_ (.A(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__nor2_4 _14772_ (.A(_09190_),
    .B(_10799_),
    .Y(_10800_));
 sky130_fd_sc_hd__nor2_1 _14773_ (.A(_09625_),
    .B(_10799_),
    .Y(_10801_));
 sky130_fd_sc_hd__inv_2 _14774_ (.A(_10801_),
    .Y(_10802_));
 sky130_fd_sc_hd__buf_4 _14775_ (.A(_10802_),
    .X(_10803_));
 sky130_fd_sc_hd__nand2_1 _14776_ (.A(_10750_),
    .B(net3166),
    .Y(_10804_));
 sky130_fd_sc_hd__a22o_1 _14777_ (.A1(_10800_),
    .A2(_09451_),
    .B1(_10803_),
    .B2(_10804_),
    .X(_10805_));
 sky130_fd_sc_hd__inv_2 _14778_ (.A(_10805_),
    .Y(_01024_));
 sky130_fd_sc_hd__buf_4 _14779_ (.A(_10802_),
    .X(_10806_));
 sky130_fd_sc_hd__nor2_1 _14780_ (.A(_10746_),
    .B(_10803_),
    .Y(_10807_));
 sky130_fd_sc_hd__a31o_1 _14781_ (.A1(_10759_),
    .A2(net2392),
    .A3(_10806_),
    .B1(_10807_),
    .X(_01025_));
 sky130_fd_sc_hd__nor2_1 _14782_ (.A(_10698_),
    .B(_10803_),
    .Y(_10808_));
 sky130_fd_sc_hd__a31o_1 _14783_ (.A1(_10759_),
    .A2(net2634),
    .A3(_10806_),
    .B1(_10808_),
    .X(_01026_));
 sky130_fd_sc_hd__buf_4 _14784_ (.A(_10645_),
    .X(_10809_));
 sky130_fd_sc_hd__and3_1 _14785_ (.A(_10798_),
    .B(_09463_),
    .C(_10687_),
    .X(_10810_));
 sky130_fd_sc_hd__a31o_1 _14786_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net2552),
    .B1(_10810_),
    .X(_01027_));
 sky130_fd_sc_hd__and3_1 _14787_ (.A(_10798_),
    .B(_10587_),
    .C(_10687_),
    .X(_10811_));
 sky130_fd_sc_hd__a31o_1 _14788_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net1939),
    .B1(_10811_),
    .X(_01028_));
 sky130_fd_sc_hd__clkbuf_4 _14789_ (.A(_09359_),
    .X(_10812_));
 sky130_fd_sc_hd__and3_1 _14790_ (.A(_10798_),
    .B(_09395_),
    .C(_10812_),
    .X(_10813_));
 sky130_fd_sc_hd__a31o_1 _14791_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net2504),
    .B1(_10813_),
    .X(_01029_));
 sky130_fd_sc_hd__buf_4 _14792_ (.A(_10349_),
    .X(_10814_));
 sky130_fd_sc_hd__nand2_1 _14793_ (.A(_10814_),
    .B(net3866),
    .Y(_10815_));
 sky130_fd_sc_hd__a22o_1 _14794_ (.A1(_10800_),
    .A2(_09398_),
    .B1(_10803_),
    .B2(_10815_),
    .X(_10816_));
 sky130_fd_sc_hd__inv_2 _14795_ (.A(_10816_),
    .Y(_01030_));
 sky130_fd_sc_hd__and3_1 _14796_ (.A(_10798_),
    .B(_09326_),
    .C(_10812_),
    .X(_10817_));
 sky130_fd_sc_hd__a31o_1 _14797_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net1525),
    .B1(_10817_),
    .X(_01031_));
 sky130_fd_sc_hd__nor2_1 _14798_ (.A(_10760_),
    .B(_10803_),
    .Y(_10818_));
 sky130_fd_sc_hd__a31o_1 _14799_ (.A1(_10759_),
    .A2(net759),
    .A3(_10806_),
    .B1(_10818_),
    .X(_01016_));
 sky130_fd_sc_hd__nand2_1 _14800_ (.A(_10814_),
    .B(net2792),
    .Y(_10819_));
 sky130_fd_sc_hd__a22o_1 _14801_ (.A1(_10800_),
    .A2(_10122_),
    .B1(_10803_),
    .B2(_10819_),
    .X(_10820_));
 sky130_fd_sc_hd__inv_2 _14802_ (.A(_10820_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _14803_ (.A(_10814_),
    .B(net3117),
    .Y(_10821_));
 sky130_fd_sc_hd__a22o_1 _14804_ (.A1(_10800_),
    .A2(_10195_),
    .B1(_10803_),
    .B2(_10821_),
    .X(_10822_));
 sky130_fd_sc_hd__inv_2 _14805_ (.A(_10822_),
    .Y(_01018_));
 sky130_fd_sc_hd__nor2_1 _14806_ (.A(_10657_),
    .B(_10803_),
    .Y(_10823_));
 sky130_fd_sc_hd__a31o_1 _14807_ (.A1(_10759_),
    .A2(net455),
    .A3(_10806_),
    .B1(_10823_),
    .X(_01019_));
 sky130_fd_sc_hd__nor2_1 _14808_ (.A(_10767_),
    .B(_10803_),
    .Y(_10824_));
 sky130_fd_sc_hd__a31o_1 _14809_ (.A1(_10759_),
    .A2(net601),
    .A3(_10806_),
    .B1(_10824_),
    .X(_01020_));
 sky130_fd_sc_hd__nor2_1 _14810_ (.A(_10602_),
    .B(_10803_),
    .Y(_10825_));
 sky130_fd_sc_hd__a31o_1 _14811_ (.A1(_10759_),
    .A2(net449),
    .A3(_10803_),
    .B1(_10825_),
    .X(_01021_));
 sky130_fd_sc_hd__and3_1 _14812_ (.A(_10798_),
    .B(_09341_),
    .C(_10812_),
    .X(_10826_));
 sky130_fd_sc_hd__a31o_1 _14813_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net1837),
    .B1(_10826_),
    .X(_01022_));
 sky130_fd_sc_hd__nor2_1 _14814_ (.A(_10663_),
    .B(_10803_),
    .Y(_10827_));
 sky130_fd_sc_hd__a31o_1 _14815_ (.A1(_10759_),
    .A2(net421),
    .A3(_10803_),
    .B1(_10827_),
    .X(_01023_));
 sky130_fd_sc_hd__nand2_1 _14816_ (.A(_10814_),
    .B(net2968),
    .Y(_10828_));
 sky130_fd_sc_hd__a22o_1 _14817_ (.A1(_10800_),
    .A2(net137),
    .B1(_10803_),
    .B2(_10828_),
    .X(_10829_));
 sky130_fd_sc_hd__inv_2 _14818_ (.A(_10829_),
    .Y(_01008_));
 sky130_fd_sc_hd__and3_1 _14819_ (.A(_10798_),
    .B(_10667_),
    .C(_10812_),
    .X(_10830_));
 sky130_fd_sc_hd__a31o_1 _14820_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net555),
    .B1(_10830_),
    .X(_01009_));
 sky130_fd_sc_hd__nand2_1 _14821_ (.A(_10814_),
    .B(net3211),
    .Y(_10831_));
 sky130_fd_sc_hd__a22o_1 _14822_ (.A1(_10800_),
    .A2(_09348_),
    .B1(_10802_),
    .B2(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__inv_2 _14823_ (.A(_10832_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_1 _14824_ (.A(_10814_),
    .B(net2883),
    .Y(_10833_));
 sky130_fd_sc_hd__a22o_1 _14825_ (.A1(_10800_),
    .A2(_09256_),
    .B1(_10802_),
    .B2(_10833_),
    .X(_10834_));
 sky130_fd_sc_hd__inv_2 _14826_ (.A(_10834_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand2_1 _14827_ (.A(_10814_),
    .B(net3073),
    .Y(_10835_));
 sky130_fd_sc_hd__a22o_1 _14828_ (.A1(_10800_),
    .A2(_09354_),
    .B1(_10802_),
    .B2(_10835_),
    .X(_10836_));
 sky130_fd_sc_hd__inv_2 _14829_ (.A(_10836_),
    .Y(_01012_));
 sky130_fd_sc_hd__nand2_1 _14830_ (.A(_10814_),
    .B(net3120),
    .Y(_10837_));
 sky130_fd_sc_hd__a22o_1 _14831_ (.A1(_10800_),
    .A2(_10149_),
    .B1(_10802_),
    .B2(_10837_),
    .X(_10838_));
 sky130_fd_sc_hd__inv_2 _14832_ (.A(_10838_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _14833_ (.A(_10814_),
    .B(net2774),
    .Y(_10839_));
 sky130_fd_sc_hd__a22o_1 _14834_ (.A1(_10800_),
    .A2(_09425_),
    .B1(_10802_),
    .B2(_10839_),
    .X(_10840_));
 sky130_fd_sc_hd__inv_2 _14835_ (.A(_10840_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _14836_ (.A(_10814_),
    .B(net2835),
    .Y(_10841_));
 sky130_fd_sc_hd__a22o_1 _14837_ (.A1(_10800_),
    .A2(_10154_),
    .B1(_10802_),
    .B2(_10841_),
    .X(_10842_));
 sky130_fd_sc_hd__inv_2 _14838_ (.A(_10842_),
    .Y(_01015_));
 sky130_fd_sc_hd__and3_1 _14839_ (.A(_10798_),
    .B(_10679_),
    .C(_10812_),
    .X(_10843_));
 sky130_fd_sc_hd__a31o_1 _14840_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net547),
    .B1(_10843_),
    .X(_01000_));
 sky130_fd_sc_hd__nor2_1 _14841_ (.A(_10681_),
    .B(_10803_),
    .Y(_10844_));
 sky130_fd_sc_hd__a31o_1 _14842_ (.A1(_10759_),
    .A2(net1155),
    .A3(_10803_),
    .B1(_10844_),
    .X(_01001_));
 sky130_fd_sc_hd__and3_1 _14843_ (.A(_10798_),
    .B(_10728_),
    .C(_10812_),
    .X(_10845_));
 sky130_fd_sc_hd__a31o_1 _14844_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net533),
    .B1(_10845_),
    .X(_01002_));
 sky130_fd_sc_hd__nand2_1 _14845_ (.A(_10814_),
    .B(net2769),
    .Y(_10846_));
 sky130_fd_sc_hd__a22o_1 _14846_ (.A1(_10800_),
    .A2(_10164_),
    .B1(_10802_),
    .B2(_10846_),
    .X(_10847_));
 sky130_fd_sc_hd__inv_2 _14847_ (.A(_10847_),
    .Y(_01003_));
 sky130_fd_sc_hd__buf_12 _14848_ (.A(net77),
    .X(_10848_));
 sky130_fd_sc_hd__and3_1 _14849_ (.A(_10798_),
    .B(_10848_),
    .C(_10812_),
    .X(_10849_));
 sky130_fd_sc_hd__a31o_1 _14850_ (.A1(_10806_),
    .A2(_10809_),
    .A3(net579),
    .B1(_10849_),
    .X(_01004_));
 sky130_fd_sc_hd__nand2_1 _14851_ (.A(_10814_),
    .B(net2880),
    .Y(_10850_));
 sky130_fd_sc_hd__a22o_1 _14852_ (.A1(_10800_),
    .A2(_09504_),
    .B1(_10802_),
    .B2(_10850_),
    .X(_10851_));
 sky130_fd_sc_hd__inv_2 _14853_ (.A(_10851_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _14854_ (.A(_10721_),
    .B(net3300),
    .Y(_10852_));
 sky130_fd_sc_hd__o2bb2a_1 _14855_ (.A1_N(_10852_),
    .A2_N(_10806_),
    .B1(_10289_),
    .B2(_10799_),
    .X(_01006_));
 sky130_fd_sc_hd__nand2_1 _14856_ (.A(_10721_),
    .B(net3547),
    .Y(_10853_));
 sky130_fd_sc_hd__o2bb2a_1 _14857_ (.A1_N(_10853_),
    .A2_N(_10806_),
    .B1(_09442_),
    .B2(_10799_),
    .X(_01007_));
 sky130_fd_sc_hd__nor2_4 _14858_ (.A(_10691_),
    .B(_10411_),
    .Y(_10854_));
 sky130_fd_sc_hd__inv_2 _14859_ (.A(_10854_),
    .Y(_10855_));
 sky130_fd_sc_hd__nor2_4 _14860_ (.A(_08795_),
    .B(_10855_),
    .Y(_10856_));
 sky130_fd_sc_hd__nor2_1 _14861_ (.A(_09304_),
    .B(_10855_),
    .Y(_10857_));
 sky130_fd_sc_hd__inv_2 _14862_ (.A(_10857_),
    .Y(_10858_));
 sky130_fd_sc_hd__buf_4 _14863_ (.A(_10858_),
    .X(_10859_));
 sky130_fd_sc_hd__nand2_1 _14864_ (.A(_10814_),
    .B(net3497),
    .Y(_10860_));
 sky130_fd_sc_hd__a22o_1 _14865_ (.A1(_10856_),
    .A2(_10239_),
    .B1(_10859_),
    .B2(_10860_),
    .X(_10861_));
 sky130_fd_sc_hd__inv_2 _14866_ (.A(_10861_),
    .Y(_00992_));
 sky130_fd_sc_hd__buf_4 _14867_ (.A(_10858_),
    .X(_10862_));
 sky130_fd_sc_hd__nor2_1 _14868_ (.A(_10746_),
    .B(_10859_),
    .Y(_10863_));
 sky130_fd_sc_hd__a31o_1 _14869_ (.A1(_10759_),
    .A2(net445),
    .A3(_10862_),
    .B1(_10863_),
    .X(_00993_));
 sky130_fd_sc_hd__buf_4 _14870_ (.A(_08776_),
    .X(_10864_));
 sky130_fd_sc_hd__buf_4 _14871_ (.A(_10864_),
    .X(_10865_));
 sky130_fd_sc_hd__nor2_1 _14872_ (.A(_10698_),
    .B(_10859_),
    .Y(_10866_));
 sky130_fd_sc_hd__a31o_1 _14873_ (.A1(_10865_),
    .A2(net1233),
    .A3(_10862_),
    .B1(_10866_),
    .X(_00994_));
 sky130_fd_sc_hd__and3_1 _14874_ (.A(_10854_),
    .B(_09463_),
    .C(_10812_),
    .X(_10867_));
 sky130_fd_sc_hd__a31o_1 _14875_ (.A1(_10862_),
    .A2(_10809_),
    .A3(net1053),
    .B1(_10867_),
    .X(_00995_));
 sky130_fd_sc_hd__and3_1 _14876_ (.A(_10854_),
    .B(_10587_),
    .C(_10812_),
    .X(_10868_));
 sky130_fd_sc_hd__a31o_1 _14877_ (.A1(_10862_),
    .A2(_10809_),
    .A3(net719),
    .B1(_10868_),
    .X(_00996_));
 sky130_fd_sc_hd__clkbuf_16 _14878_ (.A(_09204_),
    .X(_10869_));
 sky130_fd_sc_hd__nand2_1 _14879_ (.A(_10814_),
    .B(net3704),
    .Y(_10870_));
 sky130_fd_sc_hd__a22o_1 _14880_ (.A1(_10856_),
    .A2(_10869_),
    .B1(_10859_),
    .B2(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__inv_2 _14881_ (.A(_10871_),
    .Y(_00997_));
 sky130_fd_sc_hd__clkbuf_16 _14882_ (.A(_09208_),
    .X(_10872_));
 sky130_fd_sc_hd__nor2_1 _14883_ (.A(_10872_),
    .B(_10859_),
    .Y(_10873_));
 sky130_fd_sc_hd__a31o_1 _14884_ (.A1(_10865_),
    .A2(net465),
    .A3(_10862_),
    .B1(_10873_),
    .X(_00998_));
 sky130_fd_sc_hd__clkbuf_16 _14885_ (.A(net74),
    .X(_10874_));
 sky130_fd_sc_hd__and3_1 _14886_ (.A(_10854_),
    .B(_10874_),
    .C(_10812_),
    .X(_10875_));
 sky130_fd_sc_hd__a31o_1 _14887_ (.A1(_10862_),
    .A2(_10809_),
    .A3(net559),
    .B1(_10875_),
    .X(_00999_));
 sky130_fd_sc_hd__nor2_1 _14888_ (.A(_10760_),
    .B(_10859_),
    .Y(_10876_));
 sky130_fd_sc_hd__a31o_1 _14889_ (.A1(_10865_),
    .A2(net1977),
    .A3(_10862_),
    .B1(_10876_),
    .X(_00984_));
 sky130_fd_sc_hd__nand2_1 _14890_ (.A(_10814_),
    .B(net3224),
    .Y(_10877_));
 sky130_fd_sc_hd__a22o_1 _14891_ (.A1(_10856_),
    .A2(_10122_),
    .B1(_10858_),
    .B2(_10877_),
    .X(_10878_));
 sky130_fd_sc_hd__inv_2 _14892_ (.A(_10878_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _14893_ (.A(_10814_),
    .B(net3081),
    .Y(_10879_));
 sky130_fd_sc_hd__a22o_1 _14894_ (.A1(_10856_),
    .A2(_10195_),
    .B1(_10858_),
    .B2(_10879_),
    .X(_10880_));
 sky130_fd_sc_hd__inv_2 _14895_ (.A(_10880_),
    .Y(_00986_));
 sky130_fd_sc_hd__nor2_1 _14896_ (.A(_10657_),
    .B(_10859_),
    .Y(_10881_));
 sky130_fd_sc_hd__a31o_1 _14897_ (.A1(_10865_),
    .A2(net2529),
    .A3(_10859_),
    .B1(_10881_),
    .X(_00987_));
 sky130_fd_sc_hd__nor2_1 _14898_ (.A(_10767_),
    .B(_10859_),
    .Y(_10882_));
 sky130_fd_sc_hd__a31o_1 _14899_ (.A1(_10865_),
    .A2(net1075),
    .A3(_10859_),
    .B1(_10882_),
    .X(_00988_));
 sky130_fd_sc_hd__nor2_1 _14900_ (.A(_10602_),
    .B(_10859_),
    .Y(_10883_));
 sky130_fd_sc_hd__a31o_1 _14901_ (.A1(_10865_),
    .A2(net1962),
    .A3(_10859_),
    .B1(_10883_),
    .X(_00989_));
 sky130_fd_sc_hd__buf_4 _14902_ (.A(_10349_),
    .X(_10884_));
 sky130_fd_sc_hd__nand2_1 _14903_ (.A(_10884_),
    .B(net3752),
    .Y(_10885_));
 sky130_fd_sc_hd__a22o_1 _14904_ (.A1(_10856_),
    .A2(_10202_),
    .B1(_10858_),
    .B2(_10885_),
    .X(_10886_));
 sky130_fd_sc_hd__inv_2 _14905_ (.A(_10886_),
    .Y(_00990_));
 sky130_fd_sc_hd__nor2_1 _14906_ (.A(_10663_),
    .B(_10859_),
    .Y(_10887_));
 sky130_fd_sc_hd__a31o_1 _14907_ (.A1(_10865_),
    .A2(net1959),
    .A3(_10859_),
    .B1(_10887_),
    .X(_00991_));
 sky130_fd_sc_hd__nor2_1 _14908_ (.A(_09246_),
    .B(_10859_),
    .Y(_10888_));
 sky130_fd_sc_hd__a31o_1 _14909_ (.A1(_10865_),
    .A2(net1439),
    .A3(_10859_),
    .B1(_10888_),
    .X(_00968_));
 sky130_fd_sc_hd__and3_1 _14910_ (.A(_10854_),
    .B(_10667_),
    .C(_10812_),
    .X(_10889_));
 sky130_fd_sc_hd__a31o_1 _14911_ (.A1(_10862_),
    .A2(_10809_),
    .A3(net2451),
    .B1(_10889_),
    .X(_00969_));
 sky130_fd_sc_hd__nand2_1 _14912_ (.A(_10884_),
    .B(net3405),
    .Y(_10890_));
 sky130_fd_sc_hd__a22o_1 _14913_ (.A1(_10856_),
    .A2(_09348_),
    .B1(_10858_),
    .B2(_10890_),
    .X(_10891_));
 sky130_fd_sc_hd__inv_2 _14914_ (.A(_10891_),
    .Y(_00970_));
 sky130_fd_sc_hd__and3_1 _14915_ (.A(_10854_),
    .B(_10500_),
    .C(_10812_),
    .X(_10892_));
 sky130_fd_sc_hd__a31o_1 _14916_ (.A1(_10862_),
    .A2(_10809_),
    .A3(net2487),
    .B1(_10892_),
    .X(_00971_));
 sky130_fd_sc_hd__nand2_1 _14917_ (.A(_10884_),
    .B(net3174),
    .Y(_10893_));
 sky130_fd_sc_hd__a22o_1 _14918_ (.A1(_10856_),
    .A2(_09354_),
    .B1(_10858_),
    .B2(_10893_),
    .X(_10894_));
 sky130_fd_sc_hd__inv_2 _14919_ (.A(_10894_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_1 _14920_ (.A(_10884_),
    .B(net3335),
    .Y(_10895_));
 sky130_fd_sc_hd__a22o_1 _14921_ (.A1(_10856_),
    .A2(_10149_),
    .B1(_10858_),
    .B2(_10895_),
    .X(_10896_));
 sky130_fd_sc_hd__inv_2 _14922_ (.A(_10896_),
    .Y(_00973_));
 sky130_fd_sc_hd__and3_1 _14923_ (.A(_10854_),
    .B(_10617_),
    .C(_10812_),
    .X(_10897_));
 sky130_fd_sc_hd__a31o_1 _14924_ (.A1(_10862_),
    .A2(_10809_),
    .A3(net1817),
    .B1(_10897_),
    .X(_00974_));
 sky130_fd_sc_hd__nand2_1 _14925_ (.A(_10884_),
    .B(net3739),
    .Y(_10898_));
 sky130_fd_sc_hd__a22o_1 _14926_ (.A1(_10856_),
    .A2(_10154_),
    .B1(_10858_),
    .B2(_10898_),
    .X(_10899_));
 sky130_fd_sc_hd__inv_2 _14927_ (.A(_10899_),
    .Y(_00975_));
 sky130_fd_sc_hd__and3_1 _14928_ (.A(_10854_),
    .B(_10679_),
    .C(_10812_),
    .X(_10900_));
 sky130_fd_sc_hd__a31o_1 _14929_ (.A1(_10862_),
    .A2(_10809_),
    .A3(net1943),
    .B1(_10900_),
    .X(_00960_));
 sky130_fd_sc_hd__nand2_1 _14930_ (.A(_10884_),
    .B(net3595),
    .Y(_10901_));
 sky130_fd_sc_hd__a22o_1 _14931_ (.A1(_10856_),
    .A2(_09366_),
    .B1(_10858_),
    .B2(_10901_),
    .X(_10902_));
 sky130_fd_sc_hd__inv_2 _14932_ (.A(_10902_),
    .Y(_00961_));
 sky130_fd_sc_hd__clkbuf_8 _14933_ (.A(_10645_),
    .X(_10903_));
 sky130_fd_sc_hd__and3_1 _14934_ (.A(_10854_),
    .B(_10728_),
    .C(_10812_),
    .X(_10904_));
 sky130_fd_sc_hd__a31o_1 _14935_ (.A1(_10862_),
    .A2(_10903_),
    .A3(net2323),
    .B1(_10904_),
    .X(_00962_));
 sky130_fd_sc_hd__nand2_1 _14936_ (.A(_10884_),
    .B(net3578),
    .Y(_10905_));
 sky130_fd_sc_hd__a22o_1 _14937_ (.A1(_10856_),
    .A2(_10164_),
    .B1(_10858_),
    .B2(_10905_),
    .X(_10906_));
 sky130_fd_sc_hd__inv_2 _14938_ (.A(_10906_),
    .Y(_00963_));
 sky130_fd_sc_hd__and3_1 _14939_ (.A(_10854_),
    .B(_10848_),
    .C(_10812_),
    .X(_10907_));
 sky130_fd_sc_hd__a31o_1 _14940_ (.A1(_10862_),
    .A2(_10903_),
    .A3(net1682),
    .B1(_10907_),
    .X(_00964_));
 sky130_fd_sc_hd__buf_4 _14941_ (.A(_09359_),
    .X(_10908_));
 sky130_fd_sc_hd__and3_1 _14942_ (.A(_10854_),
    .B(_09730_),
    .C(_10908_),
    .X(_10909_));
 sky130_fd_sc_hd__a31o_1 _14943_ (.A1(_10862_),
    .A2(_10903_),
    .A3(net1425),
    .B1(_10909_),
    .X(_00965_));
 sky130_fd_sc_hd__nand2_1 _14944_ (.A(_10721_),
    .B(net4016),
    .Y(_10910_));
 sky130_fd_sc_hd__o2bb2a_1 _14945_ (.A1_N(_10910_),
    .A2_N(_10862_),
    .B1(_10289_),
    .B2(_10855_),
    .X(_00966_));
 sky130_fd_sc_hd__nand2_1 _14946_ (.A(_10721_),
    .B(net3832),
    .Y(_10911_));
 sky130_fd_sc_hd__o2bb2a_1 _14947_ (.A1_N(_10911_),
    .A2_N(_10862_),
    .B1(_09442_),
    .B2(_10855_),
    .X(_00967_));
 sky130_fd_sc_hd__nand2_4 _14948_ (.A(_10466_),
    .B(_09982_),
    .Y(_10912_));
 sky130_fd_sc_hd__nor2_4 _14949_ (.A(_10912_),
    .B(_10469_),
    .Y(_10913_));
 sky130_fd_sc_hd__nand2_4 _14950_ (.A(_10913_),
    .B(_10413_),
    .Y(_10914_));
 sky130_fd_sc_hd__buf_4 _14951_ (.A(_10914_),
    .X(_10915_));
 sky130_fd_sc_hd__nor2_1 _14952_ (.A(_09181_),
    .B(_10915_),
    .Y(_10916_));
 sky130_fd_sc_hd__a31o_1 _14953_ (.A1(_10865_),
    .A2(net2190),
    .A3(_10915_),
    .B1(_10916_),
    .X(_00952_));
 sky130_fd_sc_hd__buf_4 _14954_ (.A(_10914_),
    .X(_10917_));
 sky130_fd_sc_hd__nor2_1 _14955_ (.A(_10746_),
    .B(_10917_),
    .Y(_10918_));
 sky130_fd_sc_hd__a31o_1 _14956_ (.A1(_10865_),
    .A2(net2471),
    .A3(_10915_),
    .B1(_10918_),
    .X(_00953_));
 sky130_fd_sc_hd__nor2_1 _14957_ (.A(_10698_),
    .B(_10917_),
    .Y(_10919_));
 sky130_fd_sc_hd__a31o_1 _14958_ (.A1(_10865_),
    .A2(net2473),
    .A3(_10915_),
    .B1(_10919_),
    .X(_00954_));
 sky130_fd_sc_hd__and3_1 _14959_ (.A(_10913_),
    .B(_09463_),
    .C(_10908_),
    .X(_10920_));
 sky130_fd_sc_hd__a31o_1 _14960_ (.A1(_10865_),
    .A2(net2335),
    .A3(_10915_),
    .B1(_10920_),
    .X(_00955_));
 sky130_fd_sc_hd__and3_1 _14961_ (.A(_10913_),
    .B(_10587_),
    .C(_10908_),
    .X(_10921_));
 sky130_fd_sc_hd__a31o_1 _14962_ (.A1(_10865_),
    .A2(net2001),
    .A3(_10915_),
    .B1(_10921_),
    .X(_00956_));
 sky130_fd_sc_hd__nand2_1 _14963_ (.A(_10395_),
    .B(net4169),
    .Y(_10922_));
 sky130_fd_sc_hd__and2_1 _14964_ (.A(_10913_),
    .B(_08778_),
    .X(_10923_));
 sky130_fd_sc_hd__buf_4 _14965_ (.A(_10923_),
    .X(_10924_));
 sky130_fd_sc_hd__a22o_1 _14966_ (.A1(_10917_),
    .A2(_10922_),
    .B1(_10924_),
    .B2(_09205_),
    .X(_10925_));
 sky130_fd_sc_hd__inv_2 _14967_ (.A(_10925_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_1 _14968_ (.A(_10395_),
    .B(net4118),
    .Y(_10926_));
 sky130_fd_sc_hd__a22o_1 _14969_ (.A1(_10917_),
    .A2(_10926_),
    .B1(_10924_),
    .B2(_09398_),
    .X(_10927_));
 sky130_fd_sc_hd__inv_2 _14970_ (.A(_10927_),
    .Y(_00958_));
 sky130_fd_sc_hd__and3_1 _14971_ (.A(_10913_),
    .B(_10874_),
    .C(_10908_),
    .X(_10928_));
 sky130_fd_sc_hd__a31o_1 _14972_ (.A1(_10865_),
    .A2(net2079),
    .A3(_10915_),
    .B1(_10928_),
    .X(_00959_));
 sky130_fd_sc_hd__nor2_1 _14973_ (.A(_10760_),
    .B(_10917_),
    .Y(_10929_));
 sky130_fd_sc_hd__a31o_1 _14974_ (.A1(_10865_),
    .A2(net495),
    .A3(_10915_),
    .B1(_10929_),
    .X(_00944_));
 sky130_fd_sc_hd__buf_4 _14975_ (.A(_08775_),
    .X(_10930_));
 sky130_fd_sc_hd__clkbuf_8 _14976_ (.A(_10930_),
    .X(_10931_));
 sky130_fd_sc_hd__nand2_1 _14977_ (.A(_10931_),
    .B(net4175),
    .Y(_10932_));
 sky130_fd_sc_hd__a22o_1 _14978_ (.A1(_10917_),
    .A2(_10932_),
    .B1(_10924_),
    .B2(_10313_),
    .X(_10933_));
 sky130_fd_sc_hd__inv_2 _14979_ (.A(_10933_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _14980_ (.A(_10931_),
    .B(net4144),
    .Y(_10934_));
 sky130_fd_sc_hd__a22o_1 _14981_ (.A1(_10917_),
    .A2(_10934_),
    .B1(_10924_),
    .B2(_10316_),
    .X(_10935_));
 sky130_fd_sc_hd__inv_2 _14982_ (.A(_10935_),
    .Y(_00946_));
 sky130_fd_sc_hd__nor2_1 _14983_ (.A(_10657_),
    .B(_10917_),
    .Y(_10936_));
 sky130_fd_sc_hd__a31o_1 _14984_ (.A1(_10865_),
    .A2(net823),
    .A3(_10915_),
    .B1(_10936_),
    .X(_00947_));
 sky130_fd_sc_hd__buf_4 _14985_ (.A(_10864_),
    .X(_10937_));
 sky130_fd_sc_hd__nor2_1 _14986_ (.A(_10767_),
    .B(_10917_),
    .Y(_10938_));
 sky130_fd_sc_hd__a31o_1 _14987_ (.A1(_10937_),
    .A2(net529),
    .A3(_10915_),
    .B1(_10938_),
    .X(_00948_));
 sky130_fd_sc_hd__nor2_1 _14988_ (.A(_10602_),
    .B(_10917_),
    .Y(_10939_));
 sky130_fd_sc_hd__a31o_1 _14989_ (.A1(_10937_),
    .A2(net981),
    .A3(_10915_),
    .B1(_10939_),
    .X(_00949_));
 sky130_fd_sc_hd__nand2_1 _14990_ (.A(_10931_),
    .B(net3861),
    .Y(_10940_));
 sky130_fd_sc_hd__a22o_1 _14991_ (.A1(_10917_),
    .A2(_10940_),
    .B1(_10924_),
    .B2(_09239_),
    .X(_10941_));
 sky130_fd_sc_hd__inv_2 _14992_ (.A(_10941_),
    .Y(_00950_));
 sky130_fd_sc_hd__nor2_1 _14993_ (.A(_10663_),
    .B(_10917_),
    .Y(_10942_));
 sky130_fd_sc_hd__a31o_1 _14994_ (.A1(_10937_),
    .A2(net997),
    .A3(_10915_),
    .B1(_10942_),
    .X(_00951_));
 sky130_fd_sc_hd__nand2_1 _14995_ (.A(_10931_),
    .B(net4115),
    .Y(_10943_));
 sky130_fd_sc_hd__a22o_1 _14996_ (.A1(_10914_),
    .A2(_10943_),
    .B1(_10924_),
    .B2(_09415_),
    .X(_10944_));
 sky130_fd_sc_hd__inv_2 _14997_ (.A(_10944_),
    .Y(_00936_));
 sky130_fd_sc_hd__and3_1 _14998_ (.A(_10913_),
    .B(_10667_),
    .C(_10908_),
    .X(_10945_));
 sky130_fd_sc_hd__a31o_1 _14999_ (.A1(_10937_),
    .A2(net2113),
    .A3(_10915_),
    .B1(_10945_),
    .X(_00937_));
 sky130_fd_sc_hd__nor2_1 _15000_ (.A(_10669_),
    .B(_10917_),
    .Y(_10946_));
 sky130_fd_sc_hd__a31o_1 _15001_ (.A1(_10937_),
    .A2(net1455),
    .A3(_10915_),
    .B1(_10946_),
    .X(_00938_));
 sky130_fd_sc_hd__and3_1 _15002_ (.A(_10913_),
    .B(_10500_),
    .C(_10908_),
    .X(_10947_));
 sky130_fd_sc_hd__a31o_1 _15003_ (.A1(_10937_),
    .A2(net1057),
    .A3(_10915_),
    .B1(_10947_),
    .X(_00939_));
 sky130_fd_sc_hd__nor2_1 _15004_ (.A(_09260_),
    .B(_10917_),
    .Y(_10948_));
 sky130_fd_sc_hd__a31o_1 _15005_ (.A1(_10937_),
    .A2(net2146),
    .A3(_10915_),
    .B1(_10948_),
    .X(_00940_));
 sky130_fd_sc_hd__nand2_1 _15006_ (.A(_10931_),
    .B(net4280),
    .Y(_10949_));
 sky130_fd_sc_hd__a22o_1 _15007_ (.A1(_10914_),
    .A2(_10949_),
    .B1(_10924_),
    .B2(_10331_),
    .X(_10950_));
 sky130_fd_sc_hd__inv_2 _15008_ (.A(_10950_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_1 _15009_ (.A(_10931_),
    .B(net3994),
    .Y(_10951_));
 sky130_fd_sc_hd__a22o_1 _15010_ (.A1(_10914_),
    .A2(_10951_),
    .B1(_10924_),
    .B2(_09425_),
    .X(_10952_));
 sky130_fd_sc_hd__inv_2 _15011_ (.A(_10952_),
    .Y(_00942_));
 sky130_fd_sc_hd__nand2_1 _15012_ (.A(_10931_),
    .B(net4263),
    .Y(_10953_));
 sky130_fd_sc_hd__a22o_1 _15013_ (.A1(_10914_),
    .A2(_10953_),
    .B1(_10924_),
    .B2(_10335_),
    .X(_10954_));
 sky130_fd_sc_hd__inv_2 _15014_ (.A(_10954_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _15015_ (.A(_10931_),
    .B(net3955),
    .Y(_10955_));
 sky130_fd_sc_hd__a22o_1 _15016_ (.A1(_10914_),
    .A2(_10955_),
    .B1(_10924_),
    .B2(_09495_),
    .X(_10956_));
 sky130_fd_sc_hd__inv_2 _15017_ (.A(_10956_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _15018_ (.A(_10931_),
    .B(net3892),
    .Y(_10957_));
 sky130_fd_sc_hd__a22o_1 _15019_ (.A1(_10914_),
    .A2(_10957_),
    .B1(_10924_),
    .B2(_09366_),
    .X(_10958_));
 sky130_fd_sc_hd__inv_2 _15020_ (.A(_10958_),
    .Y(_00929_));
 sky130_fd_sc_hd__nand2_1 _15021_ (.A(_10931_),
    .B(net3890),
    .Y(_10959_));
 sky130_fd_sc_hd__a22o_1 _15022_ (.A1(_10914_),
    .A2(_10959_),
    .B1(_10924_),
    .B2(_09280_),
    .X(_10960_));
 sky130_fd_sc_hd__inv_2 _15023_ (.A(_10960_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _15024_ (.A(_10931_),
    .B(net3989),
    .Y(_10961_));
 sky130_fd_sc_hd__a22o_1 _15025_ (.A1(_10914_),
    .A2(_10961_),
    .B1(_10924_),
    .B2(_10342_),
    .X(_10962_));
 sky130_fd_sc_hd__inv_2 _15026_ (.A(_10962_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _15027_ (.A(_10931_),
    .B(net3941),
    .Y(_10963_));
 sky130_fd_sc_hd__a22o_1 _15028_ (.A1(_10914_),
    .A2(_10963_),
    .B1(_10924_),
    .B2(_09288_),
    .X(_10964_));
 sky130_fd_sc_hd__inv_2 _15029_ (.A(_10964_),
    .Y(_00932_));
 sky130_fd_sc_hd__nand2_1 _15030_ (.A(_10931_),
    .B(net3980),
    .Y(_10965_));
 sky130_fd_sc_hd__a22o_1 _15031_ (.A1(_10914_),
    .A2(_10965_),
    .B1(_10924_),
    .B2(_09504_),
    .X(_10966_));
 sky130_fd_sc_hd__inv_2 _15032_ (.A(_10966_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_1 _15033_ (.A(_10884_),
    .B(net2868),
    .Y(_10967_));
 sky130_fd_sc_hd__a22o_1 _15034_ (.A1(_10348_),
    .A2(_10913_),
    .B1(_10917_),
    .B2(_10967_),
    .X(_10968_));
 sky130_fd_sc_hd__inv_2 _15035_ (.A(net2869),
    .Y(_00934_));
 sky130_fd_sc_hd__nand2_1 _15036_ (.A(_10884_),
    .B(net2859),
    .Y(_10969_));
 sky130_fd_sc_hd__a22o_1 _15037_ (.A1(net142),
    .A2(_10913_),
    .B1(_10917_),
    .B2(_10969_),
    .X(_10970_));
 sky130_fd_sc_hd__inv_2 _15038_ (.A(net2860),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_2 _15039_ (.A(_10912_),
    .B(_10292_),
    .Y(_10971_));
 sky130_fd_sc_hd__inv_2 _15040_ (.A(_10971_),
    .Y(_10972_));
 sky130_fd_sc_hd__nor2_4 _15041_ (.A(_08797_),
    .B(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__nor2_1 _15042_ (.A(_09304_),
    .B(_10972_),
    .Y(_10974_));
 sky130_fd_sc_hd__inv_2 _15043_ (.A(_10974_),
    .Y(_10975_));
 sky130_fd_sc_hd__buf_4 _15044_ (.A(_10975_),
    .X(_10976_));
 sky130_fd_sc_hd__nand2_1 _15045_ (.A(_10884_),
    .B(net3851),
    .Y(_10977_));
 sky130_fd_sc_hd__a22o_1 _15046_ (.A1(_10973_),
    .A2(_10239_),
    .B1(_10976_),
    .B2(_10977_),
    .X(_10978_));
 sky130_fd_sc_hd__inv_2 _15047_ (.A(_10978_),
    .Y(_00920_));
 sky130_fd_sc_hd__buf_4 _15048_ (.A(_10975_),
    .X(_10979_));
 sky130_fd_sc_hd__nor2_1 _15049_ (.A(_10746_),
    .B(_10976_),
    .Y(_10980_));
 sky130_fd_sc_hd__a31o_1 _15050_ (.A1(_10937_),
    .A2(net703),
    .A3(_10979_),
    .B1(_10980_),
    .X(_00921_));
 sky130_fd_sc_hd__nand2_1 _15051_ (.A(_10884_),
    .B(net3448),
    .Y(_10981_));
 sky130_fd_sc_hd__a22o_1 _15052_ (.A1(_10973_),
    .A2(_09460_),
    .B1(_10976_),
    .B2(_10981_),
    .X(_10982_));
 sky130_fd_sc_hd__inv_2 _15053_ (.A(_10982_),
    .Y(_00922_));
 sky130_fd_sc_hd__buf_12 _15054_ (.A(_09194_),
    .X(_10983_));
 sky130_fd_sc_hd__nand2_1 _15055_ (.A(_10884_),
    .B(net2939),
    .Y(_10984_));
 sky130_fd_sc_hd__a22o_1 _15056_ (.A1(_10973_),
    .A2(_10983_),
    .B1(_10976_),
    .B2(_10984_),
    .X(_10985_));
 sky130_fd_sc_hd__inv_2 _15057_ (.A(_10985_),
    .Y(_00923_));
 sky130_fd_sc_hd__and3_1 _15058_ (.A(_10971_),
    .B(_10587_),
    .C(_10908_),
    .X(_10986_));
 sky130_fd_sc_hd__a31o_1 _15059_ (.A1(_10979_),
    .A2(_10903_),
    .A3(net1293),
    .B1(_10986_),
    .X(_00924_));
 sky130_fd_sc_hd__nand2_1 _15060_ (.A(_10884_),
    .B(net3736),
    .Y(_10987_));
 sky130_fd_sc_hd__a22o_1 _15061_ (.A1(_10973_),
    .A2(_10869_),
    .B1(_10976_),
    .B2(_10987_),
    .X(_10988_));
 sky130_fd_sc_hd__inv_2 _15062_ (.A(_10988_),
    .Y(_00925_));
 sky130_fd_sc_hd__nor2_1 _15063_ (.A(_10872_),
    .B(_10976_),
    .Y(_10989_));
 sky130_fd_sc_hd__a31o_1 _15064_ (.A1(_10937_),
    .A2(net437),
    .A3(_10979_),
    .B1(_10989_),
    .X(_00926_));
 sky130_fd_sc_hd__nand2_1 _15065_ (.A(_10884_),
    .B(net3718),
    .Y(_10990_));
 sky130_fd_sc_hd__a22o_1 _15066_ (.A1(_10973_),
    .A2(_10591_),
    .B1(_10975_),
    .B2(_10990_),
    .X(_10991_));
 sky130_fd_sc_hd__inv_2 _15067_ (.A(_10991_),
    .Y(_00927_));
 sky130_fd_sc_hd__nor2_1 _15068_ (.A(_10760_),
    .B(_10976_),
    .Y(_10992_));
 sky130_fd_sc_hd__a31o_1 _15069_ (.A1(_10937_),
    .A2(net1111),
    .A3(_10979_),
    .B1(_10992_),
    .X(_00912_));
 sky130_fd_sc_hd__nand2_1 _15070_ (.A(_10884_),
    .B(net3887),
    .Y(_10993_));
 sky130_fd_sc_hd__a22o_1 _15071_ (.A1(_10973_),
    .A2(_10122_),
    .B1(_10975_),
    .B2(_10993_),
    .X(_10994_));
 sky130_fd_sc_hd__inv_2 _15072_ (.A(_10994_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand2_1 _15073_ (.A(_10884_),
    .B(net4196),
    .Y(_10995_));
 sky130_fd_sc_hd__a22o_1 _15074_ (.A1(_10973_),
    .A2(_10195_),
    .B1(_10975_),
    .B2(_10995_),
    .X(_10996_));
 sky130_fd_sc_hd__inv_2 _15075_ (.A(_10996_),
    .Y(_00914_));
 sky130_fd_sc_hd__nor2_1 _15076_ (.A(_10657_),
    .B(_10976_),
    .Y(_10997_));
 sky130_fd_sc_hd__a31o_1 _15077_ (.A1(_10937_),
    .A2(net1335),
    .A3(_10979_),
    .B1(_10997_),
    .X(_00915_));
 sky130_fd_sc_hd__nor2_1 _15078_ (.A(_10767_),
    .B(_10976_),
    .Y(_10998_));
 sky130_fd_sc_hd__a31o_1 _15079_ (.A1(_10937_),
    .A2(net1949),
    .A3(_10979_),
    .B1(_10998_),
    .X(_00916_));
 sky130_fd_sc_hd__nor2_1 _15080_ (.A(_10602_),
    .B(_10976_),
    .Y(_10999_));
 sky130_fd_sc_hd__a31o_1 _15081_ (.A1(_10937_),
    .A2(net2341),
    .A3(_10979_),
    .B1(_10999_),
    .X(_00917_));
 sky130_fd_sc_hd__and3_1 _15082_ (.A(_10971_),
    .B(_09341_),
    .C(_10908_),
    .X(_11000_));
 sky130_fd_sc_hd__a31o_1 _15083_ (.A1(_10979_),
    .A2(_10903_),
    .A3(net2380),
    .B1(_11000_),
    .X(_00918_));
 sky130_fd_sc_hd__nor2_1 _15084_ (.A(_10663_),
    .B(_10976_),
    .Y(_11001_));
 sky130_fd_sc_hd__a31o_1 _15085_ (.A1(_10937_),
    .A2(net2489),
    .A3(_10979_),
    .B1(_11001_),
    .X(_00919_));
 sky130_fd_sc_hd__clkbuf_16 _15086_ (.A(_09245_),
    .X(_11002_));
 sky130_fd_sc_hd__nor2_1 _15087_ (.A(_11002_),
    .B(_10976_),
    .Y(_11003_));
 sky130_fd_sc_hd__a31o_1 _15088_ (.A1(_10937_),
    .A2(net1775),
    .A3(_10979_),
    .B1(_11003_),
    .X(_00904_));
 sky130_fd_sc_hd__and3_1 _15089_ (.A(_10971_),
    .B(_10667_),
    .C(_10908_),
    .X(_11004_));
 sky130_fd_sc_hd__a31o_1 _15090_ (.A1(_10979_),
    .A2(_10903_),
    .A3(net2375),
    .B1(_11004_),
    .X(_00905_));
 sky130_fd_sc_hd__nor2_1 _15091_ (.A(_10669_),
    .B(_10976_),
    .Y(_11005_));
 sky130_fd_sc_hd__a31o_1 _15092_ (.A1(_10937_),
    .A2(net2296),
    .A3(_10976_),
    .B1(_11005_),
    .X(_00906_));
 sky130_fd_sc_hd__buf_4 _15093_ (.A(_10349_),
    .X(_11006_));
 sky130_fd_sc_hd__nand2_1 _15094_ (.A(_11006_),
    .B(net3741),
    .Y(_11007_));
 sky130_fd_sc_hd__a22o_1 _15095_ (.A1(_10973_),
    .A2(_09256_),
    .B1(_10975_),
    .B2(_11007_),
    .X(_11008_));
 sky130_fd_sc_hd__inv_2 _15096_ (.A(_11008_),
    .Y(_00907_));
 sky130_fd_sc_hd__clkbuf_8 _15097_ (.A(_10864_),
    .X(_11009_));
 sky130_fd_sc_hd__buf_12 _15098_ (.A(_09259_),
    .X(_11010_));
 sky130_fd_sc_hd__nor2_1 _15099_ (.A(_11010_),
    .B(_10976_),
    .Y(_11011_));
 sky130_fd_sc_hd__a31o_1 _15100_ (.A1(_11009_),
    .A2(net1035),
    .A3(_10976_),
    .B1(_11011_),
    .X(_00908_));
 sky130_fd_sc_hd__nand2_1 _15101_ (.A(_11006_),
    .B(net3697),
    .Y(_11012_));
 sky130_fd_sc_hd__a22o_1 _15102_ (.A1(_10973_),
    .A2(_10149_),
    .B1(_10975_),
    .B2(_11012_),
    .X(_11013_));
 sky130_fd_sc_hd__inv_2 _15103_ (.A(_11013_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand2_1 _15104_ (.A(_11006_),
    .B(net3464),
    .Y(_11014_));
 sky130_fd_sc_hd__a22o_1 _15105_ (.A1(_10973_),
    .A2(_09425_),
    .B1(_10975_),
    .B2(_11014_),
    .X(_11015_));
 sky130_fd_sc_hd__inv_2 _15106_ (.A(_11015_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand2_1 _15107_ (.A(_11006_),
    .B(net3755),
    .Y(_11016_));
 sky130_fd_sc_hd__a22o_1 _15108_ (.A1(_10973_),
    .A2(_10154_),
    .B1(_10975_),
    .B2(_11016_),
    .X(_11017_));
 sky130_fd_sc_hd__inv_2 _15109_ (.A(_11017_),
    .Y(_00911_));
 sky130_fd_sc_hd__and3_1 _15110_ (.A(_10971_),
    .B(_10679_),
    .C(_10908_),
    .X(_11018_));
 sky130_fd_sc_hd__a31o_1 _15111_ (.A1(_10979_),
    .A2(_10903_),
    .A3(net1285),
    .B1(_11018_),
    .X(_00896_));
 sky130_fd_sc_hd__nand2_1 _15112_ (.A(_11006_),
    .B(net3874),
    .Y(_11019_));
 sky130_fd_sc_hd__a22o_1 _15113_ (.A1(_10973_),
    .A2(_09366_),
    .B1(_10975_),
    .B2(_11019_),
    .X(_11020_));
 sky130_fd_sc_hd__inv_2 _15114_ (.A(_11020_),
    .Y(_00897_));
 sky130_fd_sc_hd__and3_1 _15115_ (.A(_10971_),
    .B(_10728_),
    .C(_10908_),
    .X(_11021_));
 sky130_fd_sc_hd__a31o_1 _15116_ (.A1(_10979_),
    .A2(_10903_),
    .A3(net1778),
    .B1(_11021_),
    .X(_00898_));
 sky130_fd_sc_hd__nand2_1 _15117_ (.A(_11006_),
    .B(net3687),
    .Y(_11022_));
 sky130_fd_sc_hd__a22o_1 _15118_ (.A1(_10973_),
    .A2(_10164_),
    .B1(_10975_),
    .B2(_11022_),
    .X(_11023_));
 sky130_fd_sc_hd__inv_2 _15119_ (.A(_11023_),
    .Y(_00899_));
 sky130_fd_sc_hd__nand2_1 _15120_ (.A(_11006_),
    .B(net3036),
    .Y(_11024_));
 sky130_fd_sc_hd__a22o_1 _15121_ (.A1(_10973_),
    .A2(net139),
    .B1(_10975_),
    .B2(_11024_),
    .X(_11025_));
 sky130_fd_sc_hd__inv_2 _15122_ (.A(_11025_),
    .Y(_00900_));
 sky130_fd_sc_hd__and3_1 _15123_ (.A(_10971_),
    .B(_09730_),
    .C(_10908_),
    .X(_11026_));
 sky130_fd_sc_hd__a31o_1 _15124_ (.A1(_10979_),
    .A2(_10903_),
    .A3(net2646),
    .B1(_11026_),
    .X(_00901_));
 sky130_fd_sc_hd__nand2_1 _15125_ (.A(_10721_),
    .B(net3760),
    .Y(_11027_));
 sky130_fd_sc_hd__o2bb2a_1 _15126_ (.A1_N(_11027_),
    .A2_N(_10979_),
    .B1(_10289_),
    .B2(_10972_),
    .X(_00902_));
 sky130_fd_sc_hd__nand2_1 _15127_ (.A(_10721_),
    .B(net3770),
    .Y(_11028_));
 sky130_fd_sc_hd__o2bb2a_1 _15128_ (.A1_N(_11028_),
    .A2_N(_10979_),
    .B1(_09442_),
    .B2(_10972_),
    .X(_00903_));
 sky130_fd_sc_hd__nor2_2 _15129_ (.A(_10912_),
    .B(_10356_),
    .Y(_11029_));
 sky130_fd_sc_hd__inv_2 _15130_ (.A(_11029_),
    .Y(_11030_));
 sky130_fd_sc_hd__nor2_4 _15131_ (.A(_08797_),
    .B(_11030_),
    .Y(_11031_));
 sky130_fd_sc_hd__nor2_1 _15132_ (.A(_09625_),
    .B(_11030_),
    .Y(_11032_));
 sky130_fd_sc_hd__inv_2 _15133_ (.A(_11032_),
    .Y(_11033_));
 sky130_fd_sc_hd__buf_4 _15134_ (.A(_11033_),
    .X(_11034_));
 sky130_fd_sc_hd__nand2_1 _15135_ (.A(_11006_),
    .B(net3834),
    .Y(_11035_));
 sky130_fd_sc_hd__a22o_1 _15136_ (.A1(_11031_),
    .A2(_10239_),
    .B1(_11034_),
    .B2(_11035_),
    .X(_11036_));
 sky130_fd_sc_hd__inv_2 _15137_ (.A(_11036_),
    .Y(_00872_));
 sky130_fd_sc_hd__buf_4 _15138_ (.A(_11033_),
    .X(_11037_));
 sky130_fd_sc_hd__nor2_1 _15139_ (.A(_10746_),
    .B(_11034_),
    .Y(_11038_));
 sky130_fd_sc_hd__a31o_1 _15140_ (.A1(_11009_),
    .A2(net1836),
    .A3(_11037_),
    .B1(_11038_),
    .X(_00873_));
 sky130_fd_sc_hd__nor2_1 _15141_ (.A(_10698_),
    .B(_11034_),
    .Y(_11039_));
 sky130_fd_sc_hd__a31o_1 _15142_ (.A1(_11009_),
    .A2(net1663),
    .A3(_11037_),
    .B1(_11039_),
    .X(_00874_));
 sky130_fd_sc_hd__buf_12 _15143_ (.A(net69),
    .X(_11040_));
 sky130_fd_sc_hd__and3_1 _15144_ (.A(_11029_),
    .B(_11040_),
    .C(_10908_),
    .X(_11041_));
 sky130_fd_sc_hd__a31o_1 _15145_ (.A1(_11037_),
    .A2(_10903_),
    .A3(net2663),
    .B1(_11041_),
    .X(_00875_));
 sky130_fd_sc_hd__nand2_1 _15146_ (.A(_11006_),
    .B(net3469),
    .Y(_11042_));
 sky130_fd_sc_hd__a22o_1 _15147_ (.A1(_11031_),
    .A2(_09201_),
    .B1(_11034_),
    .B2(_11042_),
    .X(_11043_));
 sky130_fd_sc_hd__inv_2 _15148_ (.A(_11043_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand2_1 _15149_ (.A(_11006_),
    .B(net3683),
    .Y(_11044_));
 sky130_fd_sc_hd__a22o_1 _15150_ (.A1(_11031_),
    .A2(_10869_),
    .B1(_11034_),
    .B2(_11044_),
    .X(_11045_));
 sky130_fd_sc_hd__inv_2 _15151_ (.A(_11045_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_1 _15152_ (.A(_11006_),
    .B(net3952),
    .Y(_11046_));
 sky130_fd_sc_hd__a22o_1 _15153_ (.A1(_11031_),
    .A2(_09398_),
    .B1(_11034_),
    .B2(_11046_),
    .X(_11047_));
 sky130_fd_sc_hd__inv_2 _15154_ (.A(_11047_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand2_1 _15155_ (.A(_11006_),
    .B(net3843),
    .Y(_11048_));
 sky130_fd_sc_hd__a22o_1 _15156_ (.A1(_11031_),
    .A2(_10591_),
    .B1(_11034_),
    .B2(_11048_),
    .X(_11049_));
 sky130_fd_sc_hd__inv_2 _15157_ (.A(_11049_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _15158_ (.A(_11006_),
    .B(net2831),
    .Y(_11050_));
 sky130_fd_sc_hd__a22o_1 _15159_ (.A1(_11031_),
    .A2(_09531_),
    .B1(_11034_),
    .B2(_11050_),
    .X(_11051_));
 sky130_fd_sc_hd__inv_2 _15160_ (.A(_11051_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2_1 _15161_ (.A(_11006_),
    .B(net3325),
    .Y(_11052_));
 sky130_fd_sc_hd__a22o_1 _15162_ (.A1(_11031_),
    .A2(_10122_),
    .B1(_11033_),
    .B2(_11052_),
    .X(_11053_));
 sky130_fd_sc_hd__inv_2 _15163_ (.A(_11053_),
    .Y(_00865_));
 sky130_fd_sc_hd__nand2_1 _15164_ (.A(_11006_),
    .B(net3606),
    .Y(_11054_));
 sky130_fd_sc_hd__a22o_1 _15165_ (.A1(_11031_),
    .A2(_10195_),
    .B1(_11033_),
    .B2(_11054_),
    .X(_11055_));
 sky130_fd_sc_hd__inv_2 _15166_ (.A(_11055_),
    .Y(_00866_));
 sky130_fd_sc_hd__nor2_1 _15167_ (.A(_10657_),
    .B(_11034_),
    .Y(_11056_));
 sky130_fd_sc_hd__a31o_1 _15168_ (.A1(_11009_),
    .A2(net1243),
    .A3(_11037_),
    .B1(_11056_),
    .X(_00867_));
 sky130_fd_sc_hd__nor2_1 _15169_ (.A(_10767_),
    .B(_11034_),
    .Y(_11057_));
 sky130_fd_sc_hd__a31o_1 _15170_ (.A1(_11009_),
    .A2(net871),
    .A3(_11037_),
    .B1(_11057_),
    .X(_00868_));
 sky130_fd_sc_hd__nor2_1 _15171_ (.A(_10602_),
    .B(_11034_),
    .Y(_11058_));
 sky130_fd_sc_hd__a31o_1 _15172_ (.A1(_11009_),
    .A2(net1759),
    .A3(_11037_),
    .B1(_11058_),
    .X(_00869_));
 sky130_fd_sc_hd__and3_1 _15173_ (.A(_11029_),
    .B(_09341_),
    .C(_10908_),
    .X(_11059_));
 sky130_fd_sc_hd__a31o_1 _15174_ (.A1(_11037_),
    .A2(_10903_),
    .A3(net2241),
    .B1(_11059_),
    .X(_00870_));
 sky130_fd_sc_hd__nor2_1 _15175_ (.A(_10663_),
    .B(_11034_),
    .Y(_11060_));
 sky130_fd_sc_hd__a31o_1 _15176_ (.A1(_11009_),
    .A2(net2396),
    .A3(_11037_),
    .B1(_11060_),
    .X(_00871_));
 sky130_fd_sc_hd__nor2_1 _15177_ (.A(_11002_),
    .B(_11034_),
    .Y(_11061_));
 sky130_fd_sc_hd__a31o_1 _15178_ (.A1(_11009_),
    .A2(net431),
    .A3(_11034_),
    .B1(_11061_),
    .X(_00856_));
 sky130_fd_sc_hd__and3_1 _15179_ (.A(_11029_),
    .B(_10667_),
    .C(_10908_),
    .X(_11062_));
 sky130_fd_sc_hd__a31o_1 _15180_ (.A1(_11037_),
    .A2(_10903_),
    .A3(net2459),
    .B1(_11062_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_1 _15181_ (.A(_11006_),
    .B(net3005),
    .Y(_11063_));
 sky130_fd_sc_hd__a22o_1 _15182_ (.A1(_11031_),
    .A2(_09348_),
    .B1(_11033_),
    .B2(_11063_),
    .X(_11064_));
 sky130_fd_sc_hd__inv_2 _15183_ (.A(_11064_),
    .Y(_00858_));
 sky130_fd_sc_hd__and3_1 _15184_ (.A(_11029_),
    .B(_10500_),
    .C(_10908_),
    .X(_11065_));
 sky130_fd_sc_hd__a31o_1 _15185_ (.A1(_11037_),
    .A2(_10903_),
    .A3(net2258),
    .B1(_11065_),
    .X(_00859_));
 sky130_fd_sc_hd__nor2_1 _15186_ (.A(_11010_),
    .B(_11034_),
    .Y(_11066_));
 sky130_fd_sc_hd__a31o_1 _15187_ (.A1(_11009_),
    .A2(net1844),
    .A3(_11034_),
    .B1(_11066_),
    .X(_00860_));
 sky130_fd_sc_hd__buf_4 _15188_ (.A(_10349_),
    .X(_11067_));
 sky130_fd_sc_hd__nand2_1 _15189_ (.A(_11067_),
    .B(net3318),
    .Y(_11068_));
 sky130_fd_sc_hd__a22o_1 _15190_ (.A1(_11031_),
    .A2(_10149_),
    .B1(_11033_),
    .B2(_11068_),
    .X(_11069_));
 sky130_fd_sc_hd__inv_2 _15191_ (.A(_11069_),
    .Y(_00861_));
 sky130_fd_sc_hd__nand2_1 _15192_ (.A(_11067_),
    .B(net3417),
    .Y(_11070_));
 sky130_fd_sc_hd__a22o_1 _15193_ (.A1(_11031_),
    .A2(_09425_),
    .B1(_11033_),
    .B2(_11070_),
    .X(_11071_));
 sky130_fd_sc_hd__inv_2 _15194_ (.A(_11071_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _15195_ (.A(_11067_),
    .B(net3720),
    .Y(_11072_));
 sky130_fd_sc_hd__a22o_1 _15196_ (.A1(_11031_),
    .A2(_10154_),
    .B1(_11033_),
    .B2(_11072_),
    .X(_11073_));
 sky130_fd_sc_hd__inv_2 _15197_ (.A(_11073_),
    .Y(_00863_));
 sky130_fd_sc_hd__buf_4 _15198_ (.A(_09359_),
    .X(_11074_));
 sky130_fd_sc_hd__and3_1 _15199_ (.A(_11029_),
    .B(_10679_),
    .C(_11074_),
    .X(_11075_));
 sky130_fd_sc_hd__a31o_1 _15200_ (.A1(_11037_),
    .A2(_10903_),
    .A3(net1471),
    .B1(_11075_),
    .X(_00848_));
 sky130_fd_sc_hd__nand2_1 _15201_ (.A(_11067_),
    .B(net3465),
    .Y(_11076_));
 sky130_fd_sc_hd__a22o_1 _15202_ (.A1(_11031_),
    .A2(_09366_),
    .B1(_11033_),
    .B2(_11076_),
    .X(_11077_));
 sky130_fd_sc_hd__inv_2 _15203_ (.A(_11077_),
    .Y(_00849_));
 sky130_fd_sc_hd__and3_1 _15204_ (.A(_11029_),
    .B(_10728_),
    .C(_11074_),
    .X(_11078_));
 sky130_fd_sc_hd__a31o_1 _15205_ (.A1(_11037_),
    .A2(_10903_),
    .A3(net2586),
    .B1(_11078_),
    .X(_00850_));
 sky130_fd_sc_hd__nand2_1 _15206_ (.A(_11067_),
    .B(net3753),
    .Y(_11079_));
 sky130_fd_sc_hd__a22o_1 _15207_ (.A1(_11031_),
    .A2(_10164_),
    .B1(_11033_),
    .B2(_11079_),
    .X(_11080_));
 sky130_fd_sc_hd__inv_2 _15208_ (.A(_11080_),
    .Y(_00851_));
 sky130_fd_sc_hd__and3_1 _15209_ (.A(_11029_),
    .B(_10848_),
    .C(_11074_),
    .X(_11081_));
 sky130_fd_sc_hd__a31o_1 _15210_ (.A1(_11037_),
    .A2(_10903_),
    .A3(net1539),
    .B1(_11081_),
    .X(_00852_));
 sky130_fd_sc_hd__clkbuf_8 _15211_ (.A(_10645_),
    .X(_11082_));
 sky130_fd_sc_hd__and3_1 _15212_ (.A(_11029_),
    .B(_09730_),
    .C(_11074_),
    .X(_11083_));
 sky130_fd_sc_hd__a31o_1 _15213_ (.A1(_11037_),
    .A2(_11082_),
    .A3(net2707),
    .B1(_11083_),
    .X(_00853_));
 sky130_fd_sc_hd__nand2_1 _15214_ (.A(_10721_),
    .B(net3551),
    .Y(_11084_));
 sky130_fd_sc_hd__o2bb2a_1 _15215_ (.A1_N(_11084_),
    .A2_N(_11037_),
    .B1(_10289_),
    .B2(_11030_),
    .X(_00854_));
 sky130_fd_sc_hd__nand2_1 _15216_ (.A(_10721_),
    .B(net3694),
    .Y(_11085_));
 sky130_fd_sc_hd__o2bb2a_1 _15217_ (.A1_N(_11085_),
    .A2_N(_11037_),
    .B1(_09442_),
    .B2(_11030_),
    .X(_00855_));
 sky130_fd_sc_hd__nor2_1 _15218_ (.A(_10912_),
    .B(_10411_),
    .Y(_11086_));
 sky130_fd_sc_hd__inv_2 _15219_ (.A(_11086_),
    .Y(_11087_));
 sky130_fd_sc_hd__nor2_4 _15220_ (.A(_08794_),
    .B(_11087_),
    .Y(_11088_));
 sky130_fd_sc_hd__buf_4 _15221_ (.A(_11088_),
    .X(_11089_));
 sky130_fd_sc_hd__nor2_1 _15222_ (.A(_09625_),
    .B(_11087_),
    .Y(_11090_));
 sky130_fd_sc_hd__inv_2 _15223_ (.A(_11090_),
    .Y(_11091_));
 sky130_fd_sc_hd__buf_4 _15224_ (.A(_11091_),
    .X(_11092_));
 sky130_fd_sc_hd__nand2_1 _15225_ (.A(_11067_),
    .B(net3506),
    .Y(_11093_));
 sky130_fd_sc_hd__a22o_1 _15226_ (.A1(_11089_),
    .A2(_10239_),
    .B1(_11092_),
    .B2(_11093_),
    .X(_11094_));
 sky130_fd_sc_hd__inv_2 _15227_ (.A(_11094_),
    .Y(_00840_));
 sky130_fd_sc_hd__nand2_1 _15228_ (.A(_11067_),
    .B(net3383),
    .Y(_11095_));
 sky130_fd_sc_hd__a22o_1 _15229_ (.A1(_11089_),
    .A2(_09315_),
    .B1(_11092_),
    .B2(_11095_),
    .X(_11096_));
 sky130_fd_sc_hd__inv_2 _15230_ (.A(_11096_),
    .Y(_00841_));
 sky130_fd_sc_hd__nand2_1 _15231_ (.A(_11067_),
    .B(net3772),
    .Y(_11097_));
 sky130_fd_sc_hd__a22o_1 _15232_ (.A1(_11089_),
    .A2(_09460_),
    .B1(_11092_),
    .B2(_11097_),
    .X(_11098_));
 sky130_fd_sc_hd__inv_2 _15233_ (.A(_11098_),
    .Y(_00842_));
 sky130_fd_sc_hd__nand2_1 _15234_ (.A(_11067_),
    .B(net3593),
    .Y(_11099_));
 sky130_fd_sc_hd__a22o_1 _15235_ (.A1(_11089_),
    .A2(_10983_),
    .B1(_11092_),
    .B2(_11099_),
    .X(_11100_));
 sky130_fd_sc_hd__inv_2 _15236_ (.A(_11100_),
    .Y(_00843_));
 sky130_fd_sc_hd__nand2_1 _15237_ (.A(_11067_),
    .B(net3604),
    .Y(_11101_));
 sky130_fd_sc_hd__a22o_1 _15238_ (.A1(_11089_),
    .A2(_09201_),
    .B1(_11092_),
    .B2(_11101_),
    .X(_11102_));
 sky130_fd_sc_hd__inv_2 _15239_ (.A(_11102_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _15240_ (.A(_11067_),
    .B(net3523),
    .Y(_11103_));
 sky130_fd_sc_hd__a22o_1 _15241_ (.A1(_11089_),
    .A2(_10869_),
    .B1(_11092_),
    .B2(_11103_),
    .X(_11104_));
 sky130_fd_sc_hd__inv_2 _15242_ (.A(_11104_),
    .Y(_00845_));
 sky130_fd_sc_hd__buf_12 _15243_ (.A(_09397_),
    .X(_11105_));
 sky130_fd_sc_hd__nand2_1 _15244_ (.A(_11067_),
    .B(net2960),
    .Y(_11106_));
 sky130_fd_sc_hd__a22o_1 _15245_ (.A1(_11089_),
    .A2(_11105_),
    .B1(_11092_),
    .B2(_11106_),
    .X(_11107_));
 sky130_fd_sc_hd__inv_2 _15246_ (.A(_11107_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _15247_ (.A(_11067_),
    .B(net3828),
    .Y(_11108_));
 sky130_fd_sc_hd__a22o_1 _15248_ (.A1(_11089_),
    .A2(_10591_),
    .B1(_11092_),
    .B2(_11108_),
    .X(_11109_));
 sky130_fd_sc_hd__inv_2 _15249_ (.A(_11109_),
    .Y(_00847_));
 sky130_fd_sc_hd__nand2_1 _15250_ (.A(_11067_),
    .B(net2858),
    .Y(_11110_));
 sky130_fd_sc_hd__a22o_1 _15251_ (.A1(_11089_),
    .A2(_09530_),
    .B1(_11092_),
    .B2(_11110_),
    .X(_11111_));
 sky130_fd_sc_hd__inv_2 _15252_ (.A(_11111_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand2_1 _15253_ (.A(_11067_),
    .B(net3602),
    .Y(_11112_));
 sky130_fd_sc_hd__a22o_1 _15254_ (.A1(_11089_),
    .A2(_10122_),
    .B1(_11092_),
    .B2(_11112_),
    .X(_11113_));
 sky130_fd_sc_hd__inv_2 _15255_ (.A(_11113_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand2_1 _15256_ (.A(_11067_),
    .B(net3572),
    .Y(_11114_));
 sky130_fd_sc_hd__a22o_1 _15257_ (.A1(_11089_),
    .A2(_10195_),
    .B1(_11092_),
    .B2(_11114_),
    .X(_11115_));
 sky130_fd_sc_hd__inv_2 _15258_ (.A(_11115_),
    .Y(_00834_));
 sky130_fd_sc_hd__buf_4 _15259_ (.A(_10349_),
    .X(_11116_));
 sky130_fd_sc_hd__nand2_1 _15260_ (.A(_11116_),
    .B(net2808),
    .Y(_11117_));
 sky130_fd_sc_hd__a22o_1 _15261_ (.A1(_11089_),
    .A2(_09589_),
    .B1(_11092_),
    .B2(_11117_),
    .X(_11118_));
 sky130_fd_sc_hd__inv_2 _15262_ (.A(_11118_),
    .Y(_00835_));
 sky130_fd_sc_hd__nand2_1 _15263_ (.A(_11116_),
    .B(net2847),
    .Y(_11119_));
 sky130_fd_sc_hd__a22o_1 _15264_ (.A1(_11089_),
    .A2(_09593_),
    .B1(_11092_),
    .B2(_11119_),
    .X(_11120_));
 sky130_fd_sc_hd__inv_2 _15265_ (.A(_11120_),
    .Y(_00836_));
 sky130_fd_sc_hd__nand2_1 _15266_ (.A(_11116_),
    .B(net2855),
    .Y(_11121_));
 sky130_fd_sc_hd__a22o_1 _15267_ (.A1(_11089_),
    .A2(_09338_),
    .B1(_11092_),
    .B2(_11121_),
    .X(_11122_));
 sky130_fd_sc_hd__inv_2 _15268_ (.A(_11122_),
    .Y(_00837_));
 sky130_fd_sc_hd__buf_4 _15269_ (.A(_11091_),
    .X(_11123_));
 sky130_fd_sc_hd__nand2_1 _15270_ (.A(_11116_),
    .B(net2822),
    .Y(_11124_));
 sky130_fd_sc_hd__a22o_1 _15271_ (.A1(_11089_),
    .A2(_10202_),
    .B1(_11123_),
    .B2(_11124_),
    .X(_11125_));
 sky130_fd_sc_hd__inv_2 _15272_ (.A(_11125_),
    .Y(_00838_));
 sky130_fd_sc_hd__nand2_1 _15273_ (.A(_11116_),
    .B(net2795),
    .Y(_11126_));
 sky130_fd_sc_hd__a22o_1 _15274_ (.A1(_11089_),
    .A2(_09768_),
    .B1(_11123_),
    .B2(_11126_),
    .X(_11127_));
 sky130_fd_sc_hd__inv_2 _15275_ (.A(_11127_),
    .Y(_00839_));
 sky130_fd_sc_hd__nand2_1 _15276_ (.A(_11116_),
    .B(net2854),
    .Y(_11128_));
 sky130_fd_sc_hd__a22o_1 _15277_ (.A1(_11088_),
    .A2(_09414_),
    .B1(_11123_),
    .B2(_11128_),
    .X(_11129_));
 sky130_fd_sc_hd__inv_2 _15278_ (.A(_11129_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_1 _15279_ (.A(_11116_),
    .B(net2889),
    .Y(_11130_));
 sky130_fd_sc_hd__a22o_1 _15280_ (.A1(_11088_),
    .A2(_09249_),
    .B1(_11123_),
    .B2(_11130_),
    .X(_11131_));
 sky130_fd_sc_hd__inv_2 _15281_ (.A(_11131_),
    .Y(_00825_));
 sky130_fd_sc_hd__nand2_1 _15282_ (.A(_11116_),
    .B(net3321),
    .Y(_11132_));
 sky130_fd_sc_hd__a22o_1 _15283_ (.A1(_11088_),
    .A2(_09348_),
    .B1(_11123_),
    .B2(_11132_),
    .X(_11133_));
 sky130_fd_sc_hd__inv_2 _15284_ (.A(_11133_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _15285_ (.A(_11116_),
    .B(net3273),
    .Y(_11134_));
 sky130_fd_sc_hd__a22o_1 _15286_ (.A1(_11088_),
    .A2(_09256_),
    .B1(_11123_),
    .B2(_11134_),
    .X(_11135_));
 sky130_fd_sc_hd__inv_2 _15287_ (.A(_11135_),
    .Y(_00827_));
 sky130_fd_sc_hd__buf_12 _15288_ (.A(_09353_),
    .X(_11136_));
 sky130_fd_sc_hd__nand2_1 _15289_ (.A(_11116_),
    .B(net2863),
    .Y(_11137_));
 sky130_fd_sc_hd__a22o_1 _15290_ (.A1(_11088_),
    .A2(_11136_),
    .B1(_11123_),
    .B2(_11137_),
    .X(_11138_));
 sky130_fd_sc_hd__inv_2 _15291_ (.A(_11138_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_1 _15292_ (.A(_11116_),
    .B(net3135),
    .Y(_11139_));
 sky130_fd_sc_hd__a22o_1 _15293_ (.A1(_11088_),
    .A2(_10149_),
    .B1(_11123_),
    .B2(_11139_),
    .X(_11140_));
 sky130_fd_sc_hd__inv_2 _15294_ (.A(_11140_),
    .Y(_00829_));
 sky130_fd_sc_hd__nand2_1 _15295_ (.A(_11116_),
    .B(net2836),
    .Y(_11141_));
 sky130_fd_sc_hd__a22o_1 _15296_ (.A1(_11088_),
    .A2(_09425_),
    .B1(_11123_),
    .B2(_11141_),
    .X(_11142_));
 sky130_fd_sc_hd__inv_2 _15297_ (.A(_11142_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_1 _15298_ (.A(_11116_),
    .B(net2986),
    .Y(_11143_));
 sky130_fd_sc_hd__a22o_1 _15299_ (.A1(_11088_),
    .A2(_10154_),
    .B1(_11123_),
    .B2(_11143_),
    .X(_11144_));
 sky130_fd_sc_hd__inv_2 _15300_ (.A(_11144_),
    .Y(_00831_));
 sky130_fd_sc_hd__nand2_1 _15301_ (.A(_11116_),
    .B(net2815),
    .Y(_11145_));
 sky130_fd_sc_hd__a22o_1 _15302_ (.A1(_11088_),
    .A2(_09495_),
    .B1(_11123_),
    .B2(_11145_),
    .X(_11146_));
 sky130_fd_sc_hd__inv_2 _15303_ (.A(_11146_),
    .Y(_00816_));
 sky130_fd_sc_hd__nand2_1 _15304_ (.A(_11116_),
    .B(net2830),
    .Y(_11147_));
 sky130_fd_sc_hd__a22o_1 _15305_ (.A1(_11088_),
    .A2(_09366_),
    .B1(_11123_),
    .B2(_11147_),
    .X(_11148_));
 sky130_fd_sc_hd__inv_2 _15306_ (.A(_11148_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_1 _15307_ (.A(_11116_),
    .B(net2806),
    .Y(_11149_));
 sky130_fd_sc_hd__a22o_1 _15308_ (.A1(_11088_),
    .A2(_10624_),
    .B1(_11123_),
    .B2(_11149_),
    .X(_11150_));
 sky130_fd_sc_hd__inv_2 _15309_ (.A(_11150_),
    .Y(_00818_));
 sky130_fd_sc_hd__buf_4 _15310_ (.A(_08775_),
    .X(_11151_));
 sky130_fd_sc_hd__buf_6 _15311_ (.A(_11151_),
    .X(_11152_));
 sky130_fd_sc_hd__nand2_1 _15312_ (.A(_11152_),
    .B(net2837),
    .Y(_11153_));
 sky130_fd_sc_hd__a22o_1 _15313_ (.A1(_11088_),
    .A2(_10164_),
    .B1(_11123_),
    .B2(_11153_),
    .X(_11154_));
 sky130_fd_sc_hd__inv_2 _15314_ (.A(_11154_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _15315_ (.A(_11152_),
    .B(net2805),
    .Y(_11155_));
 sky130_fd_sc_hd__a22o_1 _15316_ (.A1(_11088_),
    .A2(net139),
    .B1(_11123_),
    .B2(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__inv_2 _15317_ (.A(_11156_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand2_1 _15318_ (.A(_11152_),
    .B(net2777),
    .Y(_11157_));
 sky130_fd_sc_hd__a22o_1 _15319_ (.A1(_11088_),
    .A2(_09504_),
    .B1(_11123_),
    .B2(_11157_),
    .X(_11158_));
 sky130_fd_sc_hd__inv_2 _15320_ (.A(_11158_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand2_1 _15321_ (.A(_10721_),
    .B(net3235),
    .Y(_11159_));
 sky130_fd_sc_hd__o2bb2a_1 _15322_ (.A1_N(_11159_),
    .A2_N(_11092_),
    .B1(_10289_),
    .B2(_11087_),
    .X(_00822_));
 sky130_fd_sc_hd__nand2_1 _15323_ (.A(_10721_),
    .B(net3251),
    .Y(_11160_));
 sky130_fd_sc_hd__o2bb2a_1 _15324_ (.A1_N(_11160_),
    .A2_N(_11092_),
    .B1(_09442_),
    .B2(_11087_),
    .X(_00823_));
 sky130_fd_sc_hd__nor2_8 _15325_ (.A(net3899),
    .B(_08738_),
    .Y(_11161_));
 sky130_fd_sc_hd__nand2_4 _15326_ (.A(_11161_),
    .B(_09168_),
    .Y(_11162_));
 sky130_fd_sc_hd__nor2_1 _15327_ (.A(_11162_),
    .B(_10469_),
    .Y(_11163_));
 sky130_fd_sc_hd__nand2_4 _15328_ (.A(_11163_),
    .B(_09226_),
    .Y(_11164_));
 sky130_fd_sc_hd__buf_4 _15329_ (.A(_11164_),
    .X(_11165_));
 sky130_fd_sc_hd__buf_4 _15330_ (.A(_11164_),
    .X(_11166_));
 sky130_fd_sc_hd__nor2_1 _15331_ (.A(_09181_),
    .B(_11166_),
    .Y(_11167_));
 sky130_fd_sc_hd__a31o_1 _15332_ (.A1(_11009_),
    .A2(net2724),
    .A3(_11165_),
    .B1(_11167_),
    .X(_00808_));
 sky130_fd_sc_hd__nand2_1 _15333_ (.A(_10721_),
    .B(net4096),
    .Y(_11168_));
 sky130_fd_sc_hd__buf_4 _15334_ (.A(_11163_),
    .X(_11169_));
 sky130_fd_sc_hd__nand2_4 _15335_ (.A(_11169_),
    .B(_08778_),
    .Y(_11170_));
 sky130_fd_sc_hd__o2bb2a_1 _15336_ (.A1_N(_11168_),
    .A2_N(_11165_),
    .B1(_10475_),
    .B2(_11170_),
    .X(_00809_));
 sky130_fd_sc_hd__nor2_1 _15337_ (.A(_10698_),
    .B(_11166_),
    .Y(_11171_));
 sky130_fd_sc_hd__a31o_1 _15338_ (.A1(_11009_),
    .A2(net1379),
    .A3(_11165_),
    .B1(_11171_),
    .X(_00810_));
 sky130_fd_sc_hd__and3_1 _15339_ (.A(_11169_),
    .B(_11040_),
    .C(_11074_),
    .X(_11172_));
 sky130_fd_sc_hd__a31o_1 _15340_ (.A1(_11009_),
    .A2(net943),
    .A3(_11165_),
    .B1(_11172_),
    .X(_00811_));
 sky130_fd_sc_hd__and3_1 _15341_ (.A(_11169_),
    .B(_10587_),
    .C(_11074_),
    .X(_11173_));
 sky130_fd_sc_hd__a31o_1 _15342_ (.A1(_11009_),
    .A2(net2205),
    .A3(_11165_),
    .B1(_11173_),
    .X(_00812_));
 sky130_fd_sc_hd__clkbuf_8 _15343_ (.A(_09375_),
    .X(_11174_));
 sky130_fd_sc_hd__nand2_1 _15344_ (.A(_11174_),
    .B(net4097),
    .Y(_11175_));
 sky130_fd_sc_hd__o2bb2a_1 _15345_ (.A1_N(_11175_),
    .A2_N(_11165_),
    .B1(_10251_),
    .B2(_11170_),
    .X(_00813_));
 sky130_fd_sc_hd__nor2_1 _15346_ (.A(_10872_),
    .B(_11166_),
    .Y(_11176_));
 sky130_fd_sc_hd__a31o_1 _15347_ (.A1(_11009_),
    .A2(net2561),
    .A3(_11165_),
    .B1(_11176_),
    .X(_00814_));
 sky130_fd_sc_hd__and3_1 _15348_ (.A(_11169_),
    .B(_10874_),
    .C(_11074_),
    .X(_11177_));
 sky130_fd_sc_hd__a31o_1 _15349_ (.A1(_11009_),
    .A2(net2044),
    .A3(_11165_),
    .B1(_11177_),
    .X(_00815_));
 sky130_fd_sc_hd__nor2_1 _15350_ (.A(_10760_),
    .B(_11166_),
    .Y(_11178_));
 sky130_fd_sc_hd__a31o_1 _15351_ (.A1(_11009_),
    .A2(net2054),
    .A3(_11165_),
    .B1(_11178_),
    .X(_00800_));
 sky130_fd_sc_hd__nand2_1 _15352_ (.A(_11174_),
    .B(net4015),
    .Y(_11179_));
 sky130_fd_sc_hd__o2bb2a_1 _15353_ (.A1_N(_11179_),
    .A2_N(_11165_),
    .B1(_10257_),
    .B2(_11170_),
    .X(_00801_));
 sky130_fd_sc_hd__nand2_1 _15354_ (.A(_11174_),
    .B(net3625),
    .Y(_11180_));
 sky130_fd_sc_hd__o2bb2a_1 _15355_ (.A1_N(_11180_),
    .A2_N(_11165_),
    .B1(_10259_),
    .B2(_11170_),
    .X(_00802_));
 sky130_fd_sc_hd__a22o_1 _15356_ (.A1(_09302_),
    .A2(net3088),
    .B1(_11169_),
    .B2(_09227_),
    .X(_11181_));
 sky130_fd_sc_hd__o31a_1 _15357_ (.A1(_09193_),
    .A2(net60),
    .A3(_11170_),
    .B1(_11181_),
    .X(_00803_));
 sky130_fd_sc_hd__clkbuf_8 _15358_ (.A(_10864_),
    .X(_11182_));
 sky130_fd_sc_hd__nor2_1 _15359_ (.A(_10767_),
    .B(_11164_),
    .Y(_11183_));
 sky130_fd_sc_hd__a31o_1 _15360_ (.A1(_11182_),
    .A2(net1930),
    .A3(_11166_),
    .B1(_11183_),
    .X(_00804_));
 sky130_fd_sc_hd__nor2_1 _15361_ (.A(_10602_),
    .B(_11164_),
    .Y(_11184_));
 sky130_fd_sc_hd__a31o_1 _15362_ (.A1(_11182_),
    .A2(net2632),
    .A3(_11166_),
    .B1(_11184_),
    .X(_00805_));
 sky130_fd_sc_hd__and3_1 _15363_ (.A(_11169_),
    .B(_09341_),
    .C(_11074_),
    .X(_11185_));
 sky130_fd_sc_hd__a31o_1 _15364_ (.A1(_11182_),
    .A2(net2541),
    .A3(_11166_),
    .B1(_11185_),
    .X(_00806_));
 sky130_fd_sc_hd__a22o_1 _15365_ (.A1(_09302_),
    .A2(net2851),
    .B1(_11169_),
    .B2(_09227_),
    .X(_11186_));
 sky130_fd_sc_hd__o31a_1 _15366_ (.A1(_09193_),
    .A2(net65),
    .A3(_11170_),
    .B1(_11186_),
    .X(_00807_));
 sky130_fd_sc_hd__nor2_1 _15367_ (.A(_11002_),
    .B(_11164_),
    .Y(_11187_));
 sky130_fd_sc_hd__a31o_1 _15368_ (.A1(_11182_),
    .A2(net1255),
    .A3(_11166_),
    .B1(_11187_),
    .X(_00784_));
 sky130_fd_sc_hd__and3_1 _15369_ (.A(_11169_),
    .B(_10667_),
    .C(_11074_),
    .X(_11188_));
 sky130_fd_sc_hd__a31o_1 _15370_ (.A1(_11182_),
    .A2(net1149),
    .A3(_11166_),
    .B1(_11188_),
    .X(_00785_));
 sky130_fd_sc_hd__nor2_1 _15371_ (.A(_10669_),
    .B(_11164_),
    .Y(_11189_));
 sky130_fd_sc_hd__a31o_1 _15372_ (.A1(_11182_),
    .A2(net419),
    .A3(_11166_),
    .B1(_11189_),
    .X(_00786_));
 sky130_fd_sc_hd__and3_1 _15373_ (.A(_11169_),
    .B(_10500_),
    .C(_11074_),
    .X(_11190_));
 sky130_fd_sc_hd__a31o_1 _15374_ (.A1(_11182_),
    .A2(net2569),
    .A3(_11166_),
    .B1(_11190_),
    .X(_00787_));
 sky130_fd_sc_hd__nand2_1 _15375_ (.A(_11174_),
    .B(net4022),
    .Y(_11191_));
 sky130_fd_sc_hd__o2bb2a_1 _15376_ (.A1_N(_11191_),
    .A2_N(_11165_),
    .B1(_10503_),
    .B2(_11170_),
    .X(_00788_));
 sky130_fd_sc_hd__nand2_1 _15377_ (.A(_11174_),
    .B(net3583),
    .Y(_11192_));
 sky130_fd_sc_hd__o2bb2a_1 _15378_ (.A1_N(_11192_),
    .A2_N(_11165_),
    .B1(_10273_),
    .B2(_11170_),
    .X(_00789_));
 sky130_fd_sc_hd__and3_1 _15379_ (.A(_11169_),
    .B(_10617_),
    .C(_11074_),
    .X(_11193_));
 sky130_fd_sc_hd__a31o_1 _15380_ (.A1(_11182_),
    .A2(net845),
    .A3(_11166_),
    .B1(_11193_),
    .X(_00790_));
 sky130_fd_sc_hd__nand2_1 _15381_ (.A(_11174_),
    .B(net3396),
    .Y(_11194_));
 sky130_fd_sc_hd__o2bb2a_1 _15382_ (.A1_N(_11194_),
    .A2_N(_11165_),
    .B1(_10276_),
    .B2(_11170_),
    .X(_00791_));
 sky130_fd_sc_hd__and3_1 _15383_ (.A(_11169_),
    .B(_10679_),
    .C(_11074_),
    .X(_11195_));
 sky130_fd_sc_hd__a31o_1 _15384_ (.A1(_11182_),
    .A2(net1630),
    .A3(_11166_),
    .B1(_11195_),
    .X(_00776_));
 sky130_fd_sc_hd__nand2_1 _15385_ (.A(_11174_),
    .B(net3728),
    .Y(_11196_));
 sky130_fd_sc_hd__o2bb2a_1 _15386_ (.A1_N(_11196_),
    .A2_N(_11165_),
    .B1(_10727_),
    .B2(_11170_),
    .X(_00777_));
 sky130_fd_sc_hd__and3_1 _15387_ (.A(_11169_),
    .B(_10728_),
    .C(_11074_),
    .X(_11197_));
 sky130_fd_sc_hd__a31o_1 _15388_ (.A1(_11182_),
    .A2(net949),
    .A3(_11166_),
    .B1(_11197_),
    .X(_00778_));
 sky130_fd_sc_hd__nand2_1 _15389_ (.A(_11174_),
    .B(net4080),
    .Y(_11198_));
 sky130_fd_sc_hd__o2bb2a_1 _15390_ (.A1_N(_11198_),
    .A2_N(_11165_),
    .B1(_10285_),
    .B2(_11170_),
    .X(_00779_));
 sky130_fd_sc_hd__and3_1 _15391_ (.A(_11169_),
    .B(_10848_),
    .C(_11074_),
    .X(_11199_));
 sky130_fd_sc_hd__a31o_1 _15392_ (.A1(_11182_),
    .A2(net2574),
    .A3(_11166_),
    .B1(_11199_),
    .X(_00780_));
 sky130_fd_sc_hd__and3_1 _15393_ (.A(_11169_),
    .B(_09730_),
    .C(_11074_),
    .X(_11200_));
 sky130_fd_sc_hd__a31o_1 _15394_ (.A1(_11182_),
    .A2(net1591),
    .A3(_11166_),
    .B1(_11200_),
    .X(_00781_));
 sky130_fd_sc_hd__nand2_1 _15395_ (.A(_11152_),
    .B(net3170),
    .Y(_11201_));
 sky130_fd_sc_hd__a22o_1 _15396_ (.A1(_10348_),
    .A2(_11169_),
    .B1(_11164_),
    .B2(_11201_),
    .X(_11202_));
 sky130_fd_sc_hd__inv_2 _15397_ (.A(_11202_),
    .Y(_00782_));
 sky130_fd_sc_hd__nand2_1 _15398_ (.A(_11152_),
    .B(net3565),
    .Y(_11203_));
 sky130_fd_sc_hd__a22o_1 _15399_ (.A1(net142),
    .A2(_11169_),
    .B1(_11164_),
    .B2(_11203_),
    .X(_11204_));
 sky130_fd_sc_hd__inv_2 _15400_ (.A(_11204_),
    .Y(_00783_));
 sky130_fd_sc_hd__nor2_2 _15401_ (.A(_11162_),
    .B(_10292_),
    .Y(_11205_));
 sky130_fd_sc_hd__inv_2 _15402_ (.A(_11205_),
    .Y(_11206_));
 sky130_fd_sc_hd__nor2_1 _15403_ (.A(_09166_),
    .B(_11206_),
    .Y(_11207_));
 sky130_fd_sc_hd__clkinv_4 _15404_ (.A(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__buf_4 _15405_ (.A(_11208_),
    .X(_11209_));
 sky130_fd_sc_hd__buf_12 _15406_ (.A(_09179_),
    .X(_11210_));
 sky130_fd_sc_hd__buf_4 _15407_ (.A(_11208_),
    .X(_11211_));
 sky130_fd_sc_hd__nor2_1 _15408_ (.A(_11210_),
    .B(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__a31o_1 _15409_ (.A1(_11182_),
    .A2(net1497),
    .A3(_11209_),
    .B1(_11212_),
    .X(_00768_));
 sky130_fd_sc_hd__nor2_8 _15410_ (.A(_08797_),
    .B(_11206_),
    .Y(_11213_));
 sky130_fd_sc_hd__nand2_1 _15411_ (.A(_11152_),
    .B(net3608),
    .Y(_11214_));
 sky130_fd_sc_hd__a22o_1 _15412_ (.A1(_11213_),
    .A2(_09315_),
    .B1(_11211_),
    .B2(_11214_),
    .X(_11215_));
 sky130_fd_sc_hd__inv_2 _15413_ (.A(_11215_),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2_1 _15414_ (.A(_11152_),
    .B(net3422),
    .Y(_11216_));
 sky130_fd_sc_hd__a22o_1 _15415_ (.A1(_11213_),
    .A2(_09460_),
    .B1(_11211_),
    .B2(_11216_),
    .X(_11217_));
 sky130_fd_sc_hd__inv_2 _15416_ (.A(_11217_),
    .Y(_00770_));
 sky130_fd_sc_hd__and3_1 _15417_ (.A(_11205_),
    .B(_11040_),
    .C(_11074_),
    .X(_11218_));
 sky130_fd_sc_hd__a31o_1 _15418_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net2053),
    .B1(_11218_),
    .X(_00771_));
 sky130_fd_sc_hd__clkbuf_16 _15419_ (.A(_09225_),
    .X(_11219_));
 sky130_fd_sc_hd__clkbuf_4 _15420_ (.A(_11219_),
    .X(_11220_));
 sky130_fd_sc_hd__and3_1 _15421_ (.A(_11205_),
    .B(_10587_),
    .C(_11220_),
    .X(_11221_));
 sky130_fd_sc_hd__a31o_1 _15422_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net2213),
    .B1(_11221_),
    .X(_00772_));
 sky130_fd_sc_hd__nand2_1 _15423_ (.A(_11152_),
    .B(net3279),
    .Y(_11222_));
 sky130_fd_sc_hd__a22o_1 _15424_ (.A1(_11213_),
    .A2(_10869_),
    .B1(_11211_),
    .B2(_11222_),
    .X(_11223_));
 sky130_fd_sc_hd__inv_2 _15425_ (.A(_11223_),
    .Y(_00773_));
 sky130_fd_sc_hd__nand2_1 _15426_ (.A(_11152_),
    .B(net3162),
    .Y(_11224_));
 sky130_fd_sc_hd__a22o_1 _15427_ (.A1(_11213_),
    .A2(_11105_),
    .B1(_11211_),
    .B2(_11224_),
    .X(_11225_));
 sky130_fd_sc_hd__inv_2 _15428_ (.A(_11225_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _15429_ (.A(_11152_),
    .B(net3045),
    .Y(_11226_));
 sky130_fd_sc_hd__a22o_1 _15430_ (.A1(_11213_),
    .A2(_10591_),
    .B1(_11211_),
    .B2(_11226_),
    .X(_11227_));
 sky130_fd_sc_hd__inv_2 _15431_ (.A(_11227_),
    .Y(_00775_));
 sky130_fd_sc_hd__nor2_1 _15432_ (.A(_10760_),
    .B(_11211_),
    .Y(_11228_));
 sky130_fd_sc_hd__a31o_1 _15433_ (.A1(_11182_),
    .A2(net467),
    .A3(_11209_),
    .B1(_11228_),
    .X(_00760_));
 sky130_fd_sc_hd__nand2_1 _15434_ (.A(_11152_),
    .B(net3133),
    .Y(_11229_));
 sky130_fd_sc_hd__a22o_1 _15435_ (.A1(_11213_),
    .A2(_10122_),
    .B1(_11208_),
    .B2(_11229_),
    .X(_11230_));
 sky130_fd_sc_hd__inv_2 _15436_ (.A(_11230_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2_1 _15437_ (.A(_11152_),
    .B(net2894),
    .Y(_11231_));
 sky130_fd_sc_hd__a22o_1 _15438_ (.A1(_11213_),
    .A2(_10195_),
    .B1(_11208_),
    .B2(_11231_),
    .X(_11232_));
 sky130_fd_sc_hd__inv_2 _15439_ (.A(_11232_),
    .Y(_00762_));
 sky130_fd_sc_hd__nor2_1 _15440_ (.A(_10657_),
    .B(_11211_),
    .Y(_11233_));
 sky130_fd_sc_hd__a31o_1 _15441_ (.A1(_11182_),
    .A2(net2610),
    .A3(_11209_),
    .B1(_11233_),
    .X(_00763_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(_11152_),
    .B(net3257),
    .Y(_11234_));
 sky130_fd_sc_hd__a22o_1 _15443_ (.A1(_11213_),
    .A2(_09593_),
    .B1(_11208_),
    .B2(_11234_),
    .X(_11235_));
 sky130_fd_sc_hd__inv_2 _15444_ (.A(_11235_),
    .Y(_00764_));
 sky130_fd_sc_hd__nor2_1 _15445_ (.A(_10602_),
    .B(_11211_),
    .Y(_11236_));
 sky130_fd_sc_hd__a31o_1 _15446_ (.A1(_11182_),
    .A2(net2554),
    .A3(_11209_),
    .B1(_11236_),
    .X(_00765_));
 sky130_fd_sc_hd__and3_1 _15447_ (.A(_11205_),
    .B(_09341_),
    .C(_11220_),
    .X(_11237_));
 sky130_fd_sc_hd__a31o_1 _15448_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net2111),
    .B1(_11237_),
    .X(_00766_));
 sky130_fd_sc_hd__buf_4 _15449_ (.A(_10864_),
    .X(_11238_));
 sky130_fd_sc_hd__nor2_1 _15450_ (.A(_10663_),
    .B(_11211_),
    .Y(_11239_));
 sky130_fd_sc_hd__a31o_1 _15451_ (.A1(_11238_),
    .A2(net2333),
    .A3(_11209_),
    .B1(_11239_),
    .X(_00767_));
 sky130_fd_sc_hd__nor2_1 _15452_ (.A(_11002_),
    .B(_11211_),
    .Y(_11240_));
 sky130_fd_sc_hd__a31o_1 _15453_ (.A1(_11238_),
    .A2(net1371),
    .A3(_11209_),
    .B1(_11240_),
    .X(_00752_));
 sky130_fd_sc_hd__and3_1 _15454_ (.A(_11205_),
    .B(_10667_),
    .C(_11220_),
    .X(_11241_));
 sky130_fd_sc_hd__a31o_1 _15455_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net1810),
    .B1(_11241_),
    .X(_00753_));
 sky130_fd_sc_hd__nand2_1 _15456_ (.A(_11152_),
    .B(net3277),
    .Y(_11242_));
 sky130_fd_sc_hd__a22o_1 _15457_ (.A1(_11213_),
    .A2(_09348_),
    .B1(_11208_),
    .B2(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__inv_2 _15458_ (.A(_11243_),
    .Y(_00754_));
 sky130_fd_sc_hd__and3_1 _15459_ (.A(_11205_),
    .B(_10500_),
    .C(_11220_),
    .X(_11244_));
 sky130_fd_sc_hd__a31o_1 _15460_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net2245),
    .B1(_11244_),
    .X(_00755_));
 sky130_fd_sc_hd__nor2_1 _15461_ (.A(_11010_),
    .B(_11211_),
    .Y(_11245_));
 sky130_fd_sc_hd__a31o_1 _15462_ (.A1(_11238_),
    .A2(net1789),
    .A3(_11209_),
    .B1(_11245_),
    .X(_00756_));
 sky130_fd_sc_hd__nand2_1 _15463_ (.A(_11152_),
    .B(net3225),
    .Y(_11246_));
 sky130_fd_sc_hd__a22o_1 _15464_ (.A1(_11213_),
    .A2(_10149_),
    .B1(_11208_),
    .B2(_11246_),
    .X(_11247_));
 sky130_fd_sc_hd__inv_2 _15465_ (.A(_11247_),
    .Y(_00757_));
 sky130_fd_sc_hd__and3_1 _15466_ (.A(_11205_),
    .B(_10617_),
    .C(_11220_),
    .X(_11248_));
 sky130_fd_sc_hd__a31o_1 _15467_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net1786),
    .B1(_11248_),
    .X(_00758_));
 sky130_fd_sc_hd__nand2_1 _15468_ (.A(_11152_),
    .B(net2962),
    .Y(_11249_));
 sky130_fd_sc_hd__a22o_1 _15469_ (.A1(_11213_),
    .A2(_10154_),
    .B1(_11208_),
    .B2(_11249_),
    .X(_11250_));
 sky130_fd_sc_hd__inv_2 _15470_ (.A(_11250_),
    .Y(_00759_));
 sky130_fd_sc_hd__buf_4 _15471_ (.A(_11151_),
    .X(_11251_));
 sky130_fd_sc_hd__nand2_1 _15472_ (.A(_11251_),
    .B(net3291),
    .Y(_11252_));
 sky130_fd_sc_hd__a22o_1 _15473_ (.A1(_11213_),
    .A2(_09495_),
    .B1(_11208_),
    .B2(_11252_),
    .X(_11253_));
 sky130_fd_sc_hd__inv_2 _15474_ (.A(_11253_),
    .Y(_00744_));
 sky130_fd_sc_hd__nor2_1 _15475_ (.A(_10681_),
    .B(_11211_),
    .Y(_11254_));
 sky130_fd_sc_hd__a31o_1 _15476_ (.A1(_11238_),
    .A2(net2013),
    .A3(_11211_),
    .B1(_11254_),
    .X(_00745_));
 sky130_fd_sc_hd__and3_1 _15477_ (.A(_11205_),
    .B(_10728_),
    .C(_11220_),
    .X(_11255_));
 sky130_fd_sc_hd__a31o_1 _15478_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net2283),
    .B1(_11255_),
    .X(_00746_));
 sky130_fd_sc_hd__nand2_1 _15479_ (.A(_11251_),
    .B(net3319),
    .Y(_11256_));
 sky130_fd_sc_hd__a22o_1 _15480_ (.A1(_11213_),
    .A2(_10164_),
    .B1(_11208_),
    .B2(_11256_),
    .X(_11257_));
 sky130_fd_sc_hd__inv_2 _15481_ (.A(_11257_),
    .Y(_00747_));
 sky130_fd_sc_hd__and3_1 _15482_ (.A(_11205_),
    .B(_10848_),
    .C(_11220_),
    .X(_11258_));
 sky130_fd_sc_hd__a31o_1 _15483_ (.A1(_11209_),
    .A2(_11082_),
    .A3(net2066),
    .B1(_11258_),
    .X(_00748_));
 sky130_fd_sc_hd__nand2_1 _15484_ (.A(_11251_),
    .B(net3156),
    .Y(_11259_));
 sky130_fd_sc_hd__a22o_1 _15485_ (.A1(_11213_),
    .A2(net136),
    .B1(_11208_),
    .B2(_11259_),
    .X(_11260_));
 sky130_fd_sc_hd__inv_2 _15486_ (.A(_11260_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand2_1 _15487_ (.A(_11174_),
    .B(net3935),
    .Y(_11261_));
 sky130_fd_sc_hd__o2bb2a_1 _15488_ (.A1_N(_11261_),
    .A2_N(_11209_),
    .B1(_10289_),
    .B2(_11206_),
    .X(_00750_));
 sky130_fd_sc_hd__nor2_1 _15489_ (.A(_09300_),
    .B(_11211_),
    .Y(_11262_));
 sky130_fd_sc_hd__a31o_1 _15490_ (.A1(_11238_),
    .A2(net805),
    .A3(_11211_),
    .B1(_11262_),
    .X(_00751_));
 sky130_fd_sc_hd__nor2_2 _15491_ (.A(_11162_),
    .B(_10356_),
    .Y(_11263_));
 sky130_fd_sc_hd__inv_2 _15492_ (.A(_11263_),
    .Y(_11264_));
 sky130_fd_sc_hd__nor2_4 _15493_ (.A(_09190_),
    .B(_11264_),
    .Y(_11265_));
 sky130_fd_sc_hd__nor2_1 _15494_ (.A(_09304_),
    .B(_11264_),
    .Y(_11266_));
 sky130_fd_sc_hd__inv_2 _15495_ (.A(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__buf_4 _15496_ (.A(_11267_),
    .X(_11268_));
 sky130_fd_sc_hd__nand2_1 _15497_ (.A(_11251_),
    .B(net2890),
    .Y(_11269_));
 sky130_fd_sc_hd__a22o_1 _15498_ (.A1(_11265_),
    .A2(_10239_),
    .B1(_11268_),
    .B2(_11269_),
    .X(_11270_));
 sky130_fd_sc_hd__inv_2 _15499_ (.A(_11270_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand2_1 _15500_ (.A(_11251_),
    .B(net2911),
    .Y(_11271_));
 sky130_fd_sc_hd__a22o_1 _15501_ (.A1(_11265_),
    .A2(_09315_),
    .B1(_11268_),
    .B2(_11271_),
    .X(_11272_));
 sky130_fd_sc_hd__inv_2 _15502_ (.A(_11272_),
    .Y(_00737_));
 sky130_fd_sc_hd__buf_4 _15503_ (.A(_11267_),
    .X(_11273_));
 sky130_fd_sc_hd__nor2_1 _15504_ (.A(_10698_),
    .B(_11268_),
    .Y(_11274_));
 sky130_fd_sc_hd__a31o_1 _15505_ (.A1(_11238_),
    .A2(net1800),
    .A3(_11273_),
    .B1(_11274_),
    .X(_00738_));
 sky130_fd_sc_hd__nand2_1 _15506_ (.A(_11251_),
    .B(net3690),
    .Y(_11275_));
 sky130_fd_sc_hd__a22o_1 _15507_ (.A1(_11265_),
    .A2(_10983_),
    .B1(_11268_),
    .B2(_11275_),
    .X(_11276_));
 sky130_fd_sc_hd__inv_2 _15508_ (.A(_11276_),
    .Y(_00739_));
 sky130_fd_sc_hd__and3_1 _15509_ (.A(_11263_),
    .B(_10587_),
    .C(_11220_),
    .X(_11277_));
 sky130_fd_sc_hd__a31o_1 _15510_ (.A1(_11273_),
    .A2(_11082_),
    .A3(net2449),
    .B1(_11277_),
    .X(_00740_));
 sky130_fd_sc_hd__nand2_1 _15511_ (.A(_11251_),
    .B(net3859),
    .Y(_11278_));
 sky130_fd_sc_hd__a22o_1 _15512_ (.A1(_11265_),
    .A2(_10869_),
    .B1(_11267_),
    .B2(_11278_),
    .X(_11279_));
 sky130_fd_sc_hd__inv_2 _15513_ (.A(_11279_),
    .Y(_00741_));
 sky130_fd_sc_hd__nor2_1 _15514_ (.A(_10872_),
    .B(_11268_),
    .Y(_11280_));
 sky130_fd_sc_hd__a31o_1 _15515_ (.A1(_11238_),
    .A2(net2303),
    .A3(_11273_),
    .B1(_11280_),
    .X(_00742_));
 sky130_fd_sc_hd__and3_1 _15516_ (.A(_11263_),
    .B(_10874_),
    .C(_11220_),
    .X(_11281_));
 sky130_fd_sc_hd__a31o_1 _15517_ (.A1(_11273_),
    .A2(_11082_),
    .A3(net2413),
    .B1(_11281_),
    .X(_00743_));
 sky130_fd_sc_hd__nor2_1 _15518_ (.A(_10760_),
    .B(_11268_),
    .Y(_11282_));
 sky130_fd_sc_hd__a31o_1 _15519_ (.A1(_11238_),
    .A2(net1183),
    .A3(_11273_),
    .B1(_11282_),
    .X(_00728_));
 sky130_fd_sc_hd__nand2_1 _15520_ (.A(_11251_),
    .B(net3037),
    .Y(_11283_));
 sky130_fd_sc_hd__a22o_1 _15521_ (.A1(_11265_),
    .A2(_10122_),
    .B1(_11267_),
    .B2(_11283_),
    .X(_11284_));
 sky130_fd_sc_hd__inv_2 _15522_ (.A(_11284_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _15523_ (.A(_11251_),
    .B(net2935),
    .Y(_11285_));
 sky130_fd_sc_hd__a22o_1 _15524_ (.A1(_11265_),
    .A2(_10195_),
    .B1(_11267_),
    .B2(_11285_),
    .X(_11286_));
 sky130_fd_sc_hd__inv_2 _15525_ (.A(_11286_),
    .Y(_00730_));
 sky130_fd_sc_hd__nor2_1 _15526_ (.A(_10657_),
    .B(_11268_),
    .Y(_11287_));
 sky130_fd_sc_hd__a31o_1 _15527_ (.A1(_11238_),
    .A2(net2612),
    .A3(_11273_),
    .B1(_11287_),
    .X(_00731_));
 sky130_fd_sc_hd__nor2_1 _15528_ (.A(_10767_),
    .B(_11268_),
    .Y(_11288_));
 sky130_fd_sc_hd__a31o_1 _15529_ (.A1(_11238_),
    .A2(net2255),
    .A3(_11273_),
    .B1(_11288_),
    .X(_00732_));
 sky130_fd_sc_hd__nand2_1 _15530_ (.A(_11251_),
    .B(net3787),
    .Y(_11289_));
 sky130_fd_sc_hd__a22o_1 _15531_ (.A1(_11265_),
    .A2(_09338_),
    .B1(_11267_),
    .B2(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__inv_2 _15532_ (.A(_11290_),
    .Y(_00733_));
 sky130_fd_sc_hd__buf_8 _15533_ (.A(net64),
    .X(_11291_));
 sky130_fd_sc_hd__and3_1 _15534_ (.A(_11263_),
    .B(_11291_),
    .C(_11220_),
    .X(_11292_));
 sky130_fd_sc_hd__a31o_1 _15535_ (.A1(_11273_),
    .A2(_11082_),
    .A3(net2530),
    .B1(_11292_),
    .X(_00734_));
 sky130_fd_sc_hd__nor2_1 _15536_ (.A(_10663_),
    .B(_11268_),
    .Y(_11293_));
 sky130_fd_sc_hd__a31o_1 _15537_ (.A1(_11238_),
    .A2(net1938),
    .A3(_11268_),
    .B1(_11293_),
    .X(_00735_));
 sky130_fd_sc_hd__nor2_1 _15538_ (.A(_11002_),
    .B(_11268_),
    .Y(_11294_));
 sky130_fd_sc_hd__a31o_1 _15539_ (.A1(_11238_),
    .A2(net2189),
    .A3(_11268_),
    .B1(_11294_),
    .X(_00720_));
 sky130_fd_sc_hd__nand2_1 _15540_ (.A(_11251_),
    .B(net3290),
    .Y(_11295_));
 sky130_fd_sc_hd__a22o_1 _15541_ (.A1(_11265_),
    .A2(_09249_),
    .B1(_11267_),
    .B2(_11295_),
    .X(_11296_));
 sky130_fd_sc_hd__inv_2 _15542_ (.A(_11296_),
    .Y(_00721_));
 sky130_fd_sc_hd__nor2_1 _15543_ (.A(_10669_),
    .B(_11268_),
    .Y(_11297_));
 sky130_fd_sc_hd__a31o_1 _15544_ (.A1(_11238_),
    .A2(net1369),
    .A3(_11268_),
    .B1(_11297_),
    .X(_00722_));
 sky130_fd_sc_hd__and3_1 _15545_ (.A(_11263_),
    .B(_10500_),
    .C(_11220_),
    .X(_11298_));
 sky130_fd_sc_hd__a31o_1 _15546_ (.A1(_11273_),
    .A2(_11082_),
    .A3(net2368),
    .B1(_11298_),
    .X(_00723_));
 sky130_fd_sc_hd__nand2_1 _15547_ (.A(_11251_),
    .B(net3171),
    .Y(_11299_));
 sky130_fd_sc_hd__a22o_1 _15548_ (.A1(_11265_),
    .A2(_11136_),
    .B1(_11267_),
    .B2(_11299_),
    .X(_11300_));
 sky130_fd_sc_hd__inv_2 _15549_ (.A(_11300_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _15550_ (.A(_11251_),
    .B(net3394),
    .Y(_11301_));
 sky130_fd_sc_hd__a22o_1 _15551_ (.A1(_11265_),
    .A2(_10149_),
    .B1(_11267_),
    .B2(_11301_),
    .X(_11302_));
 sky130_fd_sc_hd__inv_2 _15552_ (.A(_11302_),
    .Y(_00725_));
 sky130_fd_sc_hd__and3_1 _15553_ (.A(_11263_),
    .B(_10617_),
    .C(_11220_),
    .X(_11303_));
 sky130_fd_sc_hd__a31o_1 _15554_ (.A1(_11273_),
    .A2(_11082_),
    .A3(net2472),
    .B1(_11303_),
    .X(_00726_));
 sky130_fd_sc_hd__nand2_1 _15555_ (.A(_11251_),
    .B(net3585),
    .Y(_11304_));
 sky130_fd_sc_hd__a22o_1 _15556_ (.A1(_11265_),
    .A2(_10154_),
    .B1(_11267_),
    .B2(_11304_),
    .X(_11305_));
 sky130_fd_sc_hd__inv_2 _15557_ (.A(_11305_),
    .Y(_00727_));
 sky130_fd_sc_hd__and3_1 _15558_ (.A(_11263_),
    .B(_10679_),
    .C(_11220_),
    .X(_11306_));
 sky130_fd_sc_hd__a31o_1 _15559_ (.A1(_11273_),
    .A2(_11082_),
    .A3(net2507),
    .B1(_11306_),
    .X(_00712_));
 sky130_fd_sc_hd__nor2_1 _15560_ (.A(_10681_),
    .B(_11268_),
    .Y(_11307_));
 sky130_fd_sc_hd__a31o_1 _15561_ (.A1(_11238_),
    .A2(net725),
    .A3(_11268_),
    .B1(_11307_),
    .X(_00713_));
 sky130_fd_sc_hd__and3_1 _15562_ (.A(_11263_),
    .B(_10728_),
    .C(_11220_),
    .X(_11308_));
 sky130_fd_sc_hd__a31o_1 _15563_ (.A1(_11273_),
    .A2(_11082_),
    .A3(net2644),
    .B1(_11308_),
    .X(_00714_));
 sky130_fd_sc_hd__nand2_1 _15564_ (.A(_11251_),
    .B(net3421),
    .Y(_11309_));
 sky130_fd_sc_hd__a22o_1 _15565_ (.A1(_11265_),
    .A2(_10164_),
    .B1(_11267_),
    .B2(_11309_),
    .X(_11310_));
 sky130_fd_sc_hd__inv_2 _15566_ (.A(_11310_),
    .Y(_00715_));
 sky130_fd_sc_hd__clkbuf_8 _15567_ (.A(_10645_),
    .X(_11311_));
 sky130_fd_sc_hd__and3_1 _15568_ (.A(_11263_),
    .B(_10848_),
    .C(_11220_),
    .X(_11312_));
 sky130_fd_sc_hd__a31o_1 _15569_ (.A1(_11273_),
    .A2(_11311_),
    .A3(net1612),
    .B1(_11312_),
    .X(_00716_));
 sky130_fd_sc_hd__and3_1 _15570_ (.A(_11263_),
    .B(_09730_),
    .C(_11220_),
    .X(_11313_));
 sky130_fd_sc_hd__a31o_1 _15571_ (.A1(_11273_),
    .A2(_11311_),
    .A3(net1453),
    .B1(_11313_),
    .X(_00717_));
 sky130_fd_sc_hd__nand2_1 _15572_ (.A(_11174_),
    .B(net3884),
    .Y(_11314_));
 sky130_fd_sc_hd__o2bb2a_1 _15573_ (.A1_N(_11314_),
    .A2_N(_11273_),
    .B1(_10289_),
    .B2(_11264_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_1 _15574_ (.A(_11174_),
    .B(net3908),
    .Y(_11315_));
 sky130_fd_sc_hd__clkbuf_16 _15575_ (.A(_09441_),
    .X(_11316_));
 sky130_fd_sc_hd__o2bb2a_1 _15576_ (.A1_N(_11315_),
    .A2_N(_11273_),
    .B1(_11316_),
    .B2(_11264_),
    .X(_00719_));
 sky130_fd_sc_hd__nor2_2 _15577_ (.A(_11162_),
    .B(_10411_),
    .Y(_11317_));
 sky130_fd_sc_hd__inv_2 _15578_ (.A(_11317_),
    .Y(_11318_));
 sky130_fd_sc_hd__nor2_1 _15579_ (.A(_09625_),
    .B(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__inv_2 _15580_ (.A(_11319_),
    .Y(_11320_));
 sky130_fd_sc_hd__buf_4 _15581_ (.A(_11320_),
    .X(_11321_));
 sky130_fd_sc_hd__buf_4 _15582_ (.A(_11320_),
    .X(_11322_));
 sky130_fd_sc_hd__nor2_1 _15583_ (.A(_11210_),
    .B(_11322_),
    .Y(_11323_));
 sky130_fd_sc_hd__a31o_1 _15584_ (.A1(_11238_),
    .A2(net1773),
    .A3(_11321_),
    .B1(_11323_),
    .X(_00696_));
 sky130_fd_sc_hd__nor2_8 _15585_ (.A(_08794_),
    .B(_11318_),
    .Y(_11324_));
 sky130_fd_sc_hd__nand2_1 _15586_ (.A(_11251_),
    .B(net3292),
    .Y(_11325_));
 sky130_fd_sc_hd__a22o_1 _15587_ (.A1(_11324_),
    .A2(_09315_),
    .B1(_11322_),
    .B2(_11325_),
    .X(_11326_));
 sky130_fd_sc_hd__inv_2 _15588_ (.A(_11326_),
    .Y(_00697_));
 sky130_fd_sc_hd__nor2_1 _15589_ (.A(_10698_),
    .B(_11322_),
    .Y(_11327_));
 sky130_fd_sc_hd__a31o_1 _15590_ (.A1(_11238_),
    .A2(net1317),
    .A3(_11321_),
    .B1(_11327_),
    .X(_00698_));
 sky130_fd_sc_hd__buf_4 _15591_ (.A(_11219_),
    .X(_11328_));
 sky130_fd_sc_hd__and3_1 _15592_ (.A(_11317_),
    .B(_11040_),
    .C(_11328_),
    .X(_11329_));
 sky130_fd_sc_hd__a31o_1 _15593_ (.A1(_11321_),
    .A2(_11311_),
    .A3(net2297),
    .B1(_11329_),
    .X(_00699_));
 sky130_fd_sc_hd__buf_12 _15594_ (.A(_09200_),
    .X(_11330_));
 sky130_fd_sc_hd__buf_4 _15595_ (.A(_11151_),
    .X(_11331_));
 sky130_fd_sc_hd__nand2_1 _15596_ (.A(_11331_),
    .B(net3181),
    .Y(_11332_));
 sky130_fd_sc_hd__a22o_1 _15597_ (.A1(_11324_),
    .A2(_11330_),
    .B1(_11322_),
    .B2(_11332_),
    .X(_11333_));
 sky130_fd_sc_hd__inv_2 _15598_ (.A(_11333_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2_1 _15599_ (.A(_11331_),
    .B(net2994),
    .Y(_11334_));
 sky130_fd_sc_hd__a22o_1 _15600_ (.A1(_11324_),
    .A2(_10869_),
    .B1(_11322_),
    .B2(_11334_),
    .X(_11335_));
 sky130_fd_sc_hd__inv_2 _15601_ (.A(_11335_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand2_1 _15602_ (.A(_11331_),
    .B(net3041),
    .Y(_11336_));
 sky130_fd_sc_hd__a22o_1 _15603_ (.A1(_11324_),
    .A2(_11105_),
    .B1(_11322_),
    .B2(_11336_),
    .X(_11337_));
 sky130_fd_sc_hd__inv_2 _15604_ (.A(_11337_),
    .Y(_00702_));
 sky130_fd_sc_hd__and3_1 _15605_ (.A(_11317_),
    .B(_10874_),
    .C(_11328_),
    .X(_11338_));
 sky130_fd_sc_hd__a31o_1 _15606_ (.A1(_11321_),
    .A2(_11311_),
    .A3(net2434),
    .B1(_11338_),
    .X(_00703_));
 sky130_fd_sc_hd__nand2_1 _15607_ (.A(_11331_),
    .B(net3131),
    .Y(_11339_));
 sky130_fd_sc_hd__a22o_1 _15608_ (.A1(_11324_),
    .A2(net135),
    .B1(_11322_),
    .B2(_11339_),
    .X(_11340_));
 sky130_fd_sc_hd__inv_2 _15609_ (.A(_11340_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _15610_ (.A(_11331_),
    .B(net3323),
    .Y(_11341_));
 sky130_fd_sc_hd__a22o_1 _15611_ (.A1(_11324_),
    .A2(_10122_),
    .B1(_11322_),
    .B2(_11341_),
    .X(_11342_));
 sky130_fd_sc_hd__inv_2 _15612_ (.A(_11342_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _15613_ (.A(_11331_),
    .B(net3080),
    .Y(_11343_));
 sky130_fd_sc_hd__a22o_1 _15614_ (.A1(_11324_),
    .A2(_10195_),
    .B1(_11322_),
    .B2(_11343_),
    .X(_11344_));
 sky130_fd_sc_hd__inv_2 _15615_ (.A(_11344_),
    .Y(_00690_));
 sky130_fd_sc_hd__clkbuf_8 _15616_ (.A(_10864_),
    .X(_11345_));
 sky130_fd_sc_hd__nor2_1 _15617_ (.A(_10657_),
    .B(_11322_),
    .Y(_11346_));
 sky130_fd_sc_hd__a31o_1 _15618_ (.A1(_11345_),
    .A2(net2024),
    .A3(_11321_),
    .B1(_11346_),
    .X(_00691_));
 sky130_fd_sc_hd__nor2_1 _15619_ (.A(_10767_),
    .B(_11322_),
    .Y(_11347_));
 sky130_fd_sc_hd__a31o_1 _15620_ (.A1(_11345_),
    .A2(net1391),
    .A3(_11321_),
    .B1(_11347_),
    .X(_00692_));
 sky130_fd_sc_hd__nor2_1 _15621_ (.A(_10602_),
    .B(_11322_),
    .Y(_11348_));
 sky130_fd_sc_hd__a31o_1 _15622_ (.A1(_11345_),
    .A2(net1033),
    .A3(_11321_),
    .B1(_11348_),
    .X(_00693_));
 sky130_fd_sc_hd__nand2_1 _15623_ (.A(_11331_),
    .B(net3381),
    .Y(_11349_));
 sky130_fd_sc_hd__a22o_1 _15624_ (.A1(_11324_),
    .A2(_10202_),
    .B1(_11320_),
    .B2(_11349_),
    .X(_11350_));
 sky130_fd_sc_hd__inv_2 _15625_ (.A(_11350_),
    .Y(_00694_));
 sky130_fd_sc_hd__nor2_1 _15626_ (.A(_10663_),
    .B(_11322_),
    .Y(_11351_));
 sky130_fd_sc_hd__a31o_1 _15627_ (.A1(_11345_),
    .A2(net1493),
    .A3(_11321_),
    .B1(_11351_),
    .X(_00695_));
 sky130_fd_sc_hd__nor2_1 _15628_ (.A(_11002_),
    .B(_11322_),
    .Y(_11352_));
 sky130_fd_sc_hd__a31o_1 _15629_ (.A1(_11345_),
    .A2(net927),
    .A3(_11321_),
    .B1(_11352_),
    .X(_00680_));
 sky130_fd_sc_hd__and3_1 _15630_ (.A(_11317_),
    .B(_10667_),
    .C(_11328_),
    .X(_11353_));
 sky130_fd_sc_hd__a31o_1 _15631_ (.A1(_11321_),
    .A2(_11311_),
    .A3(net2502),
    .B1(_11353_),
    .X(_00681_));
 sky130_fd_sc_hd__nor2_1 _15632_ (.A(_10669_),
    .B(_11322_),
    .Y(_11354_));
 sky130_fd_sc_hd__a31o_1 _15633_ (.A1(_11345_),
    .A2(net813),
    .A3(_11321_),
    .B1(_11354_),
    .X(_00682_));
 sky130_fd_sc_hd__and3_1 _15634_ (.A(_11317_),
    .B(_10500_),
    .C(_11328_),
    .X(_11355_));
 sky130_fd_sc_hd__a31o_1 _15635_ (.A1(_11321_),
    .A2(_11311_),
    .A3(net1870),
    .B1(_11355_),
    .X(_00683_));
 sky130_fd_sc_hd__nor2_1 _15636_ (.A(_11010_),
    .B(_11322_),
    .Y(_11356_));
 sky130_fd_sc_hd__a31o_1 _15637_ (.A1(_11345_),
    .A2(net1073),
    .A3(_11321_),
    .B1(_11356_),
    .X(_00684_));
 sky130_fd_sc_hd__nand2_1 _15638_ (.A(_11331_),
    .B(net2943),
    .Y(_11357_));
 sky130_fd_sc_hd__a22o_1 _15639_ (.A1(_11324_),
    .A2(_10149_),
    .B1(_11320_),
    .B2(_11357_),
    .X(_11358_));
 sky130_fd_sc_hd__inv_2 _15640_ (.A(_11358_),
    .Y(_00685_));
 sky130_fd_sc_hd__and3_1 _15641_ (.A(_11317_),
    .B(_10617_),
    .C(_11328_),
    .X(_11359_));
 sky130_fd_sc_hd__a31o_1 _15642_ (.A1(_11321_),
    .A2(_11311_),
    .A3(net1861),
    .B1(_11359_),
    .X(_00686_));
 sky130_fd_sc_hd__nand2_1 _15643_ (.A(_11331_),
    .B(net3479),
    .Y(_11360_));
 sky130_fd_sc_hd__a22o_1 _15644_ (.A1(_11324_),
    .A2(_10154_),
    .B1(_11320_),
    .B2(_11360_),
    .X(_11361_));
 sky130_fd_sc_hd__inv_2 _15645_ (.A(_11361_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand2_1 _15646_ (.A(_11331_),
    .B(net3139),
    .Y(_11362_));
 sky130_fd_sc_hd__a22o_1 _15647_ (.A1(_11324_),
    .A2(net141),
    .B1(_11320_),
    .B2(_11362_),
    .X(_11363_));
 sky130_fd_sc_hd__inv_2 _15648_ (.A(_11363_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _15649_ (.A(_11331_),
    .B(net3242),
    .Y(_11364_));
 sky130_fd_sc_hd__a22o_1 _15650_ (.A1(_11324_),
    .A2(_09366_),
    .B1(_11320_),
    .B2(_11364_),
    .X(_11365_));
 sky130_fd_sc_hd__inv_2 _15651_ (.A(_11365_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand2_1 _15652_ (.A(_11331_),
    .B(net3276),
    .Y(_11366_));
 sky130_fd_sc_hd__a22o_1 _15653_ (.A1(_11324_),
    .A2(_10624_),
    .B1(_11320_),
    .B2(_11366_),
    .X(_11367_));
 sky130_fd_sc_hd__inv_2 _15654_ (.A(_11367_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _15655_ (.A(_11331_),
    .B(net3063),
    .Y(_11368_));
 sky130_fd_sc_hd__a22o_1 _15656_ (.A1(_11324_),
    .A2(_10164_),
    .B1(_11320_),
    .B2(_11368_),
    .X(_11369_));
 sky130_fd_sc_hd__inv_2 _15657_ (.A(_11369_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_1 _15658_ (.A(_11331_),
    .B(net2899),
    .Y(_11370_));
 sky130_fd_sc_hd__a22o_1 _15659_ (.A1(_11324_),
    .A2(net139),
    .B1(_11320_),
    .B2(_11370_),
    .X(_11371_));
 sky130_fd_sc_hd__inv_2 _15660_ (.A(_11371_),
    .Y(_00676_));
 sky130_fd_sc_hd__nand2_1 _15661_ (.A(_11331_),
    .B(net3359),
    .Y(_11372_));
 sky130_fd_sc_hd__a22o_1 _15662_ (.A1(_11324_),
    .A2(net136),
    .B1(_11320_),
    .B2(_11372_),
    .X(_11373_));
 sky130_fd_sc_hd__inv_2 _15663_ (.A(_11373_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _15664_ (.A(_11174_),
    .B(net3726),
    .Y(_11374_));
 sky130_fd_sc_hd__o2bb2a_1 _15665_ (.A1_N(_11374_),
    .A2_N(_11321_),
    .B1(_10289_),
    .B2(_11318_),
    .X(_00678_));
 sky130_fd_sc_hd__nand2_1 _15666_ (.A(_11174_),
    .B(net3745),
    .Y(_11375_));
 sky130_fd_sc_hd__o2bb2a_1 _15667_ (.A1_N(_11375_),
    .A2_N(_11321_),
    .B1(_11316_),
    .B2(_11318_),
    .X(_00679_));
 sky130_fd_sc_hd__nand2_8 _15668_ (.A(_09509_),
    .B(_11161_),
    .Y(_11376_));
 sky130_fd_sc_hd__nor2_4 _15669_ (.A(_10469_),
    .B(_11376_),
    .Y(_11377_));
 sky130_fd_sc_hd__nand2_4 _15670_ (.A(_11377_),
    .B(_10413_),
    .Y(_11378_));
 sky130_fd_sc_hd__buf_4 _15671_ (.A(_11378_),
    .X(_11379_));
 sky130_fd_sc_hd__buf_4 _15672_ (.A(_11378_),
    .X(_11380_));
 sky130_fd_sc_hd__nor2_1 _15673_ (.A(_11210_),
    .B(_11380_),
    .Y(_11381_));
 sky130_fd_sc_hd__a31o_1 _15674_ (.A1(_11345_),
    .A2(net2690),
    .A3(_11379_),
    .B1(_11381_),
    .X(_00664_));
 sky130_fd_sc_hd__nand2_1 _15675_ (.A(_10931_),
    .B(net4264),
    .Y(_11382_));
 sky130_fd_sc_hd__and2_1 _15676_ (.A(_11377_),
    .B(_08778_),
    .X(_11383_));
 sky130_fd_sc_hd__clkbuf_4 _15677_ (.A(_11383_),
    .X(_11384_));
 sky130_fd_sc_hd__a22o_1 _15678_ (.A1(_11380_),
    .A2(_11382_),
    .B1(_11384_),
    .B2(_09315_),
    .X(_11385_));
 sky130_fd_sc_hd__inv_2 _15679_ (.A(_11385_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _15680_ (.A(_10931_),
    .B(net4148),
    .Y(_11386_));
 sky130_fd_sc_hd__a22o_1 _15681_ (.A1(_11378_),
    .A2(_11386_),
    .B1(_11384_),
    .B2(_09460_),
    .X(_11387_));
 sky130_fd_sc_hd__inv_2 _15682_ (.A(_11387_),
    .Y(_00666_));
 sky130_fd_sc_hd__and3_1 _15683_ (.A(_11377_),
    .B(_11040_),
    .C(_11328_),
    .X(_11388_));
 sky130_fd_sc_hd__a31o_1 _15684_ (.A1(_11345_),
    .A2(net1289),
    .A3(_11379_),
    .B1(_11388_),
    .X(_00667_));
 sky130_fd_sc_hd__nand2_1 _15685_ (.A(_10931_),
    .B(net4268),
    .Y(_11389_));
 sky130_fd_sc_hd__a22o_1 _15686_ (.A1(_11378_),
    .A2(_11389_),
    .B1(_11384_),
    .B2(_09201_),
    .X(_11390_));
 sky130_fd_sc_hd__inv_2 _15687_ (.A(_11390_),
    .Y(_00668_));
 sky130_fd_sc_hd__clkbuf_16 _15688_ (.A(net71),
    .X(_11391_));
 sky130_fd_sc_hd__and3_1 _15689_ (.A(_11377_),
    .B(_11391_),
    .C(_11328_),
    .X(_11392_));
 sky130_fd_sc_hd__a31o_1 _15690_ (.A1(_11345_),
    .A2(net1715),
    .A3(_11379_),
    .B1(_11392_),
    .X(_00669_));
 sky130_fd_sc_hd__nor2_1 _15691_ (.A(_10872_),
    .B(_11380_),
    .Y(_11393_));
 sky130_fd_sc_hd__a31o_1 _15692_ (.A1(_11345_),
    .A2(net641),
    .A3(_11379_),
    .B1(_11393_),
    .X(_00670_));
 sky130_fd_sc_hd__and3_1 _15693_ (.A(_11377_),
    .B(_10874_),
    .C(_11328_),
    .X(_11394_));
 sky130_fd_sc_hd__a31o_1 _15694_ (.A1(_11345_),
    .A2(net1091),
    .A3(_11379_),
    .B1(_11394_),
    .X(_00671_));
 sky130_fd_sc_hd__buf_4 _15695_ (.A(_10930_),
    .X(_11395_));
 sky130_fd_sc_hd__nand2_1 _15696_ (.A(_11395_),
    .B(net4192),
    .Y(_11396_));
 sky130_fd_sc_hd__a22o_1 _15697_ (.A1(_11378_),
    .A2(_11396_),
    .B1(_11384_),
    .B2(_09531_),
    .X(_11397_));
 sky130_fd_sc_hd__inv_2 _15698_ (.A(_11397_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand2_1 _15699_ (.A(_11395_),
    .B(net4262),
    .Y(_11398_));
 sky130_fd_sc_hd__a22o_1 _15700_ (.A1(_11378_),
    .A2(_11398_),
    .B1(_11384_),
    .B2(_10313_),
    .X(_11399_));
 sky130_fd_sc_hd__inv_2 _15701_ (.A(_11399_),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2_1 _15702_ (.A(_11395_),
    .B(net4099),
    .Y(_11400_));
 sky130_fd_sc_hd__a22o_1 _15703_ (.A1(_11378_),
    .A2(_11400_),
    .B1(_11384_),
    .B2(_10316_),
    .X(_11401_));
 sky130_fd_sc_hd__inv_2 _15704_ (.A(_11401_),
    .Y(_00658_));
 sky130_fd_sc_hd__nor2_1 _15705_ (.A(_10657_),
    .B(_11380_),
    .Y(_11402_));
 sky130_fd_sc_hd__a31o_1 _15706_ (.A1(_11345_),
    .A2(net1065),
    .A3(_11379_),
    .B1(_11402_),
    .X(_00659_));
 sky130_fd_sc_hd__nor2_1 _15707_ (.A(_10767_),
    .B(_11380_),
    .Y(_11403_));
 sky130_fd_sc_hd__a31o_1 _15708_ (.A1(_11345_),
    .A2(net1599),
    .A3(_11379_),
    .B1(_11403_),
    .X(_00660_));
 sky130_fd_sc_hd__nor2_1 _15709_ (.A(_10602_),
    .B(_11380_),
    .Y(_11404_));
 sky130_fd_sc_hd__a31o_1 _15710_ (.A1(_11345_),
    .A2(net1571),
    .A3(_11379_),
    .B1(_11404_),
    .X(_00661_));
 sky130_fd_sc_hd__and3_1 _15711_ (.A(_11377_),
    .B(_11291_),
    .C(_11328_),
    .X(_11405_));
 sky130_fd_sc_hd__a31o_1 _15712_ (.A1(_11345_),
    .A2(net1751),
    .A3(_11379_),
    .B1(_11405_),
    .X(_00662_));
 sky130_fd_sc_hd__nand2_1 _15713_ (.A(_11395_),
    .B(net4181),
    .Y(_11406_));
 sky130_fd_sc_hd__a22o_1 _15714_ (.A1(_11378_),
    .A2(_11406_),
    .B1(_11384_),
    .B2(_09768_),
    .X(_11407_));
 sky130_fd_sc_hd__inv_2 _15715_ (.A(_11407_),
    .Y(_00663_));
 sky130_fd_sc_hd__clkbuf_8 _15716_ (.A(_10864_),
    .X(_11408_));
 sky130_fd_sc_hd__nor2_1 _15717_ (.A(_11002_),
    .B(_11380_),
    .Y(_11409_));
 sky130_fd_sc_hd__a31o_1 _15718_ (.A1(_11408_),
    .A2(net1513),
    .A3(_11379_),
    .B1(_11409_),
    .X(_00648_));
 sky130_fd_sc_hd__and3_1 _15719_ (.A(_11377_),
    .B(_10667_),
    .C(_11328_),
    .X(_11410_));
 sky130_fd_sc_hd__a31o_1 _15720_ (.A1(_11408_),
    .A2(net1966),
    .A3(_11379_),
    .B1(_11410_),
    .X(_00649_));
 sky130_fd_sc_hd__nor2_1 _15721_ (.A(_10669_),
    .B(_11380_),
    .Y(_11411_));
 sky130_fd_sc_hd__a31o_1 _15722_ (.A1(_11408_),
    .A2(net793),
    .A3(_11379_),
    .B1(_11411_),
    .X(_00650_));
 sky130_fd_sc_hd__and3_1 _15723_ (.A(_11377_),
    .B(_10500_),
    .C(_11328_),
    .X(_11412_));
 sky130_fd_sc_hd__a31o_1 _15724_ (.A1(_11408_),
    .A2(net747),
    .A3(_11379_),
    .B1(_11412_),
    .X(_00651_));
 sky130_fd_sc_hd__nor2_1 _15725_ (.A(_11010_),
    .B(_11380_),
    .Y(_11413_));
 sky130_fd_sc_hd__a31o_1 _15726_ (.A1(_11408_),
    .A2(net1481),
    .A3(_11379_),
    .B1(_11413_),
    .X(_00652_));
 sky130_fd_sc_hd__nand2_1 _15727_ (.A(_11395_),
    .B(net4078),
    .Y(_11414_));
 sky130_fd_sc_hd__a22o_1 _15728_ (.A1(_11378_),
    .A2(_11414_),
    .B1(_11384_),
    .B2(_10331_),
    .X(_11415_));
 sky130_fd_sc_hd__inv_2 _15729_ (.A(_11415_),
    .Y(_00653_));
 sky130_fd_sc_hd__and3_1 _15730_ (.A(_11377_),
    .B(_10617_),
    .C(_11328_),
    .X(_11416_));
 sky130_fd_sc_hd__a31o_1 _15731_ (.A1(_11408_),
    .A2(net951),
    .A3(_11379_),
    .B1(_11416_),
    .X(_00654_));
 sky130_fd_sc_hd__nand2_1 _15732_ (.A(_11395_),
    .B(net3982),
    .Y(_11417_));
 sky130_fd_sc_hd__a22o_1 _15733_ (.A1(_11378_),
    .A2(_11417_),
    .B1(_11384_),
    .B2(_10335_),
    .X(_11418_));
 sky130_fd_sc_hd__inv_2 _15734_ (.A(_11418_),
    .Y(_00655_));
 sky130_fd_sc_hd__and3_1 _15735_ (.A(_11377_),
    .B(_10679_),
    .C(_11328_),
    .X(_11419_));
 sky130_fd_sc_hd__a31o_1 _15736_ (.A1(_11408_),
    .A2(net1069),
    .A3(_11380_),
    .B1(_11419_),
    .X(_00640_));
 sky130_fd_sc_hd__nor2_1 _15737_ (.A(_10681_),
    .B(_11380_),
    .Y(_11420_));
 sky130_fd_sc_hd__a31o_1 _15738_ (.A1(_11408_),
    .A2(net1279),
    .A3(_11380_),
    .B1(_11420_),
    .X(_00641_));
 sky130_fd_sc_hd__nand2_1 _15739_ (.A(_11395_),
    .B(net4217),
    .Y(_11421_));
 sky130_fd_sc_hd__a22o_1 _15740_ (.A1(_11378_),
    .A2(_11421_),
    .B1(_11384_),
    .B2(_09280_),
    .X(_11422_));
 sky130_fd_sc_hd__inv_2 _15741_ (.A(_11422_),
    .Y(_00642_));
 sky130_fd_sc_hd__nand2_1 _15742_ (.A(_11395_),
    .B(net3983),
    .Y(_11423_));
 sky130_fd_sc_hd__a22o_1 _15743_ (.A1(_11378_),
    .A2(_11423_),
    .B1(_11384_),
    .B2(_10342_),
    .X(_11424_));
 sky130_fd_sc_hd__inv_2 _15744_ (.A(_11424_),
    .Y(_00643_));
 sky130_fd_sc_hd__and3_1 _15745_ (.A(_11377_),
    .B(_10848_),
    .C(_11328_),
    .X(_11425_));
 sky130_fd_sc_hd__a31o_1 _15746_ (.A1(_11408_),
    .A2(net1885),
    .A3(_11380_),
    .B1(_11425_),
    .X(_00644_));
 sky130_fd_sc_hd__buf_8 _15747_ (.A(net78),
    .X(_11426_));
 sky130_fd_sc_hd__and3_1 _15748_ (.A(_11377_),
    .B(_11426_),
    .C(_11328_),
    .X(_11427_));
 sky130_fd_sc_hd__a31o_1 _15749_ (.A1(_11408_),
    .A2(net1637),
    .A3(_11380_),
    .B1(_11427_),
    .X(_00645_));
 sky130_fd_sc_hd__nand2_1 _15750_ (.A(_09196_),
    .B(net2675),
    .Y(_11428_));
 sky130_fd_sc_hd__a22oi_1 _15751_ (.A1(_11377_),
    .A2(_10348_),
    .B1(_11379_),
    .B2(_11428_),
    .Y(_00646_));
 sky130_fd_sc_hd__nor2_1 _15752_ (.A(_09300_),
    .B(_11380_),
    .Y(_11429_));
 sky130_fd_sc_hd__a31o_1 _15753_ (.A1(_11408_),
    .A2(net1505),
    .A3(_11380_),
    .B1(_11429_),
    .X(_00647_));
 sky130_fd_sc_hd__nor2_1 _15754_ (.A(_11376_),
    .B(_10292_),
    .Y(_11430_));
 sky130_fd_sc_hd__nand2_1 _15755_ (.A(_11430_),
    .B(_09359_),
    .Y(_11431_));
 sky130_fd_sc_hd__clkbuf_8 _15756_ (.A(_11431_),
    .X(_11432_));
 sky130_fd_sc_hd__nand2_1 _15757_ (.A(_11395_),
    .B(net4041),
    .Y(_11433_));
 sky130_fd_sc_hd__inv_2 _15758_ (.A(_11376_),
    .Y(_11434_));
 sky130_fd_sc_hd__and3_1 _15759_ (.A(_10291_),
    .B(_11434_),
    .C(_08725_),
    .X(_11435_));
 sky130_fd_sc_hd__clkbuf_8 _15760_ (.A(_11435_),
    .X(_11436_));
 sky130_fd_sc_hd__a22o_1 _15761_ (.A1(_11432_),
    .A2(_11433_),
    .B1(_09451_),
    .B2(_11436_),
    .X(_11437_));
 sky130_fd_sc_hd__inv_2 _15762_ (.A(_11437_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _15763_ (.A(_11395_),
    .B(net4091),
    .Y(_11438_));
 sky130_fd_sc_hd__buf_4 _15764_ (.A(_11436_),
    .X(_11439_));
 sky130_fd_sc_hd__a22o_1 _15765_ (.A1(_11432_),
    .A2(_11438_),
    .B1(_11439_),
    .B2(_09315_),
    .X(_11440_));
 sky130_fd_sc_hd__inv_2 _15766_ (.A(_11440_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _15767_ (.A(_11395_),
    .B(net4065),
    .Y(_11441_));
 sky130_fd_sc_hd__a22o_1 _15768_ (.A1(_11432_),
    .A2(_11441_),
    .B1(_11439_),
    .B2(_09460_),
    .X(_11442_));
 sky130_fd_sc_hd__inv_2 _15769_ (.A(_11442_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _15770_ (.A(_11395_),
    .B(net3967),
    .Y(_11443_));
 sky130_fd_sc_hd__a22o_1 _15771_ (.A1(_11432_),
    .A2(_11443_),
    .B1(_11439_),
    .B2(_09195_),
    .X(_11444_));
 sky130_fd_sc_hd__inv_2 _15772_ (.A(_11444_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _15773_ (.A(_11395_),
    .B(net4079),
    .Y(_11445_));
 sky130_fd_sc_hd__a22o_1 _15774_ (.A1(_11432_),
    .A2(_11445_),
    .B1(_11439_),
    .B2(_09201_),
    .X(_11446_));
 sky130_fd_sc_hd__inv_2 _15775_ (.A(_11446_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _15776_ (.A(_11395_),
    .B(net4225),
    .Y(_11447_));
 sky130_fd_sc_hd__a22o_1 _15777_ (.A1(_11432_),
    .A2(_11447_),
    .B1(_11439_),
    .B2(_09205_),
    .X(_11448_));
 sky130_fd_sc_hd__inv_2 _15778_ (.A(_11448_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _15779_ (.A(_11395_),
    .B(net4002),
    .Y(_11449_));
 sky130_fd_sc_hd__a22o_1 _15780_ (.A1(_11432_),
    .A2(_11449_),
    .B1(_11439_),
    .B2(_09398_),
    .X(_11450_));
 sky130_fd_sc_hd__inv_2 _15781_ (.A(_11450_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _15782_ (.A(_11395_),
    .B(net4200),
    .Y(_11451_));
 sky130_fd_sc_hd__a22o_1 _15783_ (.A1(_11432_),
    .A2(_11451_),
    .B1(_11439_),
    .B2(_09212_),
    .X(_11452_));
 sky130_fd_sc_hd__inv_2 _15784_ (.A(_11452_),
    .Y(_00639_));
 sky130_fd_sc_hd__buf_4 _15785_ (.A(_10930_),
    .X(_11453_));
 sky130_fd_sc_hd__nand2_1 _15786_ (.A(_11453_),
    .B(net4160),
    .Y(_11454_));
 sky130_fd_sc_hd__a22o_1 _15787_ (.A1(_11432_),
    .A2(_11454_),
    .B1(_11439_),
    .B2(_09531_),
    .X(_11455_));
 sky130_fd_sc_hd__inv_2 _15788_ (.A(_11455_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _15789_ (.A(_11453_),
    .B(net4021),
    .Y(_11456_));
 sky130_fd_sc_hd__a22o_1 _15790_ (.A1(_11432_),
    .A2(_11456_),
    .B1(_11439_),
    .B2(_10313_),
    .X(_11457_));
 sky130_fd_sc_hd__inv_2 _15791_ (.A(_11457_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _15792_ (.A(_11453_),
    .B(net3932),
    .Y(_11458_));
 sky130_fd_sc_hd__a22o_1 _15793_ (.A1(_11432_),
    .A2(_11458_),
    .B1(_11439_),
    .B2(_10316_),
    .X(_11459_));
 sky130_fd_sc_hd__inv_2 _15794_ (.A(_11459_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _15795_ (.A(_11453_),
    .B(net4013),
    .Y(_11460_));
 sky130_fd_sc_hd__a22o_1 _15796_ (.A1(_11432_),
    .A2(_11460_),
    .B1(_11439_),
    .B2(_09589_),
    .X(_11461_));
 sky130_fd_sc_hd__inv_2 _15797_ (.A(_11461_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _15798_ (.A(_11453_),
    .B(net3946),
    .Y(_11462_));
 sky130_fd_sc_hd__a22o_1 _15799_ (.A1(_11432_),
    .A2(_11462_),
    .B1(_11439_),
    .B2(_09593_),
    .X(_11463_));
 sky130_fd_sc_hd__inv_2 _15800_ (.A(_11463_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _15801_ (.A(_11453_),
    .B(net4259),
    .Y(_11464_));
 sky130_fd_sc_hd__a22o_1 _15802_ (.A1(_11432_),
    .A2(_11464_),
    .B1(_11439_),
    .B2(_09338_),
    .X(_11465_));
 sky130_fd_sc_hd__inv_2 _15803_ (.A(_11465_),
    .Y(_00629_));
 sky130_fd_sc_hd__buf_4 _15804_ (.A(_11431_),
    .X(_11466_));
 sky130_fd_sc_hd__nand2_1 _15805_ (.A(_11453_),
    .B(net3977),
    .Y(_11467_));
 sky130_fd_sc_hd__a22o_1 _15806_ (.A1(_11466_),
    .A2(_11467_),
    .B1(_11439_),
    .B2(_09239_),
    .X(_11468_));
 sky130_fd_sc_hd__inv_2 _15807_ (.A(_11468_),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _15808_ (.A(_11453_),
    .B(net4045),
    .Y(_11469_));
 sky130_fd_sc_hd__a22o_1 _15809_ (.A1(_11466_),
    .A2(_11469_),
    .B1(_11439_),
    .B2(_09768_),
    .X(_11470_));
 sky130_fd_sc_hd__inv_2 _15810_ (.A(_11470_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _15811_ (.A(_11453_),
    .B(net4228),
    .Y(_11471_));
 sky130_fd_sc_hd__a22o_1 _15812_ (.A1(_11466_),
    .A2(_11471_),
    .B1(_11439_),
    .B2(_09415_),
    .X(_11472_));
 sky130_fd_sc_hd__inv_2 _15813_ (.A(_11472_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _15814_ (.A(_11453_),
    .B(net4020),
    .Y(_11473_));
 sky130_fd_sc_hd__a22o_1 _15815_ (.A1(_11466_),
    .A2(_11473_),
    .B1(_11436_),
    .B2(_09249_),
    .X(_11474_));
 sky130_fd_sc_hd__inv_2 _15816_ (.A(_11474_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _15817_ (.A(_11453_),
    .B(net3993),
    .Y(_11475_));
 sky130_fd_sc_hd__a22o_1 _15818_ (.A1(_11466_),
    .A2(_11475_),
    .B1(_11436_),
    .B2(_09348_),
    .X(_11476_));
 sky130_fd_sc_hd__inv_2 _15819_ (.A(_11476_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _15820_ (.A(_11453_),
    .B(net3981),
    .Y(_11477_));
 sky130_fd_sc_hd__a22o_1 _15821_ (.A1(_11466_),
    .A2(_11477_),
    .B1(_11436_),
    .B2(_09256_),
    .X(_11478_));
 sky130_fd_sc_hd__inv_2 _15822_ (.A(_11478_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _15823_ (.A(_11453_),
    .B(net3877),
    .Y(_11479_));
 sky130_fd_sc_hd__a22o_1 _15824_ (.A1(_11466_),
    .A2(_11479_),
    .B1(_11436_),
    .B2(_09354_),
    .X(_11480_));
 sky130_fd_sc_hd__inv_2 _15825_ (.A(_11480_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _15826_ (.A(_11453_),
    .B(net3975),
    .Y(_11481_));
 sky130_fd_sc_hd__a22o_1 _15827_ (.A1(_11466_),
    .A2(_11481_),
    .B1(_11436_),
    .B2(_10331_),
    .X(_11482_));
 sky130_fd_sc_hd__inv_2 _15828_ (.A(_11482_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _15829_ (.A(_11453_),
    .B(net4139),
    .Y(_11483_));
 sky130_fd_sc_hd__a22o_1 _15830_ (.A1(_11466_),
    .A2(_11483_),
    .B1(_11436_),
    .B2(_09425_),
    .X(_11484_));
 sky130_fd_sc_hd__inv_2 _15831_ (.A(_11484_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _15832_ (.A(_11453_),
    .B(net3976),
    .Y(_11485_));
 sky130_fd_sc_hd__a22o_1 _15833_ (.A1(_11466_),
    .A2(_11485_),
    .B1(_11436_),
    .B2(_10335_),
    .X(_11486_));
 sky130_fd_sc_hd__inv_2 _15834_ (.A(_11486_),
    .Y(_00615_));
 sky130_fd_sc_hd__clkbuf_8 _15835_ (.A(_10930_),
    .X(_11487_));
 sky130_fd_sc_hd__nand2_1 _15836_ (.A(_11487_),
    .B(net3956),
    .Y(_11488_));
 sky130_fd_sc_hd__a22o_1 _15837_ (.A1(_11466_),
    .A2(_11488_),
    .B1(_11436_),
    .B2(_09495_),
    .X(_11489_));
 sky130_fd_sc_hd__inv_2 _15838_ (.A(_11489_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _15839_ (.A(_11487_),
    .B(net3945),
    .Y(_11490_));
 sky130_fd_sc_hd__a22o_1 _15840_ (.A1(_11466_),
    .A2(_11490_),
    .B1(_11436_),
    .B2(_09366_),
    .X(_11491_));
 sky130_fd_sc_hd__inv_2 _15841_ (.A(_11491_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _15842_ (.A(_11487_),
    .B(net4110),
    .Y(_11492_));
 sky130_fd_sc_hd__a22o_1 _15843_ (.A1(_11466_),
    .A2(_11492_),
    .B1(_11436_),
    .B2(_09280_),
    .X(_11493_));
 sky130_fd_sc_hd__inv_2 _15844_ (.A(_11493_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _15845_ (.A(_11487_),
    .B(net3968),
    .Y(_11494_));
 sky130_fd_sc_hd__a22o_1 _15846_ (.A1(_11466_),
    .A2(_11494_),
    .B1(_11436_),
    .B2(_10342_),
    .X(_11495_));
 sky130_fd_sc_hd__inv_2 _15847_ (.A(_11495_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _15848_ (.A(_11487_),
    .B(net4172),
    .Y(_11496_));
 sky130_fd_sc_hd__a22o_1 _15849_ (.A1(_11466_),
    .A2(_11496_),
    .B1(_11436_),
    .B2(_09288_),
    .X(_11497_));
 sky130_fd_sc_hd__inv_2 _15850_ (.A(_11497_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _15851_ (.A(_11487_),
    .B(net4092),
    .Y(_11498_));
 sky130_fd_sc_hd__a22o_1 _15852_ (.A1(_11466_),
    .A2(_11498_),
    .B1(_11436_),
    .B2(net136),
    .X(_11499_));
 sky130_fd_sc_hd__inv_2 _15853_ (.A(_11499_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _15854_ (.A(_11331_),
    .B(net4159),
    .Y(_11500_));
 sky130_fd_sc_hd__a22o_1 _15855_ (.A1(_10348_),
    .A2(_11430_),
    .B1(_11432_),
    .B2(_11500_),
    .X(_11501_));
 sky130_fd_sc_hd__inv_2 _15856_ (.A(_11501_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _15857_ (.A(_08777_),
    .B(net4252),
    .Y(_11502_));
 sky130_fd_sc_hd__a32o_1 _15858_ (.A1(_11436_),
    .A2(_08791_),
    .A3(_09299_),
    .B1(_11432_),
    .B2(_11502_),
    .X(_11503_));
 sky130_fd_sc_hd__inv_2 _15859_ (.A(net4253),
    .Y(_00607_));
 sky130_fd_sc_hd__nor2_4 _15860_ (.A(_11376_),
    .B(_10356_),
    .Y(_11504_));
 sky130_fd_sc_hd__nand2_4 _15861_ (.A(_11504_),
    .B(_09225_),
    .Y(_11505_));
 sky130_fd_sc_hd__buf_4 _15862_ (.A(_11505_),
    .X(_11506_));
 sky130_fd_sc_hd__buf_4 _15863_ (.A(_11505_),
    .X(_11507_));
 sky130_fd_sc_hd__nor2_1 _15864_ (.A(_11210_),
    .B(_11507_),
    .Y(_11508_));
 sky130_fd_sc_hd__a31o_1 _15865_ (.A1(_11408_),
    .A2(net1301),
    .A3(_11506_),
    .B1(_11508_),
    .X(_00592_));
 sky130_fd_sc_hd__nor2_1 _15866_ (.A(_10746_),
    .B(_11507_),
    .Y(_11509_));
 sky130_fd_sc_hd__a31o_1 _15867_ (.A1(_11408_),
    .A2(net1007),
    .A3(_11506_),
    .B1(_11509_),
    .X(_00593_));
 sky130_fd_sc_hd__nor2_1 _15868_ (.A(_10698_),
    .B(_11507_),
    .Y(_11510_));
 sky130_fd_sc_hd__a31o_1 _15869_ (.A1(_11408_),
    .A2(net1421),
    .A3(_11506_),
    .B1(_11510_),
    .X(_00594_));
 sky130_fd_sc_hd__nand2_1 _15870_ (.A(_11487_),
    .B(net4012),
    .Y(_11511_));
 sky130_fd_sc_hd__and3_1 _15871_ (.A(_10355_),
    .B(_11434_),
    .C(_08778_),
    .X(_11512_));
 sky130_fd_sc_hd__buf_4 _15872_ (.A(_11512_),
    .X(_11513_));
 sky130_fd_sc_hd__a22o_1 _15873_ (.A1(_11507_),
    .A2(_11511_),
    .B1(_11513_),
    .B2(_09195_),
    .X(_11514_));
 sky130_fd_sc_hd__inv_2 _15874_ (.A(_11514_),
    .Y(_00595_));
 sky130_fd_sc_hd__and3_1 _15875_ (.A(_11504_),
    .B(_10587_),
    .C(_11328_),
    .X(_11515_));
 sky130_fd_sc_hd__a31o_1 _15876_ (.A1(_11408_),
    .A2(net893),
    .A3(_11506_),
    .B1(_11515_),
    .X(_00596_));
 sky130_fd_sc_hd__buf_4 _15877_ (.A(_11219_),
    .X(_11516_));
 sky130_fd_sc_hd__and3_1 _15878_ (.A(_11504_),
    .B(_11391_),
    .C(_11516_),
    .X(_11517_));
 sky130_fd_sc_hd__a31o_1 _15879_ (.A1(_11408_),
    .A2(net715),
    .A3(_11506_),
    .B1(_11517_),
    .X(_00597_));
 sky130_fd_sc_hd__buf_4 _15880_ (.A(_10864_),
    .X(_11518_));
 sky130_fd_sc_hd__nor2_1 _15881_ (.A(_10872_),
    .B(_11507_),
    .Y(_11519_));
 sky130_fd_sc_hd__a31o_1 _15882_ (.A1(_11518_),
    .A2(net2057),
    .A3(_11506_),
    .B1(_11519_),
    .X(_00598_));
 sky130_fd_sc_hd__and3_1 _15883_ (.A(_11504_),
    .B(_10874_),
    .C(_11516_),
    .X(_11520_));
 sky130_fd_sc_hd__a31o_1 _15884_ (.A1(_11518_),
    .A2(net689),
    .A3(_11506_),
    .B1(_11520_),
    .X(_00599_));
 sky130_fd_sc_hd__nand2_1 _15885_ (.A(_11487_),
    .B(net4011),
    .Y(_11521_));
 sky130_fd_sc_hd__a22o_1 _15886_ (.A1(_11507_),
    .A2(_11521_),
    .B1(_11513_),
    .B2(_09531_),
    .X(_11522_));
 sky130_fd_sc_hd__inv_2 _15887_ (.A(_11522_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _15888_ (.A(_11487_),
    .B(net4049),
    .Y(_11523_));
 sky130_fd_sc_hd__a22o_1 _15889_ (.A1(_11507_),
    .A2(_11523_),
    .B1(_11513_),
    .B2(_10313_),
    .X(_11524_));
 sky130_fd_sc_hd__inv_2 _15890_ (.A(_11524_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_1 _15891_ (.A(_11487_),
    .B(net4103),
    .Y(_11525_));
 sky130_fd_sc_hd__a22o_1 _15892_ (.A1(_11507_),
    .A2(_11525_),
    .B1(_11513_),
    .B2(_10316_),
    .X(_11526_));
 sky130_fd_sc_hd__inv_2 _15893_ (.A(_11526_),
    .Y(_00586_));
 sky130_fd_sc_hd__nor2_1 _15894_ (.A(_10657_),
    .B(_11507_),
    .Y(_11527_));
 sky130_fd_sc_hd__a31o_1 _15895_ (.A1(_11518_),
    .A2(net903),
    .A3(_11506_),
    .B1(_11527_),
    .X(_00587_));
 sky130_fd_sc_hd__nand2_1 _15896_ (.A(_11487_),
    .B(net4034),
    .Y(_11528_));
 sky130_fd_sc_hd__a22o_1 _15897_ (.A1(_11505_),
    .A2(_11528_),
    .B1(_11513_),
    .B2(_09593_),
    .X(_11529_));
 sky130_fd_sc_hd__inv_2 _15898_ (.A(_11529_),
    .Y(_00588_));
 sky130_fd_sc_hd__nor2_1 _15899_ (.A(_10602_),
    .B(_11507_),
    .Y(_11530_));
 sky130_fd_sc_hd__a31o_1 _15900_ (.A1(_11518_),
    .A2(net1127),
    .A3(_11506_),
    .B1(_11530_),
    .X(_00589_));
 sky130_fd_sc_hd__nand2_1 _15901_ (.A(_11487_),
    .B(net4077),
    .Y(_11531_));
 sky130_fd_sc_hd__a22o_1 _15902_ (.A1(_11505_),
    .A2(_11531_),
    .B1(_11513_),
    .B2(_09239_),
    .X(_11532_));
 sky130_fd_sc_hd__inv_2 _15903_ (.A(_11532_),
    .Y(_00590_));
 sky130_fd_sc_hd__nor2_1 _15904_ (.A(_10663_),
    .B(_11507_),
    .Y(_11533_));
 sky130_fd_sc_hd__a31o_1 _15905_ (.A1(_11518_),
    .A2(net721),
    .A3(_11506_),
    .B1(_11533_),
    .X(_00591_));
 sky130_fd_sc_hd__nand2_1 _15906_ (.A(_11487_),
    .B(net4095),
    .Y(_11534_));
 sky130_fd_sc_hd__a22o_1 _15907_ (.A1(_11505_),
    .A2(_11534_),
    .B1(_11513_),
    .B2(_09415_),
    .X(_11535_));
 sky130_fd_sc_hd__inv_2 _15908_ (.A(_11535_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _15909_ (.A(_11487_),
    .B(net4035),
    .Y(_11536_));
 sky130_fd_sc_hd__a22o_1 _15910_ (.A1(_11505_),
    .A2(_11536_),
    .B1(_11513_),
    .B2(_09249_),
    .X(_11537_));
 sky130_fd_sc_hd__inv_2 _15911_ (.A(_11537_),
    .Y(_00577_));
 sky130_fd_sc_hd__nor2_1 _15912_ (.A(_10669_),
    .B(_11507_),
    .Y(_11538_));
 sky130_fd_sc_hd__a31o_1 _15913_ (.A1(_11518_),
    .A2(net1189),
    .A3(_11506_),
    .B1(_11538_),
    .X(_00578_));
 sky130_fd_sc_hd__and3_1 _15914_ (.A(_11504_),
    .B(_10500_),
    .C(_11516_),
    .X(_11539_));
 sky130_fd_sc_hd__a31o_1 _15915_ (.A1(_11518_),
    .A2(net921),
    .A3(_11506_),
    .B1(_11539_),
    .X(_00579_));
 sky130_fd_sc_hd__nor2_1 _15916_ (.A(_11010_),
    .B(_11507_),
    .Y(_11540_));
 sky130_fd_sc_hd__a31o_1 _15917_ (.A1(_11518_),
    .A2(net1231),
    .A3(_11506_),
    .B1(_11540_),
    .X(_00580_));
 sky130_fd_sc_hd__nand2_1 _15918_ (.A(_11487_),
    .B(net4174),
    .Y(_11541_));
 sky130_fd_sc_hd__a22o_1 _15919_ (.A1(_11505_),
    .A2(_11541_),
    .B1(_11513_),
    .B2(_10331_),
    .X(_11542_));
 sky130_fd_sc_hd__inv_2 _15920_ (.A(_11542_),
    .Y(_00581_));
 sky130_fd_sc_hd__and3_1 _15921_ (.A(_11504_),
    .B(_10617_),
    .C(_11516_),
    .X(_11543_));
 sky130_fd_sc_hd__a31o_1 _15922_ (.A1(_11518_),
    .A2(net2075),
    .A3(_11506_),
    .B1(_11543_),
    .X(_00582_));
 sky130_fd_sc_hd__nand2_1 _15923_ (.A(_11487_),
    .B(net4241),
    .Y(_11544_));
 sky130_fd_sc_hd__a22o_1 _15924_ (.A1(_11505_),
    .A2(_11544_),
    .B1(_11513_),
    .B2(_10335_),
    .X(_11545_));
 sky130_fd_sc_hd__inv_2 _15925_ (.A(_11545_),
    .Y(_00583_));
 sky130_fd_sc_hd__and3_1 _15926_ (.A(_11504_),
    .B(_10679_),
    .C(_11516_),
    .X(_11546_));
 sky130_fd_sc_hd__a31o_1 _15927_ (.A1(_11518_),
    .A2(net1427),
    .A3(_11506_),
    .B1(_11546_),
    .X(_00568_));
 sky130_fd_sc_hd__buf_4 _15928_ (.A(_10930_),
    .X(_11547_));
 sky130_fd_sc_hd__nand2_1 _15929_ (.A(_11547_),
    .B(net4043),
    .Y(_11548_));
 sky130_fd_sc_hd__a22o_1 _15930_ (.A1(_11505_),
    .A2(_11548_),
    .B1(_11513_),
    .B2(_09366_),
    .X(_11549_));
 sky130_fd_sc_hd__inv_2 _15931_ (.A(_11549_),
    .Y(_00569_));
 sky130_fd_sc_hd__and3_1 _15932_ (.A(_11504_),
    .B(_10728_),
    .C(_11516_),
    .X(_11550_));
 sky130_fd_sc_hd__a31o_1 _15933_ (.A1(_11518_),
    .A2(net1157),
    .A3(_11506_),
    .B1(_11550_),
    .X(_00570_));
 sky130_fd_sc_hd__nand2_1 _15934_ (.A(_11547_),
    .B(net4138),
    .Y(_11551_));
 sky130_fd_sc_hd__a22o_1 _15935_ (.A1(_11505_),
    .A2(_11551_),
    .B1(_11513_),
    .B2(_10342_),
    .X(_11552_));
 sky130_fd_sc_hd__inv_2 _15936_ (.A(_11552_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _15937_ (.A(_11547_),
    .B(net4141),
    .Y(_11553_));
 sky130_fd_sc_hd__a22o_1 _15938_ (.A1(_11505_),
    .A2(_11553_),
    .B1(_11513_),
    .B2(_09288_),
    .X(_11554_));
 sky130_fd_sc_hd__inv_2 _15939_ (.A(_11554_),
    .Y(_00572_));
 sky130_fd_sc_hd__and3_1 _15940_ (.A(_11504_),
    .B(_11426_),
    .C(_11516_),
    .X(_11555_));
 sky130_fd_sc_hd__a31o_1 _15941_ (.A1(_11518_),
    .A2(net711),
    .A3(_11507_),
    .B1(_11555_),
    .X(_00573_));
 sky130_fd_sc_hd__buf_4 _15942_ (.A(_11151_),
    .X(_11556_));
 sky130_fd_sc_hd__nand2_1 _15943_ (.A(_11556_),
    .B(net3568),
    .Y(_11557_));
 sky130_fd_sc_hd__a22o_1 _15944_ (.A1(_10348_),
    .A2(_11504_),
    .B1(_11507_),
    .B2(_11557_),
    .X(_11558_));
 sky130_fd_sc_hd__inv_2 _15945_ (.A(net3569),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(_11556_),
    .B(net2990),
    .Y(_11559_));
 sky130_fd_sc_hd__a22o_1 _15947_ (.A1(_09440_),
    .A2(_11504_),
    .B1(_11507_),
    .B2(_11559_),
    .X(_11560_));
 sky130_fd_sc_hd__inv_2 _15948_ (.A(net2991),
    .Y(_00575_));
 sky130_fd_sc_hd__nor2_2 _15949_ (.A(_11376_),
    .B(_10411_),
    .Y(_11561_));
 sky130_fd_sc_hd__inv_2 _15950_ (.A(_11561_),
    .Y(_11562_));
 sky130_fd_sc_hd__nor2_1 _15951_ (.A(_08797_),
    .B(_11562_),
    .Y(_11563_));
 sky130_fd_sc_hd__buf_4 _15952_ (.A(_11563_),
    .X(_11564_));
 sky130_fd_sc_hd__nor2_1 _15953_ (.A(_08728_),
    .B(_11562_),
    .Y(_11565_));
 sky130_fd_sc_hd__inv_2 _15954_ (.A(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__buf_4 _15955_ (.A(_11566_),
    .X(_11567_));
 sky130_fd_sc_hd__nand2_1 _15956_ (.A(_11556_),
    .B(net3447),
    .Y(_11568_));
 sky130_fd_sc_hd__a22o_1 _15957_ (.A1(_11564_),
    .A2(_10239_),
    .B1(_11567_),
    .B2(_11568_),
    .X(_11569_));
 sky130_fd_sc_hd__inv_2 _15958_ (.A(_11569_),
    .Y(_00560_));
 sky130_fd_sc_hd__buf_4 _15959_ (.A(_11566_),
    .X(_11570_));
 sky130_fd_sc_hd__nor2_1 _15960_ (.A(_10746_),
    .B(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__a31o_1 _15961_ (.A1(_11518_),
    .A2(net2133),
    .A3(_11570_),
    .B1(_11571_),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_1 _15962_ (.A(_11556_),
    .B(net3730),
    .Y(_11572_));
 sky130_fd_sc_hd__a22o_1 _15963_ (.A1(_11564_),
    .A2(_09459_),
    .B1(_11567_),
    .B2(_11572_),
    .X(_11573_));
 sky130_fd_sc_hd__inv_2 _15964_ (.A(_11573_),
    .Y(_00562_));
 sky130_fd_sc_hd__nand2_1 _15965_ (.A(_11556_),
    .B(net3238),
    .Y(_11574_));
 sky130_fd_sc_hd__a22o_1 _15966_ (.A1(_11564_),
    .A2(_10983_),
    .B1(_11567_),
    .B2(_11574_),
    .X(_11575_));
 sky130_fd_sc_hd__inv_2 _15967_ (.A(_11575_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _15968_ (.A(_11556_),
    .B(net3463),
    .Y(_11576_));
 sky130_fd_sc_hd__a22o_1 _15969_ (.A1(_11564_),
    .A2(_11330_),
    .B1(_11567_),
    .B2(_11576_),
    .X(_11577_));
 sky130_fd_sc_hd__inv_2 _15970_ (.A(_11577_),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_1 _15971_ (.A(_11556_),
    .B(net3475),
    .Y(_11578_));
 sky130_fd_sc_hd__a22o_1 _15972_ (.A1(_11564_),
    .A2(_10869_),
    .B1(_11567_),
    .B2(_11578_),
    .X(_11579_));
 sky130_fd_sc_hd__inv_2 _15973_ (.A(_11579_),
    .Y(_00565_));
 sky130_fd_sc_hd__nor2_1 _15974_ (.A(_10872_),
    .B(_11567_),
    .Y(_11580_));
 sky130_fd_sc_hd__a31o_1 _15975_ (.A1(_11518_),
    .A2(net1105),
    .A3(_11570_),
    .B1(_11580_),
    .X(_00566_));
 sky130_fd_sc_hd__and3_1 _15976_ (.A(_11561_),
    .B(_10874_),
    .C(_11516_),
    .X(_11581_));
 sky130_fd_sc_hd__a31o_1 _15977_ (.A1(_11570_),
    .A2(_11311_),
    .A3(net2164),
    .B1(_11581_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _15978_ (.A(_10760_),
    .B(_11567_),
    .Y(_11582_));
 sky130_fd_sc_hd__a31o_1 _15979_ (.A1(_11518_),
    .A2(net411),
    .A3(_11570_),
    .B1(_11582_),
    .X(_00552_));
 sky130_fd_sc_hd__nand2_1 _15980_ (.A(_11556_),
    .B(net3346),
    .Y(_11583_));
 sky130_fd_sc_hd__a22o_1 _15981_ (.A1(_11564_),
    .A2(_10122_),
    .B1(_11567_),
    .B2(_11583_),
    .X(_11584_));
 sky130_fd_sc_hd__inv_2 _15982_ (.A(_11584_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_1 _15983_ (.A(_11556_),
    .B(net3261),
    .Y(_11585_));
 sky130_fd_sc_hd__a22o_1 _15984_ (.A1(_11564_),
    .A2(_10195_),
    .B1(_11567_),
    .B2(_11585_),
    .X(_11586_));
 sky130_fd_sc_hd__inv_2 _15985_ (.A(_11586_),
    .Y(_00554_));
 sky130_fd_sc_hd__nor2_1 _15986_ (.A(_10657_),
    .B(_11567_),
    .Y(_11587_));
 sky130_fd_sc_hd__a31o_1 _15987_ (.A1(_11518_),
    .A2(net1593),
    .A3(_11570_),
    .B1(_11587_),
    .X(_00555_));
 sky130_fd_sc_hd__buf_4 _15988_ (.A(_10864_),
    .X(_11588_));
 sky130_fd_sc_hd__nor2_1 _15989_ (.A(_10767_),
    .B(_11567_),
    .Y(_11589_));
 sky130_fd_sc_hd__a31o_1 _15990_ (.A1(_11588_),
    .A2(net1213),
    .A3(_11570_),
    .B1(_11589_),
    .X(_00556_));
 sky130_fd_sc_hd__nor2_1 _15991_ (.A(_10602_),
    .B(_11567_),
    .Y(_11590_));
 sky130_fd_sc_hd__a31o_1 _15992_ (.A1(_11588_),
    .A2(net1821),
    .A3(_11570_),
    .B1(_11590_),
    .X(_00557_));
 sky130_fd_sc_hd__nand2_1 _15993_ (.A(_11556_),
    .B(net3875),
    .Y(_11591_));
 sky130_fd_sc_hd__a22o_1 _15994_ (.A1(_11564_),
    .A2(_10202_),
    .B1(_11567_),
    .B2(_11591_),
    .X(_11592_));
 sky130_fd_sc_hd__inv_2 _15995_ (.A(_11592_),
    .Y(_00558_));
 sky130_fd_sc_hd__nor2_1 _15996_ (.A(_10663_),
    .B(_11567_),
    .Y(_11593_));
 sky130_fd_sc_hd__a31o_1 _15997_ (.A1(_11588_),
    .A2(net891),
    .A3(_11570_),
    .B1(_11593_),
    .X(_00559_));
 sky130_fd_sc_hd__nand2_1 _15998_ (.A(_11556_),
    .B(net3013),
    .Y(_11594_));
 sky130_fd_sc_hd__a22o_1 _15999_ (.A1(_11564_),
    .A2(net137),
    .B1(_11567_),
    .B2(_11594_),
    .X(_11595_));
 sky130_fd_sc_hd__inv_2 _16000_ (.A(_11595_),
    .Y(_00544_));
 sky130_fd_sc_hd__and3_1 _16001_ (.A(_11561_),
    .B(_10667_),
    .C(_11516_),
    .X(_11596_));
 sky130_fd_sc_hd__a31o_1 _16002_ (.A1(_11570_),
    .A2(_11311_),
    .A3(net2266),
    .B1(_11596_),
    .X(_00545_));
 sky130_fd_sc_hd__nand2_1 _16003_ (.A(_11556_),
    .B(net3556),
    .Y(_11597_));
 sky130_fd_sc_hd__a22o_1 _16004_ (.A1(_11564_),
    .A2(_09347_),
    .B1(_11566_),
    .B2(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__inv_2 _16005_ (.A(_11598_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _16006_ (.A(_11556_),
    .B(net3116),
    .Y(_11599_));
 sky130_fd_sc_hd__a22o_1 _16007_ (.A1(_11564_),
    .A2(_09256_),
    .B1(_11566_),
    .B2(_11599_),
    .X(_11600_));
 sky130_fd_sc_hd__inv_2 _16008_ (.A(_11600_),
    .Y(_00547_));
 sky130_fd_sc_hd__nor2_1 _16009_ (.A(_11010_),
    .B(_11567_),
    .Y(_11601_));
 sky130_fd_sc_hd__a31o_1 _16010_ (.A1(_11588_),
    .A2(net731),
    .A3(_11570_),
    .B1(_11601_),
    .X(_00548_));
 sky130_fd_sc_hd__nand2_1 _16011_ (.A(_11556_),
    .B(net3445),
    .Y(_11602_));
 sky130_fd_sc_hd__a22o_1 _16012_ (.A1(_11564_),
    .A2(_10149_),
    .B1(_11566_),
    .B2(_11602_),
    .X(_11603_));
 sky130_fd_sc_hd__inv_2 _16013_ (.A(_11603_),
    .Y(_00549_));
 sky130_fd_sc_hd__and3_1 _16014_ (.A(_11561_),
    .B(_10617_),
    .C(_11516_),
    .X(_11604_));
 sky130_fd_sc_hd__a31o_1 _16015_ (.A1(_11570_),
    .A2(_11311_),
    .A3(net1894),
    .B1(_11604_),
    .X(_00550_));
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(_11556_),
    .B(net3845),
    .Y(_11605_));
 sky130_fd_sc_hd__a22o_1 _16017_ (.A1(_11564_),
    .A2(_10154_),
    .B1(_11566_),
    .B2(_11605_),
    .X(_11606_));
 sky130_fd_sc_hd__inv_2 _16018_ (.A(_11606_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _16019_ (.A(_11556_),
    .B(net3395),
    .Y(_11607_));
 sky130_fd_sc_hd__a22o_1 _16020_ (.A1(_11564_),
    .A2(net141),
    .B1(_11566_),
    .B2(_11607_),
    .X(_11608_));
 sky130_fd_sc_hd__inv_2 _16021_ (.A(_11608_),
    .Y(_00536_));
 sky130_fd_sc_hd__buf_4 _16022_ (.A(_11151_),
    .X(_11609_));
 sky130_fd_sc_hd__nand2_1 _16023_ (.A(_11609_),
    .B(net3954),
    .Y(_11610_));
 sky130_fd_sc_hd__a22o_1 _16024_ (.A1(_11564_),
    .A2(_09365_),
    .B1(_11566_),
    .B2(_11610_),
    .X(_11611_));
 sky130_fd_sc_hd__inv_2 _16025_ (.A(_11611_),
    .Y(_00537_));
 sky130_fd_sc_hd__and3_1 _16026_ (.A(_11561_),
    .B(_10728_),
    .C(_11516_),
    .X(_11612_));
 sky130_fd_sc_hd__a31o_1 _16027_ (.A1(_11570_),
    .A2(_11311_),
    .A3(net1983),
    .B1(_11612_),
    .X(_00538_));
 sky130_fd_sc_hd__nand2_1 _16028_ (.A(_11609_),
    .B(net3634),
    .Y(_11613_));
 sky130_fd_sc_hd__a22o_1 _16029_ (.A1(_11564_),
    .A2(_10164_),
    .B1(_11566_),
    .B2(_11613_),
    .X(_11614_));
 sky130_fd_sc_hd__inv_2 _16030_ (.A(_11614_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand2_1 _16031_ (.A(_11609_),
    .B(net3856),
    .Y(_11615_));
 sky130_fd_sc_hd__a22o_1 _16032_ (.A1(_11563_),
    .A2(net139),
    .B1(_11566_),
    .B2(_11615_),
    .X(_11616_));
 sky130_fd_sc_hd__inv_2 _16033_ (.A(_11616_),
    .Y(_00540_));
 sky130_fd_sc_hd__and3_1 _16034_ (.A(_11561_),
    .B(_11426_),
    .C(_11516_),
    .X(_11617_));
 sky130_fd_sc_hd__a31o_1 _16035_ (.A1(_11570_),
    .A2(_11311_),
    .A3(net2064),
    .B1(_11617_),
    .X(_00541_));
 sky130_fd_sc_hd__nand2_1 _16036_ (.A(_11174_),
    .B(net4038),
    .Y(_11618_));
 sky130_fd_sc_hd__o2bb2a_1 _16037_ (.A1_N(_11618_),
    .A2_N(_11570_),
    .B1(_10289_),
    .B2(_11562_),
    .X(_00542_));
 sky130_fd_sc_hd__nand2_1 _16038_ (.A(_11174_),
    .B(net4070),
    .Y(_11619_));
 sky130_fd_sc_hd__o2bb2a_1 _16039_ (.A1_N(_11619_),
    .A2_N(_11570_),
    .B1(_11316_),
    .B2(_11562_),
    .X(_00543_));
 sky130_fd_sc_hd__nand2_8 _16040_ (.A(_09735_),
    .B(_11161_),
    .Y(_11620_));
 sky130_fd_sc_hd__nor2_2 _16041_ (.A(_10469_),
    .B(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__inv_2 _16042_ (.A(_11621_),
    .Y(_11622_));
 sky130_fd_sc_hd__nor2_1 _16043_ (.A(_08727_),
    .B(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__clkinv_4 _16044_ (.A(_11623_),
    .Y(_11624_));
 sky130_fd_sc_hd__buf_4 _16045_ (.A(_11624_),
    .X(_11625_));
 sky130_fd_sc_hd__buf_4 _16046_ (.A(_11624_),
    .X(_11626_));
 sky130_fd_sc_hd__nor2_1 _16047_ (.A(_11210_),
    .B(_11626_),
    .Y(_11627_));
 sky130_fd_sc_hd__a31o_1 _16048_ (.A1(_11588_),
    .A2(net2445),
    .A3(_11625_),
    .B1(_11627_),
    .X(_00520_));
 sky130_fd_sc_hd__nor2_1 _16049_ (.A(_10746_),
    .B(_11626_),
    .Y(_11628_));
 sky130_fd_sc_hd__a31o_1 _16050_ (.A1(_11588_),
    .A2(net589),
    .A3(_11625_),
    .B1(_11628_),
    .X(_00521_));
 sky130_fd_sc_hd__nor2_1 _16051_ (.A(_10698_),
    .B(_11626_),
    .Y(_11629_));
 sky130_fd_sc_hd__a31o_1 _16052_ (.A1(_11588_),
    .A2(net889),
    .A3(_11625_),
    .B1(_11629_),
    .X(_00522_));
 sky130_fd_sc_hd__and3_1 _16053_ (.A(_11621_),
    .B(_11040_),
    .C(_11516_),
    .X(_11630_));
 sky130_fd_sc_hd__a31o_1 _16054_ (.A1(_11625_),
    .A2(_11311_),
    .A3(net2353),
    .B1(_11630_),
    .X(_00523_));
 sky130_fd_sc_hd__and3_1 _16055_ (.A(_11621_),
    .B(_10587_),
    .C(_11516_),
    .X(_11631_));
 sky130_fd_sc_hd__a31o_1 _16056_ (.A1(_11625_),
    .A2(_11311_),
    .A3(net2309),
    .B1(_11631_),
    .X(_00524_));
 sky130_fd_sc_hd__nor2_4 _16057_ (.A(_09190_),
    .B(_11622_),
    .Y(_11632_));
 sky130_fd_sc_hd__nand2_1 _16058_ (.A(_11609_),
    .B(net3498),
    .Y(_11633_));
 sky130_fd_sc_hd__a22o_1 _16059_ (.A1(_11632_),
    .A2(_10869_),
    .B1(_11626_),
    .B2(_11633_),
    .X(_11634_));
 sky130_fd_sc_hd__inv_2 _16060_ (.A(_11634_),
    .Y(_00525_));
 sky130_fd_sc_hd__nor2_1 _16061_ (.A(_10872_),
    .B(_11626_),
    .Y(_11635_));
 sky130_fd_sc_hd__a31o_1 _16062_ (.A1(_11588_),
    .A2(net1299),
    .A3(_11625_),
    .B1(_11635_),
    .X(_00526_));
 sky130_fd_sc_hd__nand2_1 _16063_ (.A(_11609_),
    .B(net3685),
    .Y(_11636_));
 sky130_fd_sc_hd__a22o_1 _16064_ (.A1(_11632_),
    .A2(_10591_),
    .B1(_11624_),
    .B2(_11636_),
    .X(_11637_));
 sky130_fd_sc_hd__inv_2 _16065_ (.A(_11637_),
    .Y(_00527_));
 sky130_fd_sc_hd__nor2_1 _16066_ (.A(_10760_),
    .B(_11626_),
    .Y(_11638_));
 sky130_fd_sc_hd__a31o_1 _16067_ (.A1(_11588_),
    .A2(net1855),
    .A3(_11625_),
    .B1(_11638_),
    .X(_00512_));
 sky130_fd_sc_hd__nand2_1 _16068_ (.A(_11609_),
    .B(net3492),
    .Y(_11639_));
 sky130_fd_sc_hd__a22o_1 _16069_ (.A1(_11632_),
    .A2(_10122_),
    .B1(_11624_),
    .B2(_11639_),
    .X(_11640_));
 sky130_fd_sc_hd__inv_2 _16070_ (.A(_11640_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(_11609_),
    .B(net3586),
    .Y(_11641_));
 sky130_fd_sc_hd__a22o_1 _16072_ (.A1(_11632_),
    .A2(_10195_),
    .B1(_11624_),
    .B2(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__inv_2 _16073_ (.A(_11642_),
    .Y(_00514_));
 sky130_fd_sc_hd__nor2_1 _16074_ (.A(_10657_),
    .B(_11626_),
    .Y(_11643_));
 sky130_fd_sc_hd__a31o_1 _16075_ (.A1(_11588_),
    .A2(net1951),
    .A3(_11625_),
    .B1(_11643_),
    .X(_00515_));
 sky130_fd_sc_hd__nor2_1 _16076_ (.A(_10767_),
    .B(_11626_),
    .Y(_02733_));
 sky130_fd_sc_hd__a31o_1 _16077_ (.A1(_11588_),
    .A2(net1941),
    .A3(_11625_),
    .B1(_02733_),
    .X(_00516_));
 sky130_fd_sc_hd__nor2_1 _16078_ (.A(_10602_),
    .B(_11626_),
    .Y(_02734_));
 sky130_fd_sc_hd__a31o_1 _16079_ (.A1(_11588_),
    .A2(net933),
    .A3(_11625_),
    .B1(_02734_),
    .X(_00517_));
 sky130_fd_sc_hd__and3_1 _16080_ (.A(_11621_),
    .B(_11291_),
    .C(_11516_),
    .X(_02735_));
 sky130_fd_sc_hd__a31o_1 _16081_ (.A1(_11625_),
    .A2(_11311_),
    .A3(net2128),
    .B1(_02735_),
    .X(_00518_));
 sky130_fd_sc_hd__nor2_1 _16082_ (.A(_10663_),
    .B(_11626_),
    .Y(_02736_));
 sky130_fd_sc_hd__a31o_1 _16083_ (.A1(_11588_),
    .A2(net965),
    .A3(_11625_),
    .B1(_02736_),
    .X(_00519_));
 sky130_fd_sc_hd__nor2_1 _16084_ (.A(_11002_),
    .B(_11626_),
    .Y(_02737_));
 sky130_fd_sc_hd__a31o_1 _16085_ (.A1(_11588_),
    .A2(net1529),
    .A3(_11626_),
    .B1(_02737_),
    .X(_00504_));
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(_11609_),
    .B(net3458),
    .Y(_02738_));
 sky130_fd_sc_hd__a22o_1 _16087_ (.A1(_11632_),
    .A2(_09249_),
    .B1(_11624_),
    .B2(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__inv_2 _16088_ (.A(_02739_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _16089_ (.A(_11609_),
    .B(net2936),
    .Y(_02740_));
 sky130_fd_sc_hd__a22o_1 _16090_ (.A1(_11632_),
    .A2(_09347_),
    .B1(_11624_),
    .B2(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__inv_2 _16091_ (.A(_02741_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _16092_ (.A(_11609_),
    .B(net3382),
    .Y(_02742_));
 sky130_fd_sc_hd__a22o_1 _16093_ (.A1(_11632_),
    .A2(_09256_),
    .B1(_11624_),
    .B2(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__inv_2 _16094_ (.A(_02743_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _16095_ (.A(_11609_),
    .B(net3531),
    .Y(_02744_));
 sky130_fd_sc_hd__a22o_1 _16096_ (.A1(_11632_),
    .A2(_11136_),
    .B1(_11624_),
    .B2(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__inv_2 _16097_ (.A(_02745_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _16098_ (.A(_11609_),
    .B(net3332),
    .Y(_02746_));
 sky130_fd_sc_hd__a22o_1 _16099_ (.A1(_11632_),
    .A2(_10149_),
    .B1(_11624_),
    .B2(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__inv_2 _16100_ (.A(_02747_),
    .Y(_00509_));
 sky130_fd_sc_hd__and3_1 _16101_ (.A(_11621_),
    .B(_10617_),
    .C(_11516_),
    .X(_02748_));
 sky130_fd_sc_hd__a31o_1 _16102_ (.A1(_11625_),
    .A2(_11311_),
    .A3(net2274),
    .B1(_02748_),
    .X(_00510_));
 sky130_fd_sc_hd__nand2_1 _16103_ (.A(_11609_),
    .B(net3780),
    .Y(_02749_));
 sky130_fd_sc_hd__a22o_1 _16104_ (.A1(_11632_),
    .A2(_10154_),
    .B1(_11624_),
    .B2(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__inv_2 _16105_ (.A(_02750_),
    .Y(_00511_));
 sky130_fd_sc_hd__clkbuf_8 _16106_ (.A(_10645_),
    .X(_02751_));
 sky130_fd_sc_hd__clkbuf_4 _16107_ (.A(_11219_),
    .X(_02752_));
 sky130_fd_sc_hd__and3_1 _16108_ (.A(_11621_),
    .B(_10679_),
    .C(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__a31o_1 _16109_ (.A1(_11625_),
    .A2(_02751_),
    .A3(net2169),
    .B1(_02753_),
    .X(_00496_));
 sky130_fd_sc_hd__nor2_1 _16110_ (.A(_10681_),
    .B(_11626_),
    .Y(_02754_));
 sky130_fd_sc_hd__a31o_1 _16111_ (.A1(_11588_),
    .A2(net585),
    .A3(_11626_),
    .B1(_02754_),
    .X(_00497_));
 sky130_fd_sc_hd__nand2_1 _16112_ (.A(_11609_),
    .B(net3390),
    .Y(_02755_));
 sky130_fd_sc_hd__a22o_1 _16113_ (.A1(_11632_),
    .A2(_10624_),
    .B1(_11624_),
    .B2(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__inv_2 _16114_ (.A(_02756_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _16115_ (.A(_11609_),
    .B(net3467),
    .Y(_02757_));
 sky130_fd_sc_hd__a22o_1 _16116_ (.A1(_11632_),
    .A2(_10164_),
    .B1(_11624_),
    .B2(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__inv_2 _16117_ (.A(_02758_),
    .Y(_00499_));
 sky130_fd_sc_hd__and3_1 _16118_ (.A(_11621_),
    .B(_10848_),
    .C(_02752_),
    .X(_02759_));
 sky130_fd_sc_hd__a31o_1 _16119_ (.A1(_11625_),
    .A2(_02751_),
    .A3(net2320),
    .B1(_02759_),
    .X(_00500_));
 sky130_fd_sc_hd__nand2_1 _16120_ (.A(_11609_),
    .B(net3590),
    .Y(_02760_));
 sky130_fd_sc_hd__a22o_1 _16121_ (.A1(_11632_),
    .A2(net136),
    .B1(_11624_),
    .B2(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__inv_2 _16122_ (.A(_02761_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _16123_ (.A(_11174_),
    .B(net3839),
    .Y(_02762_));
 sky130_fd_sc_hd__o2bb2a_1 _16124_ (.A1_N(_02762_),
    .A2_N(_11625_),
    .B1(_10289_),
    .B2(_11622_),
    .X(_00502_));
 sky130_fd_sc_hd__nor2_1 _16125_ (.A(_09300_),
    .B(_11626_),
    .Y(_02763_));
 sky130_fd_sc_hd__a31o_1 _16126_ (.A1(_11588_),
    .A2(net687),
    .A3(_11626_),
    .B1(_02763_),
    .X(_00503_));
 sky130_fd_sc_hd__nor2_4 _16127_ (.A(_11620_),
    .B(_10292_),
    .Y(_02764_));
 sky130_fd_sc_hd__nand2_4 _16128_ (.A(_02764_),
    .B(_10413_),
    .Y(_02765_));
 sky130_fd_sc_hd__buf_4 _16129_ (.A(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__nand2_1 _16130_ (.A(_11547_),
    .B(net4101),
    .Y(_02767_));
 sky130_fd_sc_hd__inv_2 _16131_ (.A(_11620_),
    .Y(_02768_));
 sky130_fd_sc_hd__and3_1 _16132_ (.A(_10291_),
    .B(_02768_),
    .C(_08725_),
    .X(_02769_));
 sky130_fd_sc_hd__buf_4 _16133_ (.A(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__a22o_1 _16134_ (.A1(_02766_),
    .A2(_02767_),
    .B1(_09451_),
    .B2(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__inv_2 _16135_ (.A(_02771_),
    .Y(_00488_));
 sky130_fd_sc_hd__buf_4 _16136_ (.A(_08776_),
    .X(_02772_));
 sky130_fd_sc_hd__buf_4 _16137_ (.A(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__buf_4 _16138_ (.A(_02765_),
    .X(_02774_));
 sky130_fd_sc_hd__nor2_1 _16139_ (.A(_10746_),
    .B(_02766_),
    .Y(_02775_));
 sky130_fd_sc_hd__a31o_1 _16140_ (.A1(_02773_),
    .A2(net1581),
    .A3(_02774_),
    .B1(_02775_),
    .X(_00489_));
 sky130_fd_sc_hd__nor2_1 _16141_ (.A(_10698_),
    .B(_02766_),
    .Y(_02776_));
 sky130_fd_sc_hd__a31o_1 _16142_ (.A1(_02773_),
    .A2(net1461),
    .A3(_02774_),
    .B1(_02776_),
    .X(_00490_));
 sky130_fd_sc_hd__and3_1 _16143_ (.A(_02764_),
    .B(_11040_),
    .C(_02752_),
    .X(_02777_));
 sky130_fd_sc_hd__a31o_1 _16144_ (.A1(_02773_),
    .A2(net1479),
    .A3(_02774_),
    .B1(_02777_),
    .X(_00491_));
 sky130_fd_sc_hd__and3_1 _16145_ (.A(_02764_),
    .B(_10587_),
    .C(_02752_),
    .X(_02778_));
 sky130_fd_sc_hd__a31o_1 _16146_ (.A1(_02773_),
    .A2(net1622),
    .A3(_02774_),
    .B1(_02778_),
    .X(_00492_));
 sky130_fd_sc_hd__and3_1 _16147_ (.A(_02764_),
    .B(_11391_),
    .C(_02752_),
    .X(_02779_));
 sky130_fd_sc_hd__a31o_1 _16148_ (.A1(_02773_),
    .A2(net939),
    .A3(_02774_),
    .B1(_02779_),
    .X(_00493_));
 sky130_fd_sc_hd__nor2_1 _16149_ (.A(_10872_),
    .B(_02766_),
    .Y(_02780_));
 sky130_fd_sc_hd__a31o_1 _16150_ (.A1(_02773_),
    .A2(net1485),
    .A3(_02774_),
    .B1(_02780_),
    .X(_00494_));
 sky130_fd_sc_hd__nand2_1 _16151_ (.A(_11547_),
    .B(net3912),
    .Y(_02781_));
 sky130_fd_sc_hd__a22o_1 _16152_ (.A1(_02766_),
    .A2(_02781_),
    .B1(_02770_),
    .B2(_09212_),
    .X(_02782_));
 sky130_fd_sc_hd__inv_2 _16153_ (.A(_02782_),
    .Y(_00495_));
 sky130_fd_sc_hd__nor2_1 _16154_ (.A(_10760_),
    .B(_02766_),
    .Y(_02783_));
 sky130_fd_sc_hd__a31o_1 _16155_ (.A1(_02773_),
    .A2(net2718),
    .A3(_02774_),
    .B1(_02783_),
    .X(_00480_));
 sky130_fd_sc_hd__nand2_1 _16156_ (.A(_11547_),
    .B(net4071),
    .Y(_02784_));
 sky130_fd_sc_hd__a22o_1 _16157_ (.A1(_02766_),
    .A2(_02784_),
    .B1(_02770_),
    .B2(_10313_),
    .X(_02785_));
 sky130_fd_sc_hd__inv_2 _16158_ (.A(_02785_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _16159_ (.A(_11547_),
    .B(net4060),
    .Y(_02786_));
 sky130_fd_sc_hd__a22o_1 _16160_ (.A1(_02765_),
    .A2(_02786_),
    .B1(_02770_),
    .B2(_10316_),
    .X(_02787_));
 sky130_fd_sc_hd__inv_2 _16161_ (.A(_02787_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _16162_ (.A(_11547_),
    .B(net4000),
    .Y(_02788_));
 sky130_fd_sc_hd__a22o_1 _16163_ (.A1(_02765_),
    .A2(_02788_),
    .B1(_02770_),
    .B2(_09589_),
    .X(_02789_));
 sky130_fd_sc_hd__inv_2 _16164_ (.A(_02789_),
    .Y(_00483_));
 sky130_fd_sc_hd__nor2_1 _16165_ (.A(_10767_),
    .B(_02766_),
    .Y(_02790_));
 sky130_fd_sc_hd__a31o_1 _16166_ (.A1(_02773_),
    .A2(net1659),
    .A3(_02774_),
    .B1(_02790_),
    .X(_00484_));
 sky130_fd_sc_hd__nand2_1 _16167_ (.A(_11547_),
    .B(net4190),
    .Y(_02791_));
 sky130_fd_sc_hd__a22o_1 _16168_ (.A1(_02765_),
    .A2(_02791_),
    .B1(_02770_),
    .B2(_09338_),
    .X(_02792_));
 sky130_fd_sc_hd__inv_2 _16169_ (.A(_02792_),
    .Y(_00485_));
 sky130_fd_sc_hd__and3_1 _16170_ (.A(_02764_),
    .B(_11291_),
    .C(_02752_),
    .X(_02793_));
 sky130_fd_sc_hd__a31o_1 _16171_ (.A1(_02773_),
    .A2(net2371),
    .A3(_02774_),
    .B1(_02793_),
    .X(_00486_));
 sky130_fd_sc_hd__nand2_1 _16172_ (.A(_11547_),
    .B(net4128),
    .Y(_02794_));
 sky130_fd_sc_hd__a22o_1 _16173_ (.A1(_02765_),
    .A2(_02794_),
    .B1(_02770_),
    .B2(_09768_),
    .X(_02795_));
 sky130_fd_sc_hd__inv_2 _16174_ (.A(_02795_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_1 _16175_ (.A(_11002_),
    .B(_02766_),
    .Y(_02796_));
 sky130_fd_sc_hd__a31o_1 _16176_ (.A1(_02773_),
    .A2(net801),
    .A3(_02774_),
    .B1(_02796_),
    .X(_00472_));
 sky130_fd_sc_hd__and3_1 _16177_ (.A(_02764_),
    .B(_10667_),
    .C(_02752_),
    .X(_02797_));
 sky130_fd_sc_hd__a31o_1 _16178_ (.A1(_02773_),
    .A2(net1881),
    .A3(_02774_),
    .B1(_02797_),
    .X(_00473_));
 sky130_fd_sc_hd__nor2_1 _16179_ (.A(_10669_),
    .B(_02766_),
    .Y(_02798_));
 sky130_fd_sc_hd__a31o_1 _16180_ (.A1(_02773_),
    .A2(net1915),
    .A3(_02774_),
    .B1(_02798_),
    .X(_00474_));
 sky130_fd_sc_hd__nand2_1 _16181_ (.A(_11547_),
    .B(net4076),
    .Y(_02799_));
 sky130_fd_sc_hd__a22o_1 _16182_ (.A1(_02765_),
    .A2(_02799_),
    .B1(_02770_),
    .B2(_09256_),
    .X(_02800_));
 sky130_fd_sc_hd__inv_2 _16183_ (.A(_02800_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _16184_ (.A(_11010_),
    .B(_02766_),
    .Y(_02801_));
 sky130_fd_sc_hd__a31o_1 _16185_ (.A1(_02773_),
    .A2(net1163),
    .A3(_02774_),
    .B1(_02801_),
    .X(_00476_));
 sky130_fd_sc_hd__nand2_1 _16186_ (.A(_11547_),
    .B(net4156),
    .Y(_02802_));
 sky130_fd_sc_hd__a22o_1 _16187_ (.A1(_02765_),
    .A2(_02802_),
    .B1(_02770_),
    .B2(_10331_),
    .X(_02803_));
 sky130_fd_sc_hd__inv_2 _16188_ (.A(_02803_),
    .Y(_00477_));
 sky130_fd_sc_hd__and3_1 _16189_ (.A(_02764_),
    .B(_10617_),
    .C(_02752_),
    .X(_02804_));
 sky130_fd_sc_hd__a31o_1 _16190_ (.A1(_02773_),
    .A2(net1133),
    .A3(_02774_),
    .B1(_02804_),
    .X(_00478_));
 sky130_fd_sc_hd__nand2_1 _16191_ (.A(_11547_),
    .B(net4094),
    .Y(_02805_));
 sky130_fd_sc_hd__a22o_1 _16192_ (.A1(_02765_),
    .A2(_02805_),
    .B1(_02770_),
    .B2(_10335_),
    .X(_02806_));
 sky130_fd_sc_hd__inv_2 _16193_ (.A(_02806_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _16194_ (.A(_11547_),
    .B(net4147),
    .Y(_02807_));
 sky130_fd_sc_hd__a22o_1 _16195_ (.A1(_02765_),
    .A2(_02807_),
    .B1(_02770_),
    .B2(_09495_),
    .X(_02808_));
 sky130_fd_sc_hd__inv_2 _16196_ (.A(_02808_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_1 _16197_ (.A(_10681_),
    .B(_02766_),
    .Y(_02809_));
 sky130_fd_sc_hd__a31o_1 _16198_ (.A1(_02773_),
    .A2(net1721),
    .A3(_02774_),
    .B1(_02809_),
    .X(_00465_));
 sky130_fd_sc_hd__and3_1 _16199_ (.A(_02764_),
    .B(_10728_),
    .C(_02752_),
    .X(_02810_));
 sky130_fd_sc_hd__a31o_1 _16200_ (.A1(_02773_),
    .A2(net1235),
    .A3(_02774_),
    .B1(_02810_),
    .X(_00466_));
 sky130_fd_sc_hd__nand2_1 _16201_ (.A(_11547_),
    .B(net4089),
    .Y(_02811_));
 sky130_fd_sc_hd__a22o_1 _16202_ (.A1(_02765_),
    .A2(_02811_),
    .B1(_02770_),
    .B2(_10342_),
    .X(_02812_));
 sky130_fd_sc_hd__inv_2 _16203_ (.A(_02812_),
    .Y(_00467_));
 sky130_fd_sc_hd__buf_4 _16204_ (.A(_02772_),
    .X(_02813_));
 sky130_fd_sc_hd__and3_1 _16205_ (.A(_02764_),
    .B(_10848_),
    .C(_02752_),
    .X(_02814_));
 sky130_fd_sc_hd__a31o_1 _16206_ (.A1(_02813_),
    .A2(net1707),
    .A3(_02766_),
    .B1(_02814_),
    .X(_00468_));
 sky130_fd_sc_hd__nand2_1 _16207_ (.A(_11547_),
    .B(net4033),
    .Y(_02815_));
 sky130_fd_sc_hd__a22o_1 _16208_ (.A1(_02765_),
    .A2(_02815_),
    .B1(_02770_),
    .B2(net136),
    .X(_02816_));
 sky130_fd_sc_hd__inv_2 _16209_ (.A(_02816_),
    .Y(_00469_));
 sky130_fd_sc_hd__clkbuf_8 _16210_ (.A(_11151_),
    .X(_02817_));
 sky130_fd_sc_hd__nand2_1 _16211_ (.A(_02817_),
    .B(net3234),
    .Y(_02818_));
 sky130_fd_sc_hd__a22o_1 _16212_ (.A1(_10348_),
    .A2(_02764_),
    .B1(_02766_),
    .B2(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__inv_2 _16213_ (.A(_02819_),
    .Y(_00470_));
 sky130_fd_sc_hd__nor2_1 _16214_ (.A(_09300_),
    .B(_02766_),
    .Y(_02820_));
 sky130_fd_sc_hd__a31o_1 _16215_ (.A1(_02813_),
    .A2(net1620),
    .A3(_02766_),
    .B1(_02820_),
    .X(_00471_));
 sky130_fd_sc_hd__nor2_4 _16216_ (.A(_11620_),
    .B(_10356_),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_4 _16217_ (.A(_02821_),
    .B(_09225_),
    .Y(_02822_));
 sky130_fd_sc_hd__buf_4 _16218_ (.A(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__buf_4 _16219_ (.A(_02822_),
    .X(_02824_));
 sky130_fd_sc_hd__nor2_1 _16220_ (.A(_11210_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__a31o_1 _16221_ (.A1(_02813_),
    .A2(net1719),
    .A3(_02823_),
    .B1(_02825_),
    .X(_00456_));
 sky130_fd_sc_hd__nor2_1 _16222_ (.A(_10746_),
    .B(_02824_),
    .Y(_02826_));
 sky130_fd_sc_hd__a31o_1 _16223_ (.A1(_02813_),
    .A2(net2551),
    .A3(_02823_),
    .B1(_02826_),
    .X(_00457_));
 sky130_fd_sc_hd__nor2_1 _16224_ (.A(_10698_),
    .B(_02824_),
    .Y(_02827_));
 sky130_fd_sc_hd__a31o_1 _16225_ (.A1(_02813_),
    .A2(net2611),
    .A3(_02823_),
    .B1(_02827_),
    .X(_00458_));
 sky130_fd_sc_hd__and3_1 _16226_ (.A(_02821_),
    .B(_11040_),
    .C(_02752_),
    .X(_02828_));
 sky130_fd_sc_hd__a31o_1 _16227_ (.A1(_02813_),
    .A2(net2555),
    .A3(_02823_),
    .B1(_02828_),
    .X(_00459_));
 sky130_fd_sc_hd__and3_1 _16228_ (.A(_02821_),
    .B(_10587_),
    .C(_02752_),
    .X(_02829_));
 sky130_fd_sc_hd__a31o_1 _16229_ (.A1(_02813_),
    .A2(net991),
    .A3(_02823_),
    .B1(_02829_),
    .X(_00460_));
 sky130_fd_sc_hd__and3_1 _16230_ (.A(_02821_),
    .B(_11391_),
    .C(_02752_),
    .X(_02830_));
 sky130_fd_sc_hd__a31o_1 _16231_ (.A1(_02813_),
    .A2(net2542),
    .A3(_02823_),
    .B1(_02830_),
    .X(_00461_));
 sky130_fd_sc_hd__buf_4 _16232_ (.A(_10930_),
    .X(_02831_));
 sky130_fd_sc_hd__nand2_1 _16233_ (.A(_02831_),
    .B(net4072),
    .Y(_02832_));
 sky130_fd_sc_hd__and3_1 _16234_ (.A(_10355_),
    .B(_02768_),
    .C(_08725_),
    .X(_02833_));
 sky130_fd_sc_hd__buf_4 _16235_ (.A(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__a22o_1 _16236_ (.A1(_02824_),
    .A2(_02832_),
    .B1(_02834_),
    .B2(_09398_),
    .X(_02835_));
 sky130_fd_sc_hd__inv_2 _16237_ (.A(_02835_),
    .Y(_00462_));
 sky130_fd_sc_hd__and3_1 _16238_ (.A(_02821_),
    .B(_10874_),
    .C(_02752_),
    .X(_02836_));
 sky130_fd_sc_hd__a31o_1 _16239_ (.A1(_02813_),
    .A2(net2525),
    .A3(_02823_),
    .B1(_02836_),
    .X(_00463_));
 sky130_fd_sc_hd__nand2_1 _16240_ (.A(_02831_),
    .B(net4027),
    .Y(_02837_));
 sky130_fd_sc_hd__a22o_1 _16241_ (.A1(_02824_),
    .A2(_02837_),
    .B1(_02834_),
    .B2(_09531_),
    .X(_02838_));
 sky130_fd_sc_hd__inv_2 _16242_ (.A(_02838_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _16243_ (.A(_02831_),
    .B(net4246),
    .Y(_02839_));
 sky130_fd_sc_hd__a22o_1 _16244_ (.A1(_02824_),
    .A2(_02839_),
    .B1(_02834_),
    .B2(_10313_),
    .X(_02840_));
 sky130_fd_sc_hd__inv_2 _16245_ (.A(_02840_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _16246_ (.A(_02831_),
    .B(net4214),
    .Y(_02841_));
 sky130_fd_sc_hd__a22o_1 _16247_ (.A1(_02824_),
    .A2(_02841_),
    .B1(_02834_),
    .B2(_10316_),
    .X(_02842_));
 sky130_fd_sc_hd__inv_2 _16248_ (.A(_02842_),
    .Y(_00450_));
 sky130_fd_sc_hd__nor2_1 _16249_ (.A(_10657_),
    .B(_02824_),
    .Y(_02843_));
 sky130_fd_sc_hd__a31o_1 _16250_ (.A1(_02813_),
    .A2(net2596),
    .A3(_02823_),
    .B1(_02843_),
    .X(_00451_));
 sky130_fd_sc_hd__nor2_1 _16251_ (.A(_10767_),
    .B(_02824_),
    .Y(_02844_));
 sky130_fd_sc_hd__a31o_1 _16252_ (.A1(_02813_),
    .A2(net843),
    .A3(_02823_),
    .B1(_02844_),
    .X(_00452_));
 sky130_fd_sc_hd__clkbuf_16 _16253_ (.A(_09235_),
    .X(_02845_));
 sky130_fd_sc_hd__nor2_1 _16254_ (.A(_02845_),
    .B(_02824_),
    .Y(_02846_));
 sky130_fd_sc_hd__a31o_1 _16255_ (.A1(_02813_),
    .A2(net2549),
    .A3(_02823_),
    .B1(_02846_),
    .X(_00453_));
 sky130_fd_sc_hd__and3_1 _16256_ (.A(_02821_),
    .B(_11291_),
    .C(_02752_),
    .X(_02847_));
 sky130_fd_sc_hd__a31o_1 _16257_ (.A1(_02813_),
    .A2(net967),
    .A3(_02823_),
    .B1(_02847_),
    .X(_00454_));
 sky130_fd_sc_hd__nand2_1 _16258_ (.A(_02831_),
    .B(net4260),
    .Y(_02848_));
 sky130_fd_sc_hd__a22o_1 _16259_ (.A1(_02822_),
    .A2(_02848_),
    .B1(_02834_),
    .B2(_09768_),
    .X(_02849_));
 sky130_fd_sc_hd__inv_2 _16260_ (.A(_02849_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _16261_ (.A(_02831_),
    .B(net4189),
    .Y(_02850_));
 sky130_fd_sc_hd__a22o_1 _16262_ (.A1(_02822_),
    .A2(_02850_),
    .B1(_02834_),
    .B2(_09415_),
    .X(_02851_));
 sky130_fd_sc_hd__inv_2 _16263_ (.A(_02851_),
    .Y(_00432_));
 sky130_fd_sc_hd__and3_1 _16264_ (.A(_02821_),
    .B(_10667_),
    .C(_02752_),
    .X(_02852_));
 sky130_fd_sc_hd__a31o_1 _16265_ (.A1(_02813_),
    .A2(net1405),
    .A3(_02823_),
    .B1(_02852_),
    .X(_00433_));
 sky130_fd_sc_hd__nor2_1 _16266_ (.A(_10669_),
    .B(_02824_),
    .Y(_02853_));
 sky130_fd_sc_hd__a31o_1 _16267_ (.A1(_02813_),
    .A2(net1181),
    .A3(_02823_),
    .B1(_02853_),
    .X(_00434_));
 sky130_fd_sc_hd__buf_4 _16268_ (.A(_11219_),
    .X(_02854_));
 sky130_fd_sc_hd__and3_1 _16269_ (.A(_02821_),
    .B(_10500_),
    .C(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__a31o_1 _16270_ (.A1(_02813_),
    .A2(net755),
    .A3(_02823_),
    .B1(_02855_),
    .X(_00435_));
 sky130_fd_sc_hd__buf_4 _16271_ (.A(_02772_),
    .X(_02856_));
 sky130_fd_sc_hd__nor2_1 _16272_ (.A(_11010_),
    .B(_02824_),
    .Y(_02857_));
 sky130_fd_sc_hd__a31o_1 _16273_ (.A1(_02856_),
    .A2(net2263),
    .A3(_02823_),
    .B1(_02857_),
    .X(_00436_));
 sky130_fd_sc_hd__nand2_1 _16274_ (.A(_02831_),
    .B(net4173),
    .Y(_02858_));
 sky130_fd_sc_hd__a22o_1 _16275_ (.A1(_02822_),
    .A2(_02858_),
    .B1(_02834_),
    .B2(_10331_),
    .X(_02859_));
 sky130_fd_sc_hd__inv_2 _16276_ (.A(_02859_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _16277_ (.A(_02831_),
    .B(net4108),
    .Y(_02860_));
 sky130_fd_sc_hd__a22o_1 _16278_ (.A1(_02822_),
    .A2(_02860_),
    .B1(_02834_),
    .B2(_09425_),
    .X(_02861_));
 sky130_fd_sc_hd__inv_2 _16279_ (.A(_02861_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _16280_ (.A(_02831_),
    .B(net4165),
    .Y(_02862_));
 sky130_fd_sc_hd__a22o_1 _16281_ (.A1(_02822_),
    .A2(_02862_),
    .B1(_02834_),
    .B2(_10335_),
    .X(_02863_));
 sky130_fd_sc_hd__inv_2 _16282_ (.A(_02863_),
    .Y(_00439_));
 sky130_fd_sc_hd__and3_1 _16283_ (.A(_02821_),
    .B(_10679_),
    .C(_02854_),
    .X(_02864_));
 sky130_fd_sc_hd__a31o_1 _16284_ (.A1(_02856_),
    .A2(net1223),
    .A3(_02823_),
    .B1(_02864_),
    .X(_00424_));
 sky130_fd_sc_hd__nor2_1 _16285_ (.A(_10681_),
    .B(_02824_),
    .Y(_02865_));
 sky130_fd_sc_hd__a31o_1 _16286_ (.A1(_02856_),
    .A2(net1125),
    .A3(_02824_),
    .B1(_02865_),
    .X(_00425_));
 sky130_fd_sc_hd__nand2_1 _16287_ (.A(_02831_),
    .B(net4114),
    .Y(_02866_));
 sky130_fd_sc_hd__a22o_1 _16288_ (.A1(_02822_),
    .A2(_02866_),
    .B1(_02834_),
    .B2(_09280_),
    .X(_02867_));
 sky130_fd_sc_hd__inv_2 _16289_ (.A(_02867_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _16290_ (.A(_02831_),
    .B(net3990),
    .Y(_02868_));
 sky130_fd_sc_hd__a22o_1 _16291_ (.A1(_02822_),
    .A2(_02868_),
    .B1(_02834_),
    .B2(_10342_),
    .X(_02869_));
 sky130_fd_sc_hd__inv_2 _16292_ (.A(_02869_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _16293_ (.A(_02831_),
    .B(net3948),
    .Y(_02870_));
 sky130_fd_sc_hd__a22o_1 _16294_ (.A1(_02822_),
    .A2(_02870_),
    .B1(_02834_),
    .B2(_09288_),
    .X(_02871_));
 sky130_fd_sc_hd__inv_2 _16295_ (.A(_02871_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _16296_ (.A(_02831_),
    .B(net4111),
    .Y(_02872_));
 sky130_fd_sc_hd__a22o_1 _16297_ (.A1(_02822_),
    .A2(_02872_),
    .B1(_02834_),
    .B2(net136),
    .X(_02873_));
 sky130_fd_sc_hd__inv_2 _16298_ (.A(_02873_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _16299_ (.A(_02817_),
    .B(net3541),
    .Y(_02874_));
 sky130_fd_sc_hd__a22o_1 _16300_ (.A1(_10348_),
    .A2(_02821_),
    .B1(_02824_),
    .B2(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__inv_2 _16301_ (.A(net3542),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _16302_ (.A(_02817_),
    .B(net3812),
    .Y(_02876_));
 sky130_fd_sc_hd__a22o_1 _16303_ (.A1(_09440_),
    .A2(_02821_),
    .B1(_02824_),
    .B2(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__inv_2 _16304_ (.A(net3813),
    .Y(_00431_));
 sky130_fd_sc_hd__nor2_2 _16305_ (.A(_11620_),
    .B(_10411_),
    .Y(_02878_));
 sky130_fd_sc_hd__inv_2 _16306_ (.A(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__nor2_8 _16307_ (.A(_08797_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__nor2_1 _16308_ (.A(_09304_),
    .B(_02879_),
    .Y(_02881_));
 sky130_fd_sc_hd__clkinv_4 _16309_ (.A(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__buf_4 _16310_ (.A(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__nand2_1 _16311_ (.A(_02817_),
    .B(net3440),
    .Y(_02884_));
 sky130_fd_sc_hd__a22o_1 _16312_ (.A1(_02880_),
    .A2(_10239_),
    .B1(_02883_),
    .B2(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__inv_2 _16313_ (.A(_02885_),
    .Y(_00416_));
 sky130_fd_sc_hd__buf_4 _16314_ (.A(_02882_),
    .X(_02886_));
 sky130_fd_sc_hd__nor2_1 _16315_ (.A(_10746_),
    .B(_02883_),
    .Y(_02887_));
 sky130_fd_sc_hd__a31o_1 _16316_ (.A1(_02856_),
    .A2(net2298),
    .A3(_02886_),
    .B1(_02887_),
    .X(_00417_));
 sky130_fd_sc_hd__nand2_1 _16317_ (.A(_02817_),
    .B(net3365),
    .Y(_02888_));
 sky130_fd_sc_hd__a22o_1 _16318_ (.A1(_02880_),
    .A2(_09459_),
    .B1(_02883_),
    .B2(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__inv_2 _16319_ (.A(_02889_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _16320_ (.A(_02817_),
    .B(net3286),
    .Y(_02890_));
 sky130_fd_sc_hd__a22o_1 _16321_ (.A1(_02880_),
    .A2(_10983_),
    .B1(_02883_),
    .B2(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__inv_2 _16322_ (.A(_02891_),
    .Y(_00419_));
 sky130_fd_sc_hd__and3_1 _16323_ (.A(_02878_),
    .B(_10587_),
    .C(_02854_),
    .X(_02892_));
 sky130_fd_sc_hd__a31o_1 _16324_ (.A1(_02886_),
    .A2(_02751_),
    .A3(net2355),
    .B1(_02892_),
    .X(_00420_));
 sky130_fd_sc_hd__nand2_1 _16325_ (.A(_02817_),
    .B(net3113),
    .Y(_02893_));
 sky130_fd_sc_hd__a22o_1 _16326_ (.A1(_02880_),
    .A2(_10869_),
    .B1(_02883_),
    .B2(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__inv_2 _16327_ (.A(_02894_),
    .Y(_00421_));
 sky130_fd_sc_hd__nor2_1 _16328_ (.A(_10872_),
    .B(_02883_),
    .Y(_02895_));
 sky130_fd_sc_hd__a31o_1 _16329_ (.A1(_02856_),
    .A2(net2453),
    .A3(_02886_),
    .B1(_02895_),
    .X(_00422_));
 sky130_fd_sc_hd__nand2_1 _16330_ (.A(_02817_),
    .B(net3526),
    .Y(_02896_));
 sky130_fd_sc_hd__a22o_1 _16331_ (.A1(_02880_),
    .A2(_10591_),
    .B1(_02882_),
    .B2(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__inv_2 _16332_ (.A(_02897_),
    .Y(_00423_));
 sky130_fd_sc_hd__nor2_1 _16333_ (.A(_10760_),
    .B(_02883_),
    .Y(_02898_));
 sky130_fd_sc_hd__a31o_1 _16334_ (.A1(_02856_),
    .A2(net1161),
    .A3(_02886_),
    .B1(_02898_),
    .X(_00408_));
 sky130_fd_sc_hd__clkbuf_16 _16335_ (.A(_09218_),
    .X(_02899_));
 sky130_fd_sc_hd__nand2_1 _16336_ (.A(_02817_),
    .B(net3888),
    .Y(_02900_));
 sky130_fd_sc_hd__a22o_1 _16337_ (.A1(_02880_),
    .A2(_02899_),
    .B1(_02882_),
    .B2(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__inv_2 _16338_ (.A(_02901_),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _16339_ (.A(_02817_),
    .B(net3693),
    .Y(_02902_));
 sky130_fd_sc_hd__a22o_1 _16340_ (.A1(_02880_),
    .A2(_10195_),
    .B1(_02882_),
    .B2(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__inv_2 _16341_ (.A(_02903_),
    .Y(_00410_));
 sky130_fd_sc_hd__clkbuf_16 _16342_ (.A(_09229_),
    .X(_02904_));
 sky130_fd_sc_hd__nor2_1 _16343_ (.A(_02904_),
    .B(_02883_),
    .Y(_02905_));
 sky130_fd_sc_hd__a31o_1 _16344_ (.A1(_02856_),
    .A2(net2469),
    .A3(_02886_),
    .B1(_02905_),
    .X(_00411_));
 sky130_fd_sc_hd__nor2_1 _16345_ (.A(_10767_),
    .B(_02883_),
    .Y(_02906_));
 sky130_fd_sc_hd__a31o_1 _16346_ (.A1(_02856_),
    .A2(net1531),
    .A3(_02886_),
    .B1(_02906_),
    .X(_00412_));
 sky130_fd_sc_hd__nor2_1 _16347_ (.A(_02845_),
    .B(_02883_),
    .Y(_02907_));
 sky130_fd_sc_hd__a31o_1 _16348_ (.A1(_02856_),
    .A2(net2462),
    .A3(_02886_),
    .B1(_02907_),
    .X(_00413_));
 sky130_fd_sc_hd__and3_1 _16349_ (.A(_02878_),
    .B(_11291_),
    .C(_02854_),
    .X(_02908_));
 sky130_fd_sc_hd__a31o_1 _16350_ (.A1(_02886_),
    .A2(_02751_),
    .A3(net2032),
    .B1(_02908_),
    .X(_00414_));
 sky130_fd_sc_hd__nor2_1 _16351_ (.A(_10663_),
    .B(_02883_),
    .Y(_02909_));
 sky130_fd_sc_hd__a31o_1 _16352_ (.A1(_02856_),
    .A2(net2515),
    .A3(_02886_),
    .B1(_02909_),
    .X(_00415_));
 sky130_fd_sc_hd__nor2_1 _16353_ (.A(_11002_),
    .B(_02883_),
    .Y(_02910_));
 sky130_fd_sc_hd__a31o_1 _16354_ (.A1(_02856_),
    .A2(net2361),
    .A3(_02886_),
    .B1(_02910_),
    .X(_00400_));
 sky130_fd_sc_hd__and3_1 _16355_ (.A(_02878_),
    .B(_10667_),
    .C(_02854_),
    .X(_02911_));
 sky130_fd_sc_hd__a31o_1 _16356_ (.A1(_02886_),
    .A2(_02751_),
    .A3(net2599),
    .B1(_02911_),
    .X(_00401_));
 sky130_fd_sc_hd__nor2_1 _16357_ (.A(_10669_),
    .B(_02883_),
    .Y(_02912_));
 sky130_fd_sc_hd__a31o_1 _16358_ (.A1(_02856_),
    .A2(net1847),
    .A3(_02883_),
    .B1(_02912_),
    .X(_00402_));
 sky130_fd_sc_hd__nand2_1 _16359_ (.A(_02817_),
    .B(net4255),
    .Y(_02913_));
 sky130_fd_sc_hd__a22o_1 _16360_ (.A1(_02880_),
    .A2(_09256_),
    .B1(_02882_),
    .B2(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__inv_2 _16361_ (.A(_02914_),
    .Y(_00403_));
 sky130_fd_sc_hd__nor2_1 _16362_ (.A(_11010_),
    .B(_02883_),
    .Y(_02915_));
 sky130_fd_sc_hd__a31o_1 _16363_ (.A1(_02856_),
    .A2(net2593),
    .A3(_02883_),
    .B1(_02915_),
    .X(_00404_));
 sky130_fd_sc_hd__clkbuf_16 _16364_ (.A(net145),
    .X(_02916_));
 sky130_fd_sc_hd__nand2_1 _16365_ (.A(_02817_),
    .B(net3802),
    .Y(_02917_));
 sky130_fd_sc_hd__a22o_1 _16366_ (.A1(_02880_),
    .A2(_02916_),
    .B1(_02882_),
    .B2(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__inv_2 _16367_ (.A(_02918_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _16368_ (.A(_02817_),
    .B(net3837),
    .Y(_02919_));
 sky130_fd_sc_hd__a22o_1 _16369_ (.A1(_02880_),
    .A2(_09425_),
    .B1(_02882_),
    .B2(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__inv_2 _16370_ (.A(_02920_),
    .Y(_00406_));
 sky130_fd_sc_hd__buf_8 _16371_ (.A(net144),
    .X(_02921_));
 sky130_fd_sc_hd__nand2_1 _16372_ (.A(_02817_),
    .B(net4056),
    .Y(_02922_));
 sky130_fd_sc_hd__a22o_1 _16373_ (.A1(_02880_),
    .A2(_02921_),
    .B1(_02882_),
    .B2(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__inv_2 _16374_ (.A(_02923_),
    .Y(_00407_));
 sky130_fd_sc_hd__and3_1 _16375_ (.A(_02878_),
    .B(_10679_),
    .C(_02854_),
    .X(_02924_));
 sky130_fd_sc_hd__a31o_1 _16376_ (.A1(_02886_),
    .A2(_02751_),
    .A3(net2038),
    .B1(_02924_),
    .X(_00392_));
 sky130_fd_sc_hd__nand2_1 _16377_ (.A(_02817_),
    .B(net3897),
    .Y(_02925_));
 sky130_fd_sc_hd__a22o_1 _16378_ (.A1(_02880_),
    .A2(_09365_),
    .B1(_02882_),
    .B2(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__inv_2 _16379_ (.A(_02926_),
    .Y(_00393_));
 sky130_fd_sc_hd__and3_1 _16380_ (.A(_02878_),
    .B(_10728_),
    .C(_02854_),
    .X(_02927_));
 sky130_fd_sc_hd__a31o_1 _16381_ (.A1(_02886_),
    .A2(_02751_),
    .A3(net2015),
    .B1(_02927_),
    .X(_00394_));
 sky130_fd_sc_hd__buf_12 _16382_ (.A(net140),
    .X(_02928_));
 sky130_fd_sc_hd__nand2_1 _16383_ (.A(_02817_),
    .B(net4265),
    .Y(_02929_));
 sky130_fd_sc_hd__a22o_1 _16384_ (.A1(_02880_),
    .A2(_02928_),
    .B1(_02882_),
    .B2(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__inv_2 _16385_ (.A(_02930_),
    .Y(_00395_));
 sky130_fd_sc_hd__buf_4 _16386_ (.A(_11151_),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_1 _16387_ (.A(_02931_),
    .B(net4061),
    .Y(_02932_));
 sky130_fd_sc_hd__a22o_1 _16388_ (.A1(_02880_),
    .A2(net139),
    .B1(_02882_),
    .B2(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__inv_2 _16389_ (.A(_02933_),
    .Y(_00396_));
 sky130_fd_sc_hd__and3_1 _16390_ (.A(_02878_),
    .B(_11426_),
    .C(_02854_),
    .X(_02934_));
 sky130_fd_sc_hd__a31o_1 _16391_ (.A1(_02886_),
    .A2(_02751_),
    .A3(net2616),
    .B1(_02934_),
    .X(_00397_));
 sky130_fd_sc_hd__clkbuf_8 _16392_ (.A(_09375_),
    .X(_02935_));
 sky130_fd_sc_hd__nand2_1 _16393_ (.A(_02935_),
    .B(net4233),
    .Y(_02936_));
 sky130_fd_sc_hd__o2bb2a_1 _16394_ (.A1_N(_02936_),
    .A2_N(_02886_),
    .B1(_10289_),
    .B2(_02879_),
    .X(_00398_));
 sky130_fd_sc_hd__nand2_1 _16395_ (.A(_02935_),
    .B(net4055),
    .Y(_02937_));
 sky130_fd_sc_hd__o2bb2a_1 _16396_ (.A1_N(_02937_),
    .A2_N(_02886_),
    .B1(_11316_),
    .B2(_02879_),
    .X(_00399_));
 sky130_fd_sc_hd__nand2_8 _16397_ (.A(_11161_),
    .B(_09982_),
    .Y(_02938_));
 sky130_fd_sc_hd__nor2_2 _16398_ (.A(_02938_),
    .B(_10469_),
    .Y(_02939_));
 sky130_fd_sc_hd__inv_2 _16399_ (.A(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__nor2_1 _16400_ (.A(_09304_),
    .B(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__clkinv_4 _16401_ (.A(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__buf_4 _16402_ (.A(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__buf_4 _16403_ (.A(_02942_),
    .X(_02944_));
 sky130_fd_sc_hd__nor2_1 _16404_ (.A(_11210_),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__a31o_1 _16405_ (.A1(_02856_),
    .A2(net2136),
    .A3(_02943_),
    .B1(_02945_),
    .X(_00384_));
 sky130_fd_sc_hd__nor2_1 _16406_ (.A(_10746_),
    .B(_02944_),
    .Y(_02946_));
 sky130_fd_sc_hd__a31o_1 _16407_ (.A1(_02856_),
    .A2(net2490),
    .A3(_02943_),
    .B1(_02946_),
    .X(_00385_));
 sky130_fd_sc_hd__nor2_1 _16408_ (.A(_10698_),
    .B(_02944_),
    .Y(_02947_));
 sky130_fd_sc_hd__a31o_1 _16409_ (.A1(_02856_),
    .A2(net2584),
    .A3(_02943_),
    .B1(_02947_),
    .X(_00386_));
 sky130_fd_sc_hd__nor2_4 _16410_ (.A(_09190_),
    .B(_02940_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_1 _16411_ (.A(_02931_),
    .B(net3353),
    .Y(_02949_));
 sky130_fd_sc_hd__a22o_1 _16412_ (.A1(_02948_),
    .A2(_10983_),
    .B1(_02944_),
    .B2(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__inv_2 _16413_ (.A(_02950_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _16414_ (.A(_02931_),
    .B(net3193),
    .Y(_02951_));
 sky130_fd_sc_hd__a22o_1 _16415_ (.A1(_02948_),
    .A2(_11330_),
    .B1(_02944_),
    .B2(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__inv_2 _16416_ (.A(_02952_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _16417_ (.A(_02931_),
    .B(net3106),
    .Y(_02953_));
 sky130_fd_sc_hd__a22o_1 _16418_ (.A1(_02948_),
    .A2(_10869_),
    .B1(_02942_),
    .B2(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__inv_2 _16419_ (.A(_02954_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _16420_ (.A(_02931_),
    .B(net3441),
    .Y(_02955_));
 sky130_fd_sc_hd__a22o_1 _16421_ (.A1(_02948_),
    .A2(_11105_),
    .B1(_02942_),
    .B2(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__inv_2 _16422_ (.A(_02956_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _16423_ (.A(_02931_),
    .B(net3044),
    .Y(_02957_));
 sky130_fd_sc_hd__a22o_1 _16424_ (.A1(_02948_),
    .A2(_10591_),
    .B1(_02942_),
    .B2(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__inv_2 _16425_ (.A(_02958_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_1 _16426_ (.A(_02931_),
    .B(net3385),
    .Y(_02959_));
 sky130_fd_sc_hd__a22o_1 _16427_ (.A1(_02948_),
    .A2(net135),
    .B1(_02942_),
    .B2(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__inv_2 _16428_ (.A(_02960_),
    .Y(_00376_));
 sky130_fd_sc_hd__nand2_1 _16429_ (.A(_02931_),
    .B(net3199),
    .Y(_02961_));
 sky130_fd_sc_hd__a22o_1 _16430_ (.A1(_02948_),
    .A2(_02899_),
    .B1(_02942_),
    .B2(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__inv_2 _16431_ (.A(_02962_),
    .Y(_00377_));
 sky130_fd_sc_hd__buf_12 _16432_ (.A(_09331_),
    .X(_02963_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(_02931_),
    .B(net2842),
    .Y(_02964_));
 sky130_fd_sc_hd__a22o_1 _16434_ (.A1(_02948_),
    .A2(_02963_),
    .B1(_02942_),
    .B2(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__inv_2 _16435_ (.A(_02965_),
    .Y(_00378_));
 sky130_fd_sc_hd__buf_4 _16436_ (.A(_02772_),
    .X(_02966_));
 sky130_fd_sc_hd__nor2_1 _16437_ (.A(_02904_),
    .B(_02944_),
    .Y(_02967_));
 sky130_fd_sc_hd__a31o_1 _16438_ (.A1(_02966_),
    .A2(net1956),
    .A3(_02943_),
    .B1(_02967_),
    .X(_00379_));
 sky130_fd_sc_hd__nor2_1 _16439_ (.A(_10767_),
    .B(_02944_),
    .Y(_02968_));
 sky130_fd_sc_hd__a31o_1 _16440_ (.A1(_02966_),
    .A2(net1995),
    .A3(_02943_),
    .B1(_02968_),
    .X(_00380_));
 sky130_fd_sc_hd__nor2_1 _16441_ (.A(_02845_),
    .B(_02944_),
    .Y(_02969_));
 sky130_fd_sc_hd__a31o_1 _16442_ (.A1(_02966_),
    .A2(net1199),
    .A3(_02943_),
    .B1(_02969_),
    .X(_00381_));
 sky130_fd_sc_hd__and3_1 _16443_ (.A(_02939_),
    .B(_11291_),
    .C(_02854_),
    .X(_02970_));
 sky130_fd_sc_hd__a31o_1 _16444_ (.A1(_02943_),
    .A2(_02751_),
    .A3(net1904),
    .B1(_02970_),
    .X(_00382_));
 sky130_fd_sc_hd__nor2_1 _16445_ (.A(_10663_),
    .B(_02944_),
    .Y(_02971_));
 sky130_fd_sc_hd__a31o_1 _16446_ (.A1(_02966_),
    .A2(net1459),
    .A3(_02943_),
    .B1(_02971_),
    .X(_00383_));
 sky130_fd_sc_hd__nor2_1 _16447_ (.A(_11002_),
    .B(_02944_),
    .Y(_02972_));
 sky130_fd_sc_hd__a31o_1 _16448_ (.A1(_02966_),
    .A2(net1147),
    .A3(_02943_),
    .B1(_02972_),
    .X(_00368_));
 sky130_fd_sc_hd__and3_1 _16449_ (.A(_02939_),
    .B(_10667_),
    .C(_02854_),
    .X(_02973_));
 sky130_fd_sc_hd__a31o_1 _16450_ (.A1(_02943_),
    .A2(_02751_),
    .A3(net2439),
    .B1(_02973_),
    .X(_00369_));
 sky130_fd_sc_hd__nand2_1 _16451_ (.A(_02931_),
    .B(net3072),
    .Y(_02974_));
 sky130_fd_sc_hd__a22o_1 _16452_ (.A1(_02948_),
    .A2(_09347_),
    .B1(_02942_),
    .B2(_02974_),
    .X(_02975_));
 sky130_fd_sc_hd__inv_2 _16453_ (.A(_02975_),
    .Y(_00370_));
 sky130_fd_sc_hd__and3_1 _16454_ (.A(_02939_),
    .B(_10500_),
    .C(_02854_),
    .X(_02976_));
 sky130_fd_sc_hd__a31o_1 _16455_ (.A1(_02943_),
    .A2(_02751_),
    .A3(net2557),
    .B1(_02976_),
    .X(_00371_));
 sky130_fd_sc_hd__nor2_1 _16456_ (.A(_11010_),
    .B(_02944_),
    .Y(_02977_));
 sky130_fd_sc_hd__a31o_1 _16457_ (.A1(_02966_),
    .A2(net1027),
    .A3(_02944_),
    .B1(_02977_),
    .X(_00372_));
 sky130_fd_sc_hd__nand2_1 _16458_ (.A(_02931_),
    .B(net2871),
    .Y(_02978_));
 sky130_fd_sc_hd__a22o_1 _16459_ (.A1(_02948_),
    .A2(_02916_),
    .B1(_02942_),
    .B2(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__inv_2 _16460_ (.A(_02979_),
    .Y(_00373_));
 sky130_fd_sc_hd__and3_1 _16461_ (.A(_02939_),
    .B(_10617_),
    .C(_02854_),
    .X(_02980_));
 sky130_fd_sc_hd__a31o_1 _16462_ (.A1(_02943_),
    .A2(_02751_),
    .A3(net2346),
    .B1(_02980_),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_1 _16463_ (.A(_02931_),
    .B(net2937),
    .Y(_02981_));
 sky130_fd_sc_hd__a22o_1 _16464_ (.A1(_02948_),
    .A2(_02921_),
    .B1(_02942_),
    .B2(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__inv_2 _16465_ (.A(_02982_),
    .Y(_00375_));
 sky130_fd_sc_hd__and3_1 _16466_ (.A(_02939_),
    .B(_10679_),
    .C(_02854_),
    .X(_02983_));
 sky130_fd_sc_hd__a31o_1 _16467_ (.A1(_02943_),
    .A2(_02751_),
    .A3(net2096),
    .B1(_02983_),
    .X(_00360_));
 sky130_fd_sc_hd__nor2_1 _16468_ (.A(_10681_),
    .B(_02944_),
    .Y(_02984_));
 sky130_fd_sc_hd__a31o_1 _16469_ (.A1(_02966_),
    .A2(net1509),
    .A3(_02944_),
    .B1(_02984_),
    .X(_00361_));
 sky130_fd_sc_hd__nand2_1 _16470_ (.A(_02931_),
    .B(net2872),
    .Y(_02985_));
 sky130_fd_sc_hd__a22o_1 _16471_ (.A1(_02948_),
    .A2(_10624_),
    .B1(_02942_),
    .B2(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__inv_2 _16472_ (.A(_02986_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_1 _16473_ (.A(_02931_),
    .B(net3014),
    .Y(_02987_));
 sky130_fd_sc_hd__a22o_1 _16474_ (.A1(_02948_),
    .A2(_02928_),
    .B1(_02942_),
    .B2(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__inv_2 _16475_ (.A(_02988_),
    .Y(_00363_));
 sky130_fd_sc_hd__and3_1 _16476_ (.A(_02939_),
    .B(_10848_),
    .C(_02854_),
    .X(_02989_));
 sky130_fd_sc_hd__a31o_1 _16477_ (.A1(_02943_),
    .A2(_02751_),
    .A3(net2331),
    .B1(_02989_),
    .X(_00364_));
 sky130_fd_sc_hd__and3_1 _16478_ (.A(_02939_),
    .B(_11426_),
    .C(_02854_),
    .X(_02990_));
 sky130_fd_sc_hd__a31o_1 _16479_ (.A1(_02943_),
    .A2(_02751_),
    .A3(net2511),
    .B1(_02990_),
    .X(_00365_));
 sky130_fd_sc_hd__nand2_1 _16480_ (.A(_02935_),
    .B(net3806),
    .Y(_02991_));
 sky130_fd_sc_hd__buf_8 _16481_ (.A(_09297_),
    .X(_02992_));
 sky130_fd_sc_hd__o2bb2a_1 _16482_ (.A1_N(_02991_),
    .A2_N(_02943_),
    .B1(_02992_),
    .B2(_02940_),
    .X(_00366_));
 sky130_fd_sc_hd__nor2_1 _16483_ (.A(_09300_),
    .B(_02944_),
    .Y(_02993_));
 sky130_fd_sc_hd__a31o_1 _16484_ (.A1(_02966_),
    .A2(net1123),
    .A3(_02944_),
    .B1(_02993_),
    .X(_00367_));
 sky130_fd_sc_hd__nor2_4 _16485_ (.A(_02938_),
    .B(_10292_),
    .Y(_02994_));
 sky130_fd_sc_hd__nand2_4 _16486_ (.A(_02994_),
    .B(_10413_),
    .Y(_02995_));
 sky130_fd_sc_hd__buf_4 _16487_ (.A(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__nand2_1 _16488_ (.A(_02831_),
    .B(net3971),
    .Y(_02997_));
 sky130_fd_sc_hd__inv_2 _16489_ (.A(_02938_),
    .Y(_02998_));
 sky130_fd_sc_hd__and3_1 _16490_ (.A(_10291_),
    .B(_02998_),
    .C(_08725_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_4 _16491_ (.A(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__a22o_1 _16492_ (.A1(_02996_),
    .A2(_02997_),
    .B1(_09451_),
    .B2(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__inv_2 _16493_ (.A(_03001_),
    .Y(_00344_));
 sky130_fd_sc_hd__buf_4 _16494_ (.A(_02995_),
    .X(_03002_));
 sky130_fd_sc_hd__nor2_1 _16495_ (.A(_10746_),
    .B(_02996_),
    .Y(_03003_));
 sky130_fd_sc_hd__a31o_1 _16496_ (.A1(_02966_),
    .A2(net749),
    .A3(_03002_),
    .B1(_03003_),
    .X(_00345_));
 sky130_fd_sc_hd__nor2_1 _16497_ (.A(_10698_),
    .B(_02996_),
    .Y(_03004_));
 sky130_fd_sc_hd__a31o_1 _16498_ (.A1(_02966_),
    .A2(net1237),
    .A3(_03002_),
    .B1(_03004_),
    .X(_00346_));
 sky130_fd_sc_hd__and3_1 _16499_ (.A(_02994_),
    .B(_11040_),
    .C(_02854_),
    .X(_03005_));
 sky130_fd_sc_hd__a31o_1 _16500_ (.A1(_02966_),
    .A2(net1723),
    .A3(_03002_),
    .B1(_03005_),
    .X(_00347_));
 sky130_fd_sc_hd__clkbuf_4 _16501_ (.A(_11219_),
    .X(_03006_));
 sky130_fd_sc_hd__and3_1 _16502_ (.A(_02994_),
    .B(_10587_),
    .C(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__a31o_1 _16503_ (.A1(_02966_),
    .A2(net1635),
    .A3(_03002_),
    .B1(_03007_),
    .X(_00348_));
 sky130_fd_sc_hd__and3_1 _16504_ (.A(_02994_),
    .B(_11391_),
    .C(_03006_),
    .X(_03008_));
 sky130_fd_sc_hd__a31o_1 _16505_ (.A1(_02966_),
    .A2(net651),
    .A3(_03002_),
    .B1(_03008_),
    .X(_00349_));
 sky130_fd_sc_hd__nor2_1 _16506_ (.A(_10872_),
    .B(_02996_),
    .Y(_03009_));
 sky130_fd_sc_hd__a31o_1 _16507_ (.A1(_02966_),
    .A2(net621),
    .A3(_03002_),
    .B1(_03009_),
    .X(_00350_));
 sky130_fd_sc_hd__nand2_1 _16508_ (.A(_02831_),
    .B(net4197),
    .Y(_03010_));
 sky130_fd_sc_hd__a22o_1 _16509_ (.A1(_02995_),
    .A2(_03010_),
    .B1(_03000_),
    .B2(_09212_),
    .X(_03011_));
 sky130_fd_sc_hd__inv_2 _16510_ (.A(_03011_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _16511_ (.A(_02831_),
    .B(net4213),
    .Y(_03012_));
 sky130_fd_sc_hd__a22o_1 _16512_ (.A1(_02995_),
    .A2(_03012_),
    .B1(_03000_),
    .B2(_09531_),
    .X(_03013_));
 sky130_fd_sc_hd__inv_2 _16513_ (.A(_03013_),
    .Y(_00336_));
 sky130_fd_sc_hd__buf_4 _16514_ (.A(_10930_),
    .X(_03014_));
 sky130_fd_sc_hd__nand2_1 _16515_ (.A(_03014_),
    .B(net4054),
    .Y(_03015_));
 sky130_fd_sc_hd__a22o_1 _16516_ (.A1(_02995_),
    .A2(_03015_),
    .B1(_03000_),
    .B2(_10313_),
    .X(_03016_));
 sky130_fd_sc_hd__inv_2 _16517_ (.A(_03016_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _16518_ (.A(_03014_),
    .B(net3984),
    .Y(_03017_));
 sky130_fd_sc_hd__a22o_1 _16519_ (.A1(_02995_),
    .A2(_03017_),
    .B1(_03000_),
    .B2(_10316_),
    .X(_03018_));
 sky130_fd_sc_hd__inv_2 _16520_ (.A(_03018_),
    .Y(_00338_));
 sky130_fd_sc_hd__nor2_1 _16521_ (.A(_02904_),
    .B(_02996_),
    .Y(_03019_));
 sky130_fd_sc_hd__a31o_1 _16522_ (.A1(_02966_),
    .A2(net1517),
    .A3(_03002_),
    .B1(_03019_),
    .X(_00339_));
 sky130_fd_sc_hd__clkbuf_16 _16523_ (.A(_09232_),
    .X(_03020_));
 sky130_fd_sc_hd__nor2_1 _16524_ (.A(_03020_),
    .B(_02996_),
    .Y(_03021_));
 sky130_fd_sc_hd__a31o_1 _16525_ (.A1(_02966_),
    .A2(net1061),
    .A3(_03002_),
    .B1(_03021_),
    .X(_00340_));
 sky130_fd_sc_hd__nand2_1 _16526_ (.A(_03014_),
    .B(net4158),
    .Y(_03022_));
 sky130_fd_sc_hd__a22o_1 _16527_ (.A1(_02995_),
    .A2(_03022_),
    .B1(_03000_),
    .B2(_09338_),
    .X(_03023_));
 sky130_fd_sc_hd__inv_2 _16528_ (.A(_03023_),
    .Y(_00341_));
 sky130_fd_sc_hd__buf_4 _16529_ (.A(_02772_),
    .X(_03024_));
 sky130_fd_sc_hd__and3_1 _16530_ (.A(_02994_),
    .B(_11291_),
    .C(_03006_),
    .X(_03025_));
 sky130_fd_sc_hd__a31o_1 _16531_ (.A1(_03024_),
    .A2(net2073),
    .A3(_03002_),
    .B1(_03025_),
    .X(_00342_));
 sky130_fd_sc_hd__buf_8 _16532_ (.A(_09242_),
    .X(_03026_));
 sky130_fd_sc_hd__nor2_1 _16533_ (.A(_03026_),
    .B(_02996_),
    .Y(_03027_));
 sky130_fd_sc_hd__a31o_1 _16534_ (.A1(_03024_),
    .A2(net1017),
    .A3(_03002_),
    .B1(_03027_),
    .X(_00343_));
 sky130_fd_sc_hd__nor2_1 _16535_ (.A(_11002_),
    .B(_02996_),
    .Y(_03028_));
 sky130_fd_sc_hd__a31o_1 _16536_ (.A1(_03024_),
    .A2(net679),
    .A3(_03002_),
    .B1(_03028_),
    .X(_00328_));
 sky130_fd_sc_hd__buf_8 _16537_ (.A(net82),
    .X(_03029_));
 sky130_fd_sc_hd__and3_1 _16538_ (.A(_02994_),
    .B(_03029_),
    .C(_03006_),
    .X(_03030_));
 sky130_fd_sc_hd__a31o_1 _16539_ (.A1(_03024_),
    .A2(net413),
    .A3(_03002_),
    .B1(_03030_),
    .X(_00329_));
 sky130_fd_sc_hd__nor2_1 _16540_ (.A(_10669_),
    .B(_02996_),
    .Y(_03031_));
 sky130_fd_sc_hd__a31o_1 _16541_ (.A1(_03024_),
    .A2(net473),
    .A3(_03002_),
    .B1(_03031_),
    .X(_00330_));
 sky130_fd_sc_hd__buf_8 _16542_ (.A(net52),
    .X(_03032_));
 sky130_fd_sc_hd__and3_1 _16543_ (.A(_02994_),
    .B(_03032_),
    .C(_03006_),
    .X(_03033_));
 sky130_fd_sc_hd__a31o_1 _16544_ (.A1(_03024_),
    .A2(net663),
    .A3(_03002_),
    .B1(_03033_),
    .X(_00331_));
 sky130_fd_sc_hd__nor2_1 _16545_ (.A(_11010_),
    .B(_02996_),
    .Y(_03034_));
 sky130_fd_sc_hd__a31o_1 _16546_ (.A1(_03024_),
    .A2(net1515),
    .A3(_03002_),
    .B1(_03034_),
    .X(_00332_));
 sky130_fd_sc_hd__nand2_1 _16547_ (.A(_03014_),
    .B(net4125),
    .Y(_03035_));
 sky130_fd_sc_hd__a22o_1 _16548_ (.A1(_02995_),
    .A2(_03035_),
    .B1(_03000_),
    .B2(_10331_),
    .X(_03036_));
 sky130_fd_sc_hd__inv_2 _16549_ (.A(_03036_),
    .Y(_00333_));
 sky130_fd_sc_hd__and3_1 _16550_ (.A(_02994_),
    .B(_10617_),
    .C(_03006_),
    .X(_03037_));
 sky130_fd_sc_hd__a31o_1 _16551_ (.A1(_03024_),
    .A2(net717),
    .A3(_03002_),
    .B1(_03037_),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_1 _16552_ (.A(_03014_),
    .B(net4123),
    .Y(_03038_));
 sky130_fd_sc_hd__a22o_1 _16553_ (.A1(_02995_),
    .A2(_03038_),
    .B1(_03000_),
    .B2(_10335_),
    .X(_03039_));
 sky130_fd_sc_hd__inv_2 _16554_ (.A(_03039_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _16555_ (.A(_03014_),
    .B(net3999),
    .Y(_03040_));
 sky130_fd_sc_hd__a22o_1 _16556_ (.A1(_02995_),
    .A2(_03040_),
    .B1(_03000_),
    .B2(_09495_),
    .X(_03041_));
 sky130_fd_sc_hd__inv_2 _16557_ (.A(_03041_),
    .Y(_00320_));
 sky130_fd_sc_hd__nor2_1 _16558_ (.A(_10681_),
    .B(_02996_),
    .Y(_03042_));
 sky130_fd_sc_hd__a31o_1 _16559_ (.A1(_03024_),
    .A2(net1568),
    .A3(_02996_),
    .B1(_03042_),
    .X(_00321_));
 sky130_fd_sc_hd__and3_1 _16560_ (.A(_02994_),
    .B(_10728_),
    .C(_03006_),
    .X(_03043_));
 sky130_fd_sc_hd__a31o_1 _16561_ (.A1(_03024_),
    .A2(net857),
    .A3(_02996_),
    .B1(_03043_),
    .X(_00322_));
 sky130_fd_sc_hd__nand2_1 _16562_ (.A(_03014_),
    .B(net4244),
    .Y(_03044_));
 sky130_fd_sc_hd__a22o_1 _16563_ (.A1(_02995_),
    .A2(_03044_),
    .B1(_03000_),
    .B2(_10342_),
    .X(_03045_));
 sky130_fd_sc_hd__inv_2 _16564_ (.A(_03045_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _16565_ (.A(_03014_),
    .B(net4134),
    .Y(_03046_));
 sky130_fd_sc_hd__a22o_1 _16566_ (.A1(_02995_),
    .A2(_03046_),
    .B1(_03000_),
    .B2(_09288_),
    .X(_03047_));
 sky130_fd_sc_hd__inv_2 _16567_ (.A(_03047_),
    .Y(_00324_));
 sky130_fd_sc_hd__and3_1 _16568_ (.A(_02994_),
    .B(_11426_),
    .C(_03006_),
    .X(_03048_));
 sky130_fd_sc_hd__a31o_1 _16569_ (.A1(_03024_),
    .A2(net1393),
    .A3(_02996_),
    .B1(_03048_),
    .X(_00325_));
 sky130_fd_sc_hd__nand2_1 _16570_ (.A(_02931_),
    .B(net3545),
    .Y(_03049_));
 sky130_fd_sc_hd__a22o_1 _16571_ (.A1(_10348_),
    .A2(_02994_),
    .B1(_02996_),
    .B2(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__inv_2 _16572_ (.A(net3546),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _16573_ (.A(_02931_),
    .B(net3599),
    .Y(_03051_));
 sky130_fd_sc_hd__a22o_1 _16574_ (.A1(_09440_),
    .A2(_02994_),
    .B1(_02996_),
    .B2(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__inv_2 _16575_ (.A(net3600),
    .Y(_00327_));
 sky130_fd_sc_hd__nor2_4 _16576_ (.A(_02938_),
    .B(_10356_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2_4 _16577_ (.A(_03053_),
    .B(_09226_),
    .Y(_03054_));
 sky130_fd_sc_hd__buf_4 _16578_ (.A(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__buf_4 _16579_ (.A(_03054_),
    .X(_03056_));
 sky130_fd_sc_hd__nor2_1 _16580_ (.A(_11210_),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__a31o_1 _16581_ (.A1(_03024_),
    .A2(net1185),
    .A3(_03055_),
    .B1(_03057_),
    .X(_00312_));
 sky130_fd_sc_hd__nor2_1 _16582_ (.A(_10746_),
    .B(_03056_),
    .Y(_03058_));
 sky130_fd_sc_hd__a31o_1 _16583_ (.A1(_03024_),
    .A2(net827),
    .A3(_03055_),
    .B1(_03058_),
    .X(_00313_));
 sky130_fd_sc_hd__nor2_1 _16584_ (.A(_10698_),
    .B(_03056_),
    .Y(_03059_));
 sky130_fd_sc_hd__a31o_1 _16585_ (.A1(_03024_),
    .A2(net1437),
    .A3(_03055_),
    .B1(_03059_),
    .X(_00314_));
 sky130_fd_sc_hd__and3_1 _16586_ (.A(_03053_),
    .B(_11040_),
    .C(_03006_),
    .X(_03060_));
 sky130_fd_sc_hd__a31o_1 _16587_ (.A1(_03024_),
    .A2(net741),
    .A3(_03055_),
    .B1(_03060_),
    .X(_00315_));
 sky130_fd_sc_hd__and3_1 _16588_ (.A(_03053_),
    .B(_10586_),
    .C(_03006_),
    .X(_03061_));
 sky130_fd_sc_hd__a31o_1 _16589_ (.A1(_03024_),
    .A2(net629),
    .A3(_03055_),
    .B1(_03061_),
    .X(_00316_));
 sky130_fd_sc_hd__nand2_1 _16590_ (.A(_03014_),
    .B(net4146),
    .Y(_03062_));
 sky130_fd_sc_hd__and3_2 _16591_ (.A(_10355_),
    .B(_02998_),
    .C(_08778_),
    .X(_03063_));
 sky130_fd_sc_hd__a22o_1 _16592_ (.A1(_03054_),
    .A2(_03062_),
    .B1(_03063_),
    .B2(_09205_),
    .X(_03064_));
 sky130_fd_sc_hd__inv_2 _16593_ (.A(_03064_),
    .Y(_00317_));
 sky130_fd_sc_hd__buf_4 _16594_ (.A(_02772_),
    .X(_03065_));
 sky130_fd_sc_hd__nor2_1 _16595_ (.A(_10872_),
    .B(_03056_),
    .Y(_03066_));
 sky130_fd_sc_hd__a31o_1 _16596_ (.A1(_03065_),
    .A2(net1921),
    .A3(_03055_),
    .B1(_03066_),
    .X(_00318_));
 sky130_fd_sc_hd__and3_1 _16597_ (.A(_03053_),
    .B(_10874_),
    .C(_03006_),
    .X(_03067_));
 sky130_fd_sc_hd__a31o_1 _16598_ (.A1(_03065_),
    .A2(net2028),
    .A3(_03055_),
    .B1(_03067_),
    .X(_00319_));
 sky130_fd_sc_hd__nor2_1 _16599_ (.A(_10760_),
    .B(_03056_),
    .Y(_03068_));
 sky130_fd_sc_hd__a31o_1 _16600_ (.A1(_03065_),
    .A2(net1087),
    .A3(_03055_),
    .B1(_03068_),
    .X(_00304_));
 sky130_fd_sc_hd__nand2_1 _16601_ (.A(_03014_),
    .B(net4050),
    .Y(_03069_));
 sky130_fd_sc_hd__a22o_1 _16602_ (.A1(_03054_),
    .A2(_03069_),
    .B1(_03063_),
    .B2(_10313_),
    .X(_03070_));
 sky130_fd_sc_hd__inv_2 _16603_ (.A(_03070_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _16604_ (.A(_03014_),
    .B(net4087),
    .Y(_03071_));
 sky130_fd_sc_hd__a22o_1 _16605_ (.A1(_03054_),
    .A2(_03071_),
    .B1(_03063_),
    .B2(_10316_),
    .X(_03072_));
 sky130_fd_sc_hd__inv_2 _16606_ (.A(_03072_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _16607_ (.A(_03014_),
    .B(net4130),
    .Y(_03073_));
 sky130_fd_sc_hd__a22o_1 _16608_ (.A1(_03054_),
    .A2(_03073_),
    .B1(_03063_),
    .B2(_09589_),
    .X(_03074_));
 sky130_fd_sc_hd__inv_2 _16609_ (.A(_03074_),
    .Y(_00307_));
 sky130_fd_sc_hd__nor2_1 _16610_ (.A(_03020_),
    .B(_03056_),
    .Y(_03075_));
 sky130_fd_sc_hd__a31o_1 _16611_ (.A1(_03065_),
    .A2(net1031),
    .A3(_03055_),
    .B1(_03075_),
    .X(_00308_));
 sky130_fd_sc_hd__nor2_1 _16612_ (.A(_02845_),
    .B(_03056_),
    .Y(_03076_));
 sky130_fd_sc_hd__a31o_1 _16613_ (.A1(_03065_),
    .A2(net791),
    .A3(_03055_),
    .B1(_03076_),
    .X(_00309_));
 sky130_fd_sc_hd__nand2_1 _16614_ (.A(_03014_),
    .B(net4122),
    .Y(_03077_));
 sky130_fd_sc_hd__a22o_1 _16615_ (.A1(_03054_),
    .A2(_03077_),
    .B1(_03063_),
    .B2(_09239_),
    .X(_03078_));
 sky130_fd_sc_hd__inv_2 _16616_ (.A(_03078_),
    .Y(_00310_));
 sky130_fd_sc_hd__nor2_1 _16617_ (.A(_03026_),
    .B(_03056_),
    .Y(_03079_));
 sky130_fd_sc_hd__a31o_1 _16618_ (.A1(_03065_),
    .A2(net1395),
    .A3(_03055_),
    .B1(_03079_),
    .X(_00311_));
 sky130_fd_sc_hd__nor2_1 _16619_ (.A(_11002_),
    .B(_03056_),
    .Y(_03080_));
 sky130_fd_sc_hd__a31o_1 _16620_ (.A1(_03065_),
    .A2(net1834),
    .A3(_03055_),
    .B1(_03080_),
    .X(_00296_));
 sky130_fd_sc_hd__and3_1 _16621_ (.A(_03053_),
    .B(_03029_),
    .C(_03006_),
    .X(_03081_));
 sky130_fd_sc_hd__a31o_1 _16622_ (.A1(_03065_),
    .A2(net577),
    .A3(_03055_),
    .B1(_03081_),
    .X(_00297_));
 sky130_fd_sc_hd__nor2_1 _16623_ (.A(_10669_),
    .B(_03056_),
    .Y(_03082_));
 sky130_fd_sc_hd__a31o_1 _16624_ (.A1(_03065_),
    .A2(net627),
    .A3(_03055_),
    .B1(_03082_),
    .X(_00298_));
 sky130_fd_sc_hd__and3_1 _16625_ (.A(_03053_),
    .B(_03032_),
    .C(_03006_),
    .X(_03083_));
 sky130_fd_sc_hd__a31o_1 _16626_ (.A1(_03065_),
    .A2(net515),
    .A3(_03055_),
    .B1(_03083_),
    .X(_00299_));
 sky130_fd_sc_hd__nor2_1 _16627_ (.A(_11010_),
    .B(_03054_),
    .Y(_03084_));
 sky130_fd_sc_hd__a31o_1 _16628_ (.A1(_03065_),
    .A2(net461),
    .A3(_03055_),
    .B1(_03084_),
    .X(_00300_));
 sky130_fd_sc_hd__nand2_1 _16629_ (.A(_03014_),
    .B(net3916),
    .Y(_03085_));
 sky130_fd_sc_hd__a22o_1 _16630_ (.A1(_03054_),
    .A2(_03085_),
    .B1(_03063_),
    .B2(_10331_),
    .X(_03086_));
 sky130_fd_sc_hd__inv_2 _16631_ (.A(_03086_),
    .Y(_00301_));
 sky130_fd_sc_hd__buf_8 _16632_ (.A(net55),
    .X(_03087_));
 sky130_fd_sc_hd__and3_1 _16633_ (.A(_03053_),
    .B(_03087_),
    .C(_03006_),
    .X(_03088_));
 sky130_fd_sc_hd__a31o_1 _16634_ (.A1(_03065_),
    .A2(net1139),
    .A3(_03056_),
    .B1(_03088_),
    .X(_00302_));
 sky130_fd_sc_hd__nand2_1 _16635_ (.A(_03014_),
    .B(net3959),
    .Y(_03089_));
 sky130_fd_sc_hd__a22o_1 _16636_ (.A1(_03054_),
    .A2(_03089_),
    .B1(_03063_),
    .B2(_10335_),
    .X(_03090_));
 sky130_fd_sc_hd__inv_2 _16637_ (.A(_03090_),
    .Y(_00303_));
 sky130_fd_sc_hd__and3_1 _16638_ (.A(_03053_),
    .B(_10679_),
    .C(_03006_),
    .X(_03091_));
 sky130_fd_sc_hd__a31o_1 _16639_ (.A1(_03065_),
    .A2(net945),
    .A3(_03056_),
    .B1(_03091_),
    .X(_00288_));
 sky130_fd_sc_hd__nor2_1 _16640_ (.A(_10681_),
    .B(_03054_),
    .Y(_03092_));
 sky130_fd_sc_hd__a31o_1 _16641_ (.A1(_03065_),
    .A2(net611),
    .A3(_03056_),
    .B1(_03092_),
    .X(_00289_));
 sky130_fd_sc_hd__and3_1 _16642_ (.A(_03053_),
    .B(_10728_),
    .C(_03006_),
    .X(_03093_));
 sky130_fd_sc_hd__a31o_1 _16643_ (.A1(_03065_),
    .A2(net463),
    .A3(_03056_),
    .B1(_03093_),
    .X(_00290_));
 sky130_fd_sc_hd__nand2_1 _16644_ (.A(_03014_),
    .B(net4010),
    .Y(_03094_));
 sky130_fd_sc_hd__a22o_1 _16645_ (.A1(_03054_),
    .A2(_03094_),
    .B1(_03063_),
    .B2(_10342_),
    .X(_03095_));
 sky130_fd_sc_hd__inv_2 _16646_ (.A(_03095_),
    .Y(_00291_));
 sky130_fd_sc_hd__buf_4 _16647_ (.A(_11219_),
    .X(_03096_));
 sky130_fd_sc_hd__and3_1 _16648_ (.A(_03053_),
    .B(_10848_),
    .C(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__a31o_1 _16649_ (.A1(_03065_),
    .A2(net485),
    .A3(_03056_),
    .B1(_03097_),
    .X(_00292_));
 sky130_fd_sc_hd__clkbuf_8 _16650_ (.A(_02772_),
    .X(_03098_));
 sky130_fd_sc_hd__and3_1 _16651_ (.A(_03053_),
    .B(_11426_),
    .C(_03096_),
    .X(_03099_));
 sky130_fd_sc_hd__a31o_1 _16652_ (.A1(_03098_),
    .A2(net1585),
    .A3(_03056_),
    .B1(_03099_),
    .X(_00293_));
 sky130_fd_sc_hd__buf_4 _16653_ (.A(_11151_),
    .X(_03100_));
 sky130_fd_sc_hd__nand2_1 _16654_ (.A(_03100_),
    .B(net2923),
    .Y(_03101_));
 sky130_fd_sc_hd__a22o_1 _16655_ (.A1(_10348_),
    .A2(_03053_),
    .B1(_03054_),
    .B2(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__inv_2 _16656_ (.A(net2924),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _16657_ (.A(_03100_),
    .B(net2799),
    .Y(_03103_));
 sky130_fd_sc_hd__a22o_1 _16658_ (.A1(_09440_),
    .A2(_03053_),
    .B1(_03054_),
    .B2(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__inv_2 _16659_ (.A(net2800),
    .Y(_00295_));
 sky130_fd_sc_hd__nor2_2 _16660_ (.A(_02938_),
    .B(_10411_),
    .Y(_03105_));
 sky130_fd_sc_hd__inv_2 _16661_ (.A(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nor2_8 _16662_ (.A(_08794_),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__nor2_1 _16663_ (.A(_08728_),
    .B(_03106_),
    .Y(_03108_));
 sky130_fd_sc_hd__inv_2 _16664_ (.A(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__buf_4 _16665_ (.A(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__nand2_1 _16666_ (.A(_03100_),
    .B(net3198),
    .Y(_03111_));
 sky130_fd_sc_hd__a22o_1 _16667_ (.A1(_03107_),
    .A2(_10239_),
    .B1(_03110_),
    .B2(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__inv_2 _16668_ (.A(_03112_),
    .Y(_00280_));
 sky130_fd_sc_hd__buf_4 _16669_ (.A(_03109_),
    .X(_03113_));
 sky130_fd_sc_hd__nor2_1 _16670_ (.A(_10746_),
    .B(_03110_),
    .Y(_03114_));
 sky130_fd_sc_hd__a31o_1 _16671_ (.A1(_03098_),
    .A2(net1227),
    .A3(_03113_),
    .B1(_03114_),
    .X(_00281_));
 sky130_fd_sc_hd__nand2_1 _16672_ (.A(_03100_),
    .B(net3270),
    .Y(_03115_));
 sky130_fd_sc_hd__a22o_1 _16673_ (.A1(_03107_),
    .A2(_09459_),
    .B1(_03110_),
    .B2(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__inv_2 _16674_ (.A(_03116_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _16675_ (.A(_03100_),
    .B(net3597),
    .Y(_03117_));
 sky130_fd_sc_hd__a22o_1 _16676_ (.A1(_03107_),
    .A2(_10983_),
    .B1(_03110_),
    .B2(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__inv_2 _16677_ (.A(_03118_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _16678_ (.A(_03100_),
    .B(net3052),
    .Y(_03119_));
 sky130_fd_sc_hd__a22o_1 _16679_ (.A1(_03107_),
    .A2(_11330_),
    .B1(_03110_),
    .B2(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__inv_2 _16680_ (.A(_03120_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _16681_ (.A(_03100_),
    .B(net3481),
    .Y(_03121_));
 sky130_fd_sc_hd__a22o_1 _16682_ (.A1(_03107_),
    .A2(_10869_),
    .B1(_03110_),
    .B2(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__inv_2 _16683_ (.A(_03122_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _16684_ (.A(_03100_),
    .B(net3442),
    .Y(_03123_));
 sky130_fd_sc_hd__a22o_1 _16685_ (.A1(_03107_),
    .A2(_11105_),
    .B1(_03110_),
    .B2(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__inv_2 _16686_ (.A(_03124_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _16687_ (.A(_03100_),
    .B(net3525),
    .Y(_03125_));
 sky130_fd_sc_hd__a22o_1 _16688_ (.A1(_03107_),
    .A2(_10591_),
    .B1(_03110_),
    .B2(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__inv_2 _16689_ (.A(_03126_),
    .Y(_00287_));
 sky130_fd_sc_hd__nor2_1 _16690_ (.A(_10760_),
    .B(_03110_),
    .Y(_03127_));
 sky130_fd_sc_hd__a31o_1 _16691_ (.A1(_03098_),
    .A2(net435),
    .A3(_03113_),
    .B1(_03127_),
    .X(_00272_));
 sky130_fd_sc_hd__nand2_1 _16692_ (.A(_03100_),
    .B(net3536),
    .Y(_03128_));
 sky130_fd_sc_hd__a22o_1 _16693_ (.A1(_03107_),
    .A2(_02899_),
    .B1(_03110_),
    .B2(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__inv_2 _16694_ (.A(_03129_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _16695_ (.A(_03100_),
    .B(net3115),
    .Y(_03130_));
 sky130_fd_sc_hd__a22o_1 _16696_ (.A1(_03107_),
    .A2(_02963_),
    .B1(_03110_),
    .B2(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__inv_2 _16697_ (.A(_03131_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _16698_ (.A(_03100_),
    .B(net3243),
    .Y(_03132_));
 sky130_fd_sc_hd__a22o_1 _16699_ (.A1(_03107_),
    .A2(_09589_),
    .B1(_03109_),
    .B2(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__inv_2 _16700_ (.A(_03133_),
    .Y(_00275_));
 sky130_fd_sc_hd__nor2_1 _16701_ (.A(_03020_),
    .B(_03110_),
    .Y(_03134_));
 sky130_fd_sc_hd__a31o_1 _16702_ (.A1(_03098_),
    .A2(net2109),
    .A3(_03113_),
    .B1(_03134_),
    .X(_00276_));
 sky130_fd_sc_hd__nor2_1 _16703_ (.A(_02845_),
    .B(_03110_),
    .Y(_03135_));
 sky130_fd_sc_hd__a31o_1 _16704_ (.A1(_03098_),
    .A2(net1850),
    .A3(_03113_),
    .B1(_03135_),
    .X(_00277_));
 sky130_fd_sc_hd__nand2_1 _16705_ (.A(_03100_),
    .B(net3388),
    .Y(_03136_));
 sky130_fd_sc_hd__a22o_1 _16706_ (.A1(_03107_),
    .A2(_10202_),
    .B1(_03109_),
    .B2(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__inv_2 _16707_ (.A(_03137_),
    .Y(_00278_));
 sky130_fd_sc_hd__nor2_1 _16708_ (.A(_03026_),
    .B(_03110_),
    .Y(_03138_));
 sky130_fd_sc_hd__a31o_1 _16709_ (.A1(_03098_),
    .A2(net1355),
    .A3(_03113_),
    .B1(_03138_),
    .X(_00279_));
 sky130_fd_sc_hd__nor2_1 _16710_ (.A(_11002_),
    .B(_03110_),
    .Y(_03139_));
 sky130_fd_sc_hd__a31o_1 _16711_ (.A1(_03098_),
    .A2(net1787),
    .A3(_03113_),
    .B1(_03139_),
    .X(_00256_));
 sky130_fd_sc_hd__and3_1 _16712_ (.A(_03105_),
    .B(_03029_),
    .C(_03096_),
    .X(_03140_));
 sky130_fd_sc_hd__a31o_1 _16713_ (.A1(_03113_),
    .A2(_02751_),
    .A3(net2493),
    .B1(_03140_),
    .X(_00257_));
 sky130_fd_sc_hd__nand2_1 _16714_ (.A(_03100_),
    .B(net3462),
    .Y(_03141_));
 sky130_fd_sc_hd__a22o_1 _16715_ (.A1(_03107_),
    .A2(_09347_),
    .B1(_03109_),
    .B2(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__inv_2 _16716_ (.A(_03142_),
    .Y(_00258_));
 sky130_fd_sc_hd__buf_4 _16717_ (.A(_10645_),
    .X(_03143_));
 sky130_fd_sc_hd__and3_1 _16718_ (.A(_03105_),
    .B(_03032_),
    .C(_03096_),
    .X(_03144_));
 sky130_fd_sc_hd__a31o_1 _16719_ (.A1(_03113_),
    .A2(_03143_),
    .A3(net2483),
    .B1(_03144_),
    .X(_00259_));
 sky130_fd_sc_hd__nand2_1 _16720_ (.A(_03100_),
    .B(net3376),
    .Y(_03145_));
 sky130_fd_sc_hd__a22o_1 _16721_ (.A1(_03107_),
    .A2(_11136_),
    .B1(_03109_),
    .B2(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__inv_2 _16722_ (.A(_03146_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _16723_ (.A(_03100_),
    .B(net3472),
    .Y(_03147_));
 sky130_fd_sc_hd__a22o_1 _16724_ (.A1(_03107_),
    .A2(_02916_),
    .B1(_03109_),
    .B2(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__inv_2 _16725_ (.A(_03148_),
    .Y(_00261_));
 sky130_fd_sc_hd__and3_1 _16726_ (.A(_03105_),
    .B(_03087_),
    .C(_03096_),
    .X(_03149_));
 sky130_fd_sc_hd__a31o_1 _16727_ (.A1(_03113_),
    .A2(_03143_),
    .A3(net573),
    .B1(_03149_),
    .X(_00262_));
 sky130_fd_sc_hd__buf_4 _16728_ (.A(_11151_),
    .X(_03150_));
 sky130_fd_sc_hd__nand2_1 _16729_ (.A(_03150_),
    .B(net2832),
    .Y(_03151_));
 sky130_fd_sc_hd__a22o_1 _16730_ (.A1(_03107_),
    .A2(_02921_),
    .B1(_03109_),
    .B2(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__inv_2 _16731_ (.A(_03152_),
    .Y(_00263_));
 sky130_fd_sc_hd__and3_1 _16732_ (.A(_03105_),
    .B(_10679_),
    .C(_03096_),
    .X(_03153_));
 sky130_fd_sc_hd__a31o_1 _16733_ (.A1(_03113_),
    .A2(_03143_),
    .A3(net2048),
    .B1(_03153_),
    .X(_00248_));
 sky130_fd_sc_hd__nor2_1 _16734_ (.A(_10681_),
    .B(_03110_),
    .Y(_03154_));
 sky130_fd_sc_hd__a31o_1 _16735_ (.A1(_03098_),
    .A2(net1103),
    .A3(_03113_),
    .B1(_03154_),
    .X(_00249_));
 sky130_fd_sc_hd__and3_1 _16736_ (.A(_03105_),
    .B(_10728_),
    .C(_03096_),
    .X(_03155_));
 sky130_fd_sc_hd__a31o_1 _16737_ (.A1(_03113_),
    .A2(_03143_),
    .A3(net2116),
    .B1(_03155_),
    .X(_00250_));
 sky130_fd_sc_hd__nand2_1 _16738_ (.A(_03150_),
    .B(net3742),
    .Y(_03156_));
 sky130_fd_sc_hd__a22o_1 _16739_ (.A1(_03107_),
    .A2(_02928_),
    .B1(_03109_),
    .B2(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__inv_2 _16740_ (.A(_03157_),
    .Y(_00251_));
 sky130_fd_sc_hd__and3_1 _16741_ (.A(_03105_),
    .B(_10848_),
    .C(_03096_),
    .X(_03158_));
 sky130_fd_sc_hd__a31o_1 _16742_ (.A1(_03113_),
    .A2(_03143_),
    .A3(net2496),
    .B1(_03158_),
    .X(_00252_));
 sky130_fd_sc_hd__and3_1 _16743_ (.A(_03105_),
    .B(_11426_),
    .C(_03096_),
    .X(_03159_));
 sky130_fd_sc_hd__a31o_1 _16744_ (.A1(_03113_),
    .A2(_03143_),
    .A3(net2454),
    .B1(_03159_),
    .X(_00253_));
 sky130_fd_sc_hd__nand2_1 _16745_ (.A(_02935_),
    .B(net3611),
    .Y(_03160_));
 sky130_fd_sc_hd__o2bb2a_1 _16746_ (.A1_N(_03160_),
    .A2_N(_03113_),
    .B1(_02992_),
    .B2(_03106_),
    .X(_00254_));
 sky130_fd_sc_hd__nand2_1 _16747_ (.A(_02935_),
    .B(net3640),
    .Y(_03161_));
 sky130_fd_sc_hd__o2bb2a_1 _16748_ (.A1_N(_03161_),
    .A2_N(_03113_),
    .B1(_11316_),
    .B2(_03106_),
    .X(_00255_));
 sky130_fd_sc_hd__inv_2 _16749_ (.A(net3899),
    .Y(_03162_));
 sky130_fd_sc_hd__nor2_8 _16750_ (.A(net2927),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__nand2_4 _16751_ (.A(_03163_),
    .B(_09168_),
    .Y(_03164_));
 sky130_fd_sc_hd__nor2_4 _16752_ (.A(_03164_),
    .B(_10469_),
    .Y(_03165_));
 sky130_fd_sc_hd__nand2_4 _16753_ (.A(_03165_),
    .B(_10413_),
    .Y(_03166_));
 sky130_fd_sc_hd__buf_4 _16754_ (.A(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__buf_4 _16755_ (.A(_03166_),
    .X(_03168_));
 sky130_fd_sc_hd__nor2_1 _16756_ (.A(_11210_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__a31o_1 _16757_ (.A1(_03098_),
    .A2(net2495),
    .A3(_03167_),
    .B1(_03169_),
    .X(_00240_));
 sky130_fd_sc_hd__buf_12 _16758_ (.A(_09184_),
    .X(_03170_));
 sky130_fd_sc_hd__nor2_1 _16759_ (.A(_03170_),
    .B(_03168_),
    .Y(_03171_));
 sky130_fd_sc_hd__a31o_1 _16760_ (.A1(_03098_),
    .A2(net2219),
    .A3(_03167_),
    .B1(_03171_),
    .X(_00241_));
 sky130_fd_sc_hd__nor2_1 _16761_ (.A(_10698_),
    .B(_03166_),
    .Y(_03172_));
 sky130_fd_sc_hd__a31o_1 _16762_ (.A1(_03098_),
    .A2(net1307),
    .A3(_03167_),
    .B1(_03172_),
    .X(_00242_));
 sky130_fd_sc_hd__nand2_1 _16763_ (.A(_02935_),
    .B(net3793),
    .Y(_03173_));
 sky130_fd_sc_hd__nand2_4 _16764_ (.A(_03165_),
    .B(_08778_),
    .Y(_03174_));
 sky130_fd_sc_hd__o2bb2a_1 _16765_ (.A1_N(_03173_),
    .A2_N(_03167_),
    .B1(_10479_),
    .B2(_03174_),
    .X(_00243_));
 sky130_fd_sc_hd__a22o_1 _16766_ (.A1(_09302_),
    .A2(net2754),
    .B1(_03165_),
    .B2(_09227_),
    .X(_03175_));
 sky130_fd_sc_hd__o31a_1 _16767_ (.A1(_09193_),
    .A2(_09321_),
    .A3(_03174_),
    .B1(net2755),
    .X(_00244_));
 sky130_fd_sc_hd__and3_1 _16768_ (.A(_03165_),
    .B(_11391_),
    .C(_03096_),
    .X(_03176_));
 sky130_fd_sc_hd__a31o_1 _16769_ (.A1(_03098_),
    .A2(net1295),
    .A3(_03167_),
    .B1(_03176_),
    .X(_00245_));
 sky130_fd_sc_hd__nor2_1 _16770_ (.A(_10872_),
    .B(_03166_),
    .Y(_03177_));
 sky130_fd_sc_hd__a31o_1 _16771_ (.A1(_03098_),
    .A2(net1465),
    .A3(_03167_),
    .B1(_03177_),
    .X(_00246_));
 sky130_fd_sc_hd__and3_1 _16772_ (.A(_03165_),
    .B(_10874_),
    .C(_03096_),
    .X(_03178_));
 sky130_fd_sc_hd__a31o_1 _16773_ (.A1(_03098_),
    .A2(net2144),
    .A3(_03167_),
    .B1(_03178_),
    .X(_00247_));
 sky130_fd_sc_hd__nor2_1 _16774_ (.A(_10760_),
    .B(_03166_),
    .Y(_03179_));
 sky130_fd_sc_hd__a31o_1 _16775_ (.A1(_03098_),
    .A2(net1467),
    .A3(_03167_),
    .B1(_03179_),
    .X(_00232_));
 sky130_fd_sc_hd__nand2_1 _16776_ (.A(_02935_),
    .B(net3091),
    .Y(_03180_));
 sky130_fd_sc_hd__o2bb2a_1 _16777_ (.A1_N(_03180_),
    .A2_N(_03167_),
    .B1(_10257_),
    .B2(_03174_),
    .X(_00233_));
 sky130_fd_sc_hd__nand2_1 _16778_ (.A(_02935_),
    .B(net4168),
    .Y(_03181_));
 sky130_fd_sc_hd__o2bb2a_1 _16779_ (.A1_N(_03181_),
    .A2_N(_03167_),
    .B1(_10259_),
    .B2(_03174_),
    .X(_00234_));
 sky130_fd_sc_hd__nor2_1 _16780_ (.A(_02904_),
    .B(_03166_),
    .Y(_03182_));
 sky130_fd_sc_hd__a31o_1 _16781_ (.A1(_03098_),
    .A2(net409),
    .A3(_03168_),
    .B1(_03182_),
    .X(_00235_));
 sky130_fd_sc_hd__buf_4 _16782_ (.A(_02772_),
    .X(_03183_));
 sky130_fd_sc_hd__nor2_1 _16783_ (.A(_03020_),
    .B(_03166_),
    .Y(_03184_));
 sky130_fd_sc_hd__a31o_1 _16784_ (.A1(_03183_),
    .A2(net407),
    .A3(_03168_),
    .B1(_03184_),
    .X(_00236_));
 sky130_fd_sc_hd__nand2_1 _16785_ (.A(_02935_),
    .B(net3336),
    .Y(_03185_));
 sky130_fd_sc_hd__o2bb2a_1 _16786_ (.A1_N(_03185_),
    .A2_N(_03167_),
    .B1(_10493_),
    .B2(_03174_),
    .X(_00237_));
 sky130_fd_sc_hd__and3_1 _16787_ (.A(_03165_),
    .B(_11291_),
    .C(_03096_),
    .X(_03186_));
 sky130_fd_sc_hd__a31o_1 _16788_ (.A1(_03183_),
    .A2(net477),
    .A3(_03168_),
    .B1(_03186_),
    .X(_00238_));
 sky130_fd_sc_hd__nor2_1 _16789_ (.A(_03026_),
    .B(_03166_),
    .Y(_03187_));
 sky130_fd_sc_hd__a31o_1 _16790_ (.A1(_03183_),
    .A2(net581),
    .A3(_03168_),
    .B1(_03187_),
    .X(_00239_));
 sky130_fd_sc_hd__nor2_1 _16791_ (.A(_11002_),
    .B(_03166_),
    .Y(_03188_));
 sky130_fd_sc_hd__a31o_1 _16792_ (.A1(_03183_),
    .A2(net919),
    .A3(_03168_),
    .B1(_03188_),
    .X(_00224_));
 sky130_fd_sc_hd__and3_1 _16793_ (.A(_03165_),
    .B(_03029_),
    .C(_03096_),
    .X(_03189_));
 sky130_fd_sc_hd__a31o_1 _16794_ (.A1(_03183_),
    .A2(net917),
    .A3(_03168_),
    .B1(_03189_),
    .X(_00225_));
 sky130_fd_sc_hd__nor2_1 _16795_ (.A(_10669_),
    .B(_03166_),
    .Y(_03190_));
 sky130_fd_sc_hd__a31o_1 _16796_ (.A1(_03183_),
    .A2(net975),
    .A3(_03168_),
    .B1(_03190_),
    .X(_00226_));
 sky130_fd_sc_hd__and3_1 _16797_ (.A(_03165_),
    .B(_03032_),
    .C(_03096_),
    .X(_03191_));
 sky130_fd_sc_hd__a31o_1 _16798_ (.A1(_03183_),
    .A2(net561),
    .A3(_03168_),
    .B1(_03191_),
    .X(_00227_));
 sky130_fd_sc_hd__nand2_1 _16799_ (.A(_02935_),
    .B(net3905),
    .Y(_03192_));
 sky130_fd_sc_hd__o2bb2a_1 _16800_ (.A1_N(_03192_),
    .A2_N(_03167_),
    .B1(_10503_),
    .B2(_03174_),
    .X(_00228_));
 sky130_fd_sc_hd__nand2_1 _16801_ (.A(_02935_),
    .B(net4133),
    .Y(_03193_));
 sky130_fd_sc_hd__o2bb2a_1 _16802_ (.A1_N(_03193_),
    .A2_N(_03167_),
    .B1(_10273_),
    .B2(_03174_),
    .X(_00229_));
 sky130_fd_sc_hd__and3_1 _16803_ (.A(_03165_),
    .B(_03087_),
    .C(_03096_),
    .X(_03194_));
 sky130_fd_sc_hd__a31o_1 _16804_ (.A1(_03183_),
    .A2(net993),
    .A3(_03168_),
    .B1(_03194_),
    .X(_00230_));
 sky130_fd_sc_hd__nand2_1 _16805_ (.A(_02935_),
    .B(net3352),
    .Y(_03195_));
 sky130_fd_sc_hd__o2bb2a_1 _16806_ (.A1_N(_03195_),
    .A2_N(_03167_),
    .B1(_10276_),
    .B2(_03174_),
    .X(_00231_));
 sky130_fd_sc_hd__buf_8 _16807_ (.A(net50),
    .X(_03196_));
 sky130_fd_sc_hd__and3_1 _16808_ (.A(_03165_),
    .B(_03196_),
    .C(_03096_),
    .X(_03197_));
 sky130_fd_sc_hd__a31o_1 _16809_ (.A1(_03183_),
    .A2(net1275),
    .A3(_03168_),
    .B1(_03197_),
    .X(_00216_));
 sky130_fd_sc_hd__nand2_1 _16810_ (.A(_02935_),
    .B(net3931),
    .Y(_03198_));
 sky130_fd_sc_hd__o2bb2a_1 _16811_ (.A1_N(_03198_),
    .A2_N(_03167_),
    .B1(_10727_),
    .B2(_03174_),
    .X(_00217_));
 sky130_fd_sc_hd__buf_8 _16812_ (.A(net72),
    .X(_03199_));
 sky130_fd_sc_hd__clkbuf_4 _16813_ (.A(_11219_),
    .X(_03200_));
 sky130_fd_sc_hd__and3_1 _16814_ (.A(_03165_),
    .B(_03199_),
    .C(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__a31o_1 _16815_ (.A1(_03183_),
    .A2(net1411),
    .A3(_03168_),
    .B1(_03201_),
    .X(_00218_));
 sky130_fd_sc_hd__nand2_1 _16816_ (.A(_02935_),
    .B(net3737),
    .Y(_03202_));
 sky130_fd_sc_hd__o2bb2a_1 _16817_ (.A1_N(_03202_),
    .A2_N(_03167_),
    .B1(_10285_),
    .B2(_03174_),
    .X(_00219_));
 sky130_fd_sc_hd__and3_1 _16818_ (.A(_03165_),
    .B(_10848_),
    .C(_03200_),
    .X(_03203_));
 sky130_fd_sc_hd__a31o_1 _16819_ (.A1(_03183_),
    .A2(net1566),
    .A3(_03168_),
    .B1(_03203_),
    .X(_00220_));
 sky130_fd_sc_hd__and3_1 _16820_ (.A(_03165_),
    .B(_11426_),
    .C(_03200_),
    .X(_03204_));
 sky130_fd_sc_hd__a31o_1 _16821_ (.A1(_03183_),
    .A2(net1988),
    .A3(_03168_),
    .B1(_03204_),
    .X(_00221_));
 sky130_fd_sc_hd__nand2_1 _16822_ (.A(_03150_),
    .B(net3127),
    .Y(_03205_));
 sky130_fd_sc_hd__a22o_1 _16823_ (.A1(_10348_),
    .A2(_03165_),
    .B1(_03166_),
    .B2(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__inv_2 _16824_ (.A(_03206_),
    .Y(_00222_));
 sky130_fd_sc_hd__nor2_1 _16825_ (.A(_09299_),
    .B(_03166_),
    .Y(_03207_));
 sky130_fd_sc_hd__a31o_1 _16826_ (.A1(_03183_),
    .A2(net785),
    .A3(_03168_),
    .B1(_03207_),
    .X(_00223_));
 sky130_fd_sc_hd__nor2_2 _16827_ (.A(_03164_),
    .B(_10292_),
    .Y(_03208_));
 sky130_fd_sc_hd__inv_2 _16828_ (.A(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__nor2_4 _16829_ (.A(_08797_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__nor2_1 _16830_ (.A(_09166_),
    .B(_03209_),
    .Y(_03211_));
 sky130_fd_sc_hd__inv_2 _16831_ (.A(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__buf_4 _16832_ (.A(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__nand2_1 _16833_ (.A(_03150_),
    .B(net3338),
    .Y(_03214_));
 sky130_fd_sc_hd__a22o_1 _16834_ (.A1(_03210_),
    .A2(_10239_),
    .B1(_03213_),
    .B2(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__inv_2 _16835_ (.A(_03215_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _16836_ (.A(_03150_),
    .B(net3516),
    .Y(_03216_));
 sky130_fd_sc_hd__a22o_1 _16837_ (.A1(_03210_),
    .A2(_09314_),
    .B1(_03213_),
    .B2(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__inv_2 _16838_ (.A(_03217_),
    .Y(_00209_));
 sky130_fd_sc_hd__buf_4 _16839_ (.A(_03212_),
    .X(_03218_));
 sky130_fd_sc_hd__buf_12 _16840_ (.A(_09187_),
    .X(_03219_));
 sky130_fd_sc_hd__nor2_1 _16841_ (.A(_03219_),
    .B(_03213_),
    .Y(_03220_));
 sky130_fd_sc_hd__a31o_1 _16842_ (.A1(_03183_),
    .A2(net1793),
    .A3(_03218_),
    .B1(_03220_),
    .X(_00210_));
 sky130_fd_sc_hd__and3_1 _16843_ (.A(_03208_),
    .B(_11040_),
    .C(_03200_),
    .X(_03221_));
 sky130_fd_sc_hd__a31o_1 _16844_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net2174),
    .B1(_03221_),
    .X(_00211_));
 sky130_fd_sc_hd__and3_1 _16845_ (.A(_03208_),
    .B(_10586_),
    .C(_03200_),
    .X(_03222_));
 sky130_fd_sc_hd__a31o_1 _16846_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net1633),
    .B1(_03222_),
    .X(_00212_));
 sky130_fd_sc_hd__and3_1 _16847_ (.A(_03208_),
    .B(_11391_),
    .C(_03200_),
    .X(_03223_));
 sky130_fd_sc_hd__a31o_1 _16848_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net1657),
    .B1(_03223_),
    .X(_00213_));
 sky130_fd_sc_hd__nand2_1 _16849_ (.A(_03150_),
    .B(net3086),
    .Y(_03224_));
 sky130_fd_sc_hd__a22o_1 _16850_ (.A1(_03210_),
    .A2(_11105_),
    .B1(_03213_),
    .B2(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__inv_2 _16851_ (.A(_03225_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _16852_ (.A(_03150_),
    .B(net3429),
    .Y(_03226_));
 sky130_fd_sc_hd__a22o_1 _16853_ (.A1(_03210_),
    .A2(_10591_),
    .B1(_03213_),
    .B2(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__inv_2 _16854_ (.A(_03227_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _16855_ (.A(_03150_),
    .B(net2945),
    .Y(_03228_));
 sky130_fd_sc_hd__a22o_1 _16856_ (.A1(_03210_),
    .A2(_09530_),
    .B1(_03212_),
    .B2(_03228_),
    .X(_03229_));
 sky130_fd_sc_hd__inv_2 _16857_ (.A(_03229_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _16858_ (.A(_03150_),
    .B(net3667),
    .Y(_03230_));
 sky130_fd_sc_hd__a22o_1 _16859_ (.A1(_03210_),
    .A2(_02899_),
    .B1(_03212_),
    .B2(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__inv_2 _16860_ (.A(_03231_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _16861_ (.A(_03150_),
    .B(net3617),
    .Y(_03232_));
 sky130_fd_sc_hd__a22o_1 _16862_ (.A1(_03210_),
    .A2(_02963_),
    .B1(_03212_),
    .B2(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__inv_2 _16863_ (.A(_03233_),
    .Y(_00202_));
 sky130_fd_sc_hd__nor2_1 _16864_ (.A(_02904_),
    .B(_03213_),
    .Y(_03234_));
 sky130_fd_sc_hd__a31o_1 _16865_ (.A1(_03183_),
    .A2(net735),
    .A3(_03218_),
    .B1(_03234_),
    .X(_00203_));
 sky130_fd_sc_hd__nor2_1 _16866_ (.A(_03020_),
    .B(_03213_),
    .Y(_03235_));
 sky130_fd_sc_hd__a31o_1 _16867_ (.A1(_03183_),
    .A2(net1840),
    .A3(_03218_),
    .B1(_03235_),
    .X(_00204_));
 sky130_fd_sc_hd__clkbuf_8 _16868_ (.A(_02772_),
    .X(_03236_));
 sky130_fd_sc_hd__nor2_1 _16869_ (.A(_02845_),
    .B(_03213_),
    .Y(_03237_));
 sky130_fd_sc_hd__a31o_1 _16870_ (.A1(_03236_),
    .A2(net1896),
    .A3(_03218_),
    .B1(_03237_),
    .X(_00205_));
 sky130_fd_sc_hd__nand2_1 _16871_ (.A(_03150_),
    .B(net3501),
    .Y(_03238_));
 sky130_fd_sc_hd__a22o_1 _16872_ (.A1(_03210_),
    .A2(_10202_),
    .B1(_03212_),
    .B2(_03238_),
    .X(_03239_));
 sky130_fd_sc_hd__inv_2 _16873_ (.A(_03239_),
    .Y(_00206_));
 sky130_fd_sc_hd__nor2_1 _16874_ (.A(_03026_),
    .B(_03213_),
    .Y(_03240_));
 sky130_fd_sc_hd__a31o_1 _16875_ (.A1(_03236_),
    .A2(net2011),
    .A3(_03218_),
    .B1(_03240_),
    .X(_00207_));
 sky130_fd_sc_hd__nor2_1 _16876_ (.A(_11002_),
    .B(_03213_),
    .Y(_03241_));
 sky130_fd_sc_hd__a31o_1 _16877_ (.A1(_03236_),
    .A2(net1806),
    .A3(_03218_),
    .B1(_03241_),
    .X(_00192_));
 sky130_fd_sc_hd__and3_1 _16878_ (.A(_03208_),
    .B(_03029_),
    .C(_03200_),
    .X(_03242_));
 sky130_fd_sc_hd__a31o_1 _16879_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net2030),
    .B1(_03242_),
    .X(_00193_));
 sky130_fd_sc_hd__nor2_1 _16880_ (.A(_10669_),
    .B(_03213_),
    .Y(_03243_));
 sky130_fd_sc_hd__a31o_1 _16881_ (.A1(_03236_),
    .A2(net415),
    .A3(_03213_),
    .B1(_03243_),
    .X(_00194_));
 sky130_fd_sc_hd__nand2_1 _16882_ (.A(_03150_),
    .B(net3003),
    .Y(_03244_));
 sky130_fd_sc_hd__a22o_1 _16883_ (.A1(_03210_),
    .A2(_09256_),
    .B1(_03212_),
    .B2(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__inv_2 _16884_ (.A(_03245_),
    .Y(_00195_));
 sky130_fd_sc_hd__nor2_1 _16885_ (.A(_11010_),
    .B(_03213_),
    .Y(_03246_));
 sky130_fd_sc_hd__a31o_1 _16886_ (.A1(_03236_),
    .A2(net489),
    .A3(_03213_),
    .B1(_03246_),
    .X(_00196_));
 sky130_fd_sc_hd__nand2_1 _16887_ (.A(_03150_),
    .B(net3060),
    .Y(_03247_));
 sky130_fd_sc_hd__a22o_1 _16888_ (.A1(_03210_),
    .A2(_02916_),
    .B1(_03212_),
    .B2(_03247_),
    .X(_03248_));
 sky130_fd_sc_hd__inv_2 _16889_ (.A(_03248_),
    .Y(_00197_));
 sky130_fd_sc_hd__and3_1 _16890_ (.A(_03208_),
    .B(_03087_),
    .C(_03200_),
    .X(_03249_));
 sky130_fd_sc_hd__a31o_1 _16891_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net1445),
    .B1(_03249_),
    .X(_00198_));
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(_03150_),
    .B(net3048),
    .Y(_03250_));
 sky130_fd_sc_hd__a22o_1 _16893_ (.A1(_03210_),
    .A2(_02921_),
    .B1(_03212_),
    .B2(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__inv_2 _16894_ (.A(_03251_),
    .Y(_00199_));
 sky130_fd_sc_hd__and3_1 _16895_ (.A(_03208_),
    .B(_03196_),
    .C(_03200_),
    .X(_03252_));
 sky130_fd_sc_hd__a31o_1 _16896_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net2313),
    .B1(_03252_),
    .X(_00184_));
 sky130_fd_sc_hd__nand2_1 _16897_ (.A(_03150_),
    .B(net3488),
    .Y(_03253_));
 sky130_fd_sc_hd__a22o_1 _16898_ (.A1(_03210_),
    .A2(_09365_),
    .B1(_03212_),
    .B2(_03253_),
    .X(_03254_));
 sky130_fd_sc_hd__inv_2 _16899_ (.A(_03254_),
    .Y(_00185_));
 sky130_fd_sc_hd__and3_1 _16900_ (.A(_03208_),
    .B(_03199_),
    .C(_03200_),
    .X(_03255_));
 sky130_fd_sc_hd__a31o_1 _16901_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net2150),
    .B1(_03255_),
    .X(_00186_));
 sky130_fd_sc_hd__nand2_1 _16902_ (.A(_03150_),
    .B(net3574),
    .Y(_03256_));
 sky130_fd_sc_hd__a22o_1 _16903_ (.A1(_03210_),
    .A2(_02928_),
    .B1(_03212_),
    .B2(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__inv_2 _16904_ (.A(_03257_),
    .Y(_00187_));
 sky130_fd_sc_hd__and3_1 _16905_ (.A(_03208_),
    .B(_10848_),
    .C(_03200_),
    .X(_03258_));
 sky130_fd_sc_hd__a31o_1 _16906_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net2007),
    .B1(_03258_),
    .X(_00188_));
 sky130_fd_sc_hd__and3_1 _16907_ (.A(_03208_),
    .B(_11426_),
    .C(_03200_),
    .X(_03259_));
 sky130_fd_sc_hd__a31o_1 _16908_ (.A1(_03218_),
    .A2(_03143_),
    .A3(net2276),
    .B1(_03259_),
    .X(_00189_));
 sky130_fd_sc_hd__nand2_1 _16909_ (.A(_02935_),
    .B(net3715),
    .Y(_03260_));
 sky130_fd_sc_hd__o2bb2a_1 _16910_ (.A1_N(_03260_),
    .A2_N(_03218_),
    .B1(_02992_),
    .B2(_03209_),
    .X(_00190_));
 sky130_fd_sc_hd__nor2_1 _16911_ (.A(_09299_),
    .B(_03213_),
    .Y(_03261_));
 sky130_fd_sc_hd__a31o_1 _16912_ (.A1(_03236_),
    .A2(net693),
    .A3(_03213_),
    .B1(_03261_),
    .X(_00191_));
 sky130_fd_sc_hd__nor2_4 _16913_ (.A(_03164_),
    .B(_10356_),
    .Y(_03262_));
 sky130_fd_sc_hd__inv_2 _16914_ (.A(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_1 _16915_ (.A(_09625_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__inv_2 _16916_ (.A(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__buf_4 _16917_ (.A(_03265_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_4 _16918_ (.A(_03265_),
    .X(_03267_));
 sky130_fd_sc_hd__nor2_1 _16919_ (.A(_11210_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__a31o_1 _16920_ (.A1(_03236_),
    .A2(net2397),
    .A3(_03266_),
    .B1(_03268_),
    .X(_00168_));
 sky130_fd_sc_hd__nor2_1 _16921_ (.A(_03170_),
    .B(_03267_),
    .Y(_03269_));
 sky130_fd_sc_hd__a31o_1 _16922_ (.A1(_03236_),
    .A2(net1203),
    .A3(_03266_),
    .B1(_03269_),
    .X(_00169_));
 sky130_fd_sc_hd__nor2_4 _16923_ (.A(_09190_),
    .B(_03263_),
    .Y(_03270_));
 sky130_fd_sc_hd__buf_4 _16924_ (.A(_08775_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_8 _16925_ (.A(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__nand2_1 _16926_ (.A(_03272_),
    .B(net3363),
    .Y(_03273_));
 sky130_fd_sc_hd__a22o_1 _16927_ (.A1(_03270_),
    .A2(_09459_),
    .B1(_03267_),
    .B2(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__inv_2 _16928_ (.A(_03274_),
    .Y(_00170_));
 sky130_fd_sc_hd__and3_1 _16929_ (.A(_03262_),
    .B(_11040_),
    .C(_03200_),
    .X(_03275_));
 sky130_fd_sc_hd__a31o_1 _16930_ (.A1(_03266_),
    .A2(_03143_),
    .A3(net2588),
    .B1(_03275_),
    .X(_00171_));
 sky130_fd_sc_hd__nand2_1 _16931_ (.A(_03272_),
    .B(net2921),
    .Y(_03276_));
 sky130_fd_sc_hd__a22o_1 _16932_ (.A1(_03270_),
    .A2(_11330_),
    .B1(_03267_),
    .B2(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__inv_2 _16933_ (.A(_03277_),
    .Y(_00172_));
 sky130_fd_sc_hd__clkbuf_8 _16934_ (.A(_10645_),
    .X(_03278_));
 sky130_fd_sc_hd__and3_1 _16935_ (.A(_03262_),
    .B(_11391_),
    .C(_03200_),
    .X(_03279_));
 sky130_fd_sc_hd__a31o_1 _16936_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net1771),
    .B1(_03279_),
    .X(_00173_));
 sky130_fd_sc_hd__nor2_1 _16937_ (.A(_10872_),
    .B(_03267_),
    .Y(_03280_));
 sky130_fd_sc_hd__a31o_1 _16938_ (.A1(_03236_),
    .A2(net1704),
    .A3(_03266_),
    .B1(_03280_),
    .X(_00174_));
 sky130_fd_sc_hd__and3_1 _16939_ (.A(_03262_),
    .B(_10874_),
    .C(_03200_),
    .X(_03281_));
 sky130_fd_sc_hd__a31o_1 _16940_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net2567),
    .B1(_03281_),
    .X(_00175_));
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(_03272_),
    .B(net3294),
    .Y(_03282_));
 sky130_fd_sc_hd__a22o_1 _16942_ (.A1(_03270_),
    .A2(net135),
    .B1(_03267_),
    .B2(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__inv_2 _16943_ (.A(_03283_),
    .Y(_00160_));
 sky130_fd_sc_hd__nand2_1 _16944_ (.A(_03272_),
    .B(net3055),
    .Y(_03284_));
 sky130_fd_sc_hd__a22o_1 _16945_ (.A1(_03270_),
    .A2(_02899_),
    .B1(_03267_),
    .B2(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__inv_2 _16946_ (.A(_03285_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _16947_ (.A(_03272_),
    .B(net2913),
    .Y(_03286_));
 sky130_fd_sc_hd__a22o_1 _16948_ (.A1(_03270_),
    .A2(_02963_),
    .B1(_03265_),
    .B2(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__inv_2 _16949_ (.A(_03287_),
    .Y(_00162_));
 sky130_fd_sc_hd__nor2_1 _16950_ (.A(_02904_),
    .B(_03267_),
    .Y(_03288_));
 sky130_fd_sc_hd__a31o_1 _16951_ (.A1(_03236_),
    .A2(net1853),
    .A3(_03266_),
    .B1(_03288_),
    .X(_00163_));
 sky130_fd_sc_hd__nor2_1 _16952_ (.A(_03020_),
    .B(_03267_),
    .Y(_03289_));
 sky130_fd_sc_hd__a31o_1 _16953_ (.A1(_03236_),
    .A2(net2470),
    .A3(_03267_),
    .B1(_03289_),
    .X(_00164_));
 sky130_fd_sc_hd__nor2_1 _16954_ (.A(_02845_),
    .B(_03267_),
    .Y(_03290_));
 sky130_fd_sc_hd__a31o_1 _16955_ (.A1(_03236_),
    .A2(net2334),
    .A3(_03267_),
    .B1(_03290_),
    .X(_00165_));
 sky130_fd_sc_hd__and3_1 _16956_ (.A(_03262_),
    .B(_11291_),
    .C(_03200_),
    .X(_03291_));
 sky130_fd_sc_hd__a31o_1 _16957_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net2362),
    .B1(_03291_),
    .X(_00166_));
 sky130_fd_sc_hd__nand2_1 _16958_ (.A(_03272_),
    .B(net3411),
    .Y(_03292_));
 sky130_fd_sc_hd__a22o_1 _16959_ (.A1(_03270_),
    .A2(_09768_),
    .B1(_03265_),
    .B2(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__inv_2 _16960_ (.A(_03293_),
    .Y(_00167_));
 sky130_fd_sc_hd__buf_12 _16961_ (.A(_09245_),
    .X(_03294_));
 sky130_fd_sc_hd__nor2_1 _16962_ (.A(_03294_),
    .B(_03267_),
    .Y(_03295_));
 sky130_fd_sc_hd__a31o_1 _16963_ (.A1(_03236_),
    .A2(net1791),
    .A3(_03267_),
    .B1(_03295_),
    .X(_00152_));
 sky130_fd_sc_hd__buf_4 _16964_ (.A(_11219_),
    .X(_03296_));
 sky130_fd_sc_hd__and3_1 _16965_ (.A(_03262_),
    .B(_03029_),
    .C(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__a31o_1 _16966_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net2217),
    .B1(_03297_),
    .X(_00153_));
 sky130_fd_sc_hd__nand2_1 _16967_ (.A(_03272_),
    .B(net3309),
    .Y(_03298_));
 sky130_fd_sc_hd__a22o_1 _16968_ (.A1(_03270_),
    .A2(_09347_),
    .B1(_03265_),
    .B2(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__inv_2 _16969_ (.A(_03299_),
    .Y(_00154_));
 sky130_fd_sc_hd__and3_1 _16970_ (.A(_03262_),
    .B(_03032_),
    .C(_03296_),
    .X(_03300_));
 sky130_fd_sc_hd__a31o_1 _16971_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net2285),
    .B1(_03300_),
    .X(_00155_));
 sky130_fd_sc_hd__nand2_1 _16972_ (.A(_03272_),
    .B(net3461),
    .Y(_03301_));
 sky130_fd_sc_hd__a22o_1 _16973_ (.A1(_03270_),
    .A2(_11136_),
    .B1(_03265_),
    .B2(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__inv_2 _16974_ (.A(_03302_),
    .Y(_00156_));
 sky130_fd_sc_hd__nand2_1 _16975_ (.A(_03272_),
    .B(net3085),
    .Y(_03303_));
 sky130_fd_sc_hd__a22o_1 _16976_ (.A1(_03270_),
    .A2(_02916_),
    .B1(_03265_),
    .B2(_03303_),
    .X(_03304_));
 sky130_fd_sc_hd__inv_2 _16977_ (.A(_03304_),
    .Y(_00157_));
 sky130_fd_sc_hd__and3_1 _16978_ (.A(_03262_),
    .B(_03087_),
    .C(_03296_),
    .X(_03305_));
 sky130_fd_sc_hd__a31o_1 _16979_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net1667),
    .B1(_03305_),
    .X(_00158_));
 sky130_fd_sc_hd__nand2_1 _16980_ (.A(_03272_),
    .B(net3316),
    .Y(_03306_));
 sky130_fd_sc_hd__a22o_1 _16981_ (.A1(_03270_),
    .A2(_02921_),
    .B1(_03265_),
    .B2(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__inv_2 _16982_ (.A(_03307_),
    .Y(_00159_));
 sky130_fd_sc_hd__and3_1 _16983_ (.A(_03262_),
    .B(_03196_),
    .C(_03296_),
    .X(_03308_));
 sky130_fd_sc_hd__a31o_1 _16984_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net2005),
    .B1(_03308_),
    .X(_00144_));
 sky130_fd_sc_hd__nor2_1 _16985_ (.A(_10681_),
    .B(_03267_),
    .Y(_03309_));
 sky130_fd_sc_hd__a31o_1 _16986_ (.A1(_03236_),
    .A2(net1709),
    .A3(_03267_),
    .B1(_03309_),
    .X(_00145_));
 sky130_fd_sc_hd__nand2_1 _16987_ (.A(_03272_),
    .B(net3304),
    .Y(_03310_));
 sky130_fd_sc_hd__a22o_1 _16988_ (.A1(_03270_),
    .A2(_10624_),
    .B1(_03265_),
    .B2(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__inv_2 _16989_ (.A(_03311_),
    .Y(_00146_));
 sky130_fd_sc_hd__nand2_1 _16990_ (.A(_03272_),
    .B(net3099),
    .Y(_03312_));
 sky130_fd_sc_hd__a22o_1 _16991_ (.A1(_03270_),
    .A2(_02928_),
    .B1(_03265_),
    .B2(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__inv_2 _16992_ (.A(_03313_),
    .Y(_00147_));
 sky130_fd_sc_hd__and3_1 _16993_ (.A(_03262_),
    .B(_10848_),
    .C(_03296_),
    .X(_03314_));
 sky130_fd_sc_hd__a31o_1 _16994_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net1765),
    .B1(_03314_),
    .X(_00148_));
 sky130_fd_sc_hd__and3_1 _16995_ (.A(_03262_),
    .B(_11426_),
    .C(_03296_),
    .X(_03315_));
 sky130_fd_sc_hd__a31o_1 _16996_ (.A1(_03266_),
    .A2(_03278_),
    .A3(net1862),
    .B1(_03315_),
    .X(_00149_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(_02935_),
    .B(net3767),
    .Y(_03316_));
 sky130_fd_sc_hd__o2bb2a_1 _16998_ (.A1_N(_03316_),
    .A2_N(_03266_),
    .B1(_02992_),
    .B2(_03263_),
    .X(_00150_));
 sky130_fd_sc_hd__buf_8 _16999_ (.A(_09375_),
    .X(_03317_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_03317_),
    .B(net3577),
    .Y(_03318_));
 sky130_fd_sc_hd__o2bb2a_1 _17001_ (.A1_N(_03318_),
    .A2_N(_03266_),
    .B1(_11316_),
    .B2(_03263_),
    .X(_00151_));
 sky130_fd_sc_hd__nor2_1 _17002_ (.A(_03164_),
    .B(_10411_),
    .Y(_03319_));
 sky130_fd_sc_hd__inv_2 _17003_ (.A(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__nor2_4 _17004_ (.A(_08794_),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__buf_4 _17005_ (.A(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__nor2_1 _17006_ (.A(_09625_),
    .B(_03320_),
    .Y(_03323_));
 sky130_fd_sc_hd__inv_2 _17007_ (.A(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__buf_4 _17008_ (.A(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__nand2_1 _17009_ (.A(_03272_),
    .B(net2844),
    .Y(_03326_));
 sky130_fd_sc_hd__a22o_1 _17010_ (.A1(_03322_),
    .A2(_10239_),
    .B1(_03325_),
    .B2(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__inv_2 _17011_ (.A(_03327_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(_03272_),
    .B(net3570),
    .Y(_03328_));
 sky130_fd_sc_hd__a22o_1 _17013_ (.A1(_03322_),
    .A2(_09314_),
    .B1(_03325_),
    .B2(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__inv_2 _17014_ (.A(_03329_),
    .Y(_00137_));
 sky130_fd_sc_hd__nand2_1 _17015_ (.A(_03272_),
    .B(net3230),
    .Y(_03330_));
 sky130_fd_sc_hd__a22o_1 _17016_ (.A1(_03322_),
    .A2(_09459_),
    .B1(_03325_),
    .B2(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__inv_2 _17017_ (.A(_03331_),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(_03272_),
    .B(net3157),
    .Y(_03332_));
 sky130_fd_sc_hd__a22o_1 _17019_ (.A1(_03322_),
    .A2(_10983_),
    .B1(_03325_),
    .B2(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__inv_2 _17020_ (.A(_03333_),
    .Y(_00139_));
 sky130_fd_sc_hd__buf_4 _17021_ (.A(_03271_),
    .X(_03334_));
 sky130_fd_sc_hd__nand2_1 _17022_ (.A(_03334_),
    .B(net2964),
    .Y(_03335_));
 sky130_fd_sc_hd__a22o_1 _17023_ (.A1(_03322_),
    .A2(_11330_),
    .B1(_03325_),
    .B2(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__inv_2 _17024_ (.A(_03336_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand2_1 _17025_ (.A(_03334_),
    .B(net3042),
    .Y(_03337_));
 sky130_fd_sc_hd__a22o_1 _17026_ (.A1(_03322_),
    .A2(_10869_),
    .B1(_03325_),
    .B2(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__inv_2 _17027_ (.A(_03338_),
    .Y(_00141_));
 sky130_fd_sc_hd__nand2_1 _17028_ (.A(_03334_),
    .B(net3083),
    .Y(_03339_));
 sky130_fd_sc_hd__a22o_1 _17029_ (.A1(_03322_),
    .A2(_11105_),
    .B1(_03325_),
    .B2(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__inv_2 _17030_ (.A(_03340_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _17031_ (.A(_03334_),
    .B(net2849),
    .Y(_03341_));
 sky130_fd_sc_hd__a22o_1 _17032_ (.A1(_03322_),
    .A2(_10591_),
    .B1(_03325_),
    .B2(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__inv_2 _17033_ (.A(_03342_),
    .Y(_00143_));
 sky130_fd_sc_hd__nand2_1 _17034_ (.A(_03334_),
    .B(net3094),
    .Y(_03343_));
 sky130_fd_sc_hd__a22o_1 _17035_ (.A1(_03322_),
    .A2(net135),
    .B1(_03325_),
    .B2(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__inv_2 _17036_ (.A(_03344_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _17037_ (.A(_03334_),
    .B(net2969),
    .Y(_03345_));
 sky130_fd_sc_hd__a22o_1 _17038_ (.A1(_03322_),
    .A2(_02899_),
    .B1(_03325_),
    .B2(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__inv_2 _17039_ (.A(_03346_),
    .Y(_00129_));
 sky130_fd_sc_hd__nand2_1 _17040_ (.A(_03334_),
    .B(net2909),
    .Y(_03347_));
 sky130_fd_sc_hd__a22o_1 _17041_ (.A1(_03322_),
    .A2(_02963_),
    .B1(_03325_),
    .B2(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__inv_2 _17042_ (.A(_03348_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _17043_ (.A(_03334_),
    .B(net3389),
    .Y(_03349_));
 sky130_fd_sc_hd__a22o_1 _17044_ (.A1(_03322_),
    .A2(_09589_),
    .B1(_03325_),
    .B2(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__inv_2 _17045_ (.A(_03350_),
    .Y(_00131_));
 sky130_fd_sc_hd__nand2_1 _17046_ (.A(_03334_),
    .B(net2949),
    .Y(_03351_));
 sky130_fd_sc_hd__a22o_1 _17047_ (.A1(_03322_),
    .A2(_09593_),
    .B1(_03325_),
    .B2(_03351_),
    .X(_03352_));
 sky130_fd_sc_hd__inv_2 _17048_ (.A(_03352_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _17049_ (.A(_03334_),
    .B(net3375),
    .Y(_03353_));
 sky130_fd_sc_hd__a22o_1 _17050_ (.A1(_03322_),
    .A2(_09338_),
    .B1(_03325_),
    .B2(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__inv_2 _17051_ (.A(_03354_),
    .Y(_00133_));
 sky130_fd_sc_hd__buf_4 _17052_ (.A(_03324_),
    .X(_03355_));
 sky130_fd_sc_hd__nand2_1 _17053_ (.A(_03334_),
    .B(net2811),
    .Y(_03356_));
 sky130_fd_sc_hd__a22o_1 _17054_ (.A1(_03322_),
    .A2(_10202_),
    .B1(_03355_),
    .B2(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__inv_2 _17055_ (.A(_03357_),
    .Y(_00134_));
 sky130_fd_sc_hd__nand2_1 _17056_ (.A(_03334_),
    .B(net3024),
    .Y(_03358_));
 sky130_fd_sc_hd__a22o_1 _17057_ (.A1(_03322_),
    .A2(_09768_),
    .B1(_03355_),
    .B2(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__inv_2 _17058_ (.A(_03359_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand2_1 _17059_ (.A(_03334_),
    .B(net2972),
    .Y(_03360_));
 sky130_fd_sc_hd__a22o_1 _17060_ (.A1(_03321_),
    .A2(net138),
    .B1(_03355_),
    .B2(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__inv_2 _17061_ (.A(_03361_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _17062_ (.A(_03334_),
    .B(net3207),
    .Y(_03362_));
 sky130_fd_sc_hd__a22o_1 _17063_ (.A1(_03321_),
    .A2(_09249_),
    .B1(_03355_),
    .B2(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__inv_2 _17064_ (.A(_03363_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_1 _17065_ (.A(_03334_),
    .B(net3480),
    .Y(_03364_));
 sky130_fd_sc_hd__a22o_1 _17066_ (.A1(_03321_),
    .A2(_09347_),
    .B1(_03355_),
    .B2(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__inv_2 _17067_ (.A(_03365_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_1 _17068_ (.A(_03334_),
    .B(net3320),
    .Y(_03366_));
 sky130_fd_sc_hd__a22o_1 _17069_ (.A1(_03321_),
    .A2(_09256_),
    .B1(_03355_),
    .B2(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__inv_2 _17070_ (.A(_03367_),
    .Y(_00123_));
 sky130_fd_sc_hd__clkbuf_8 _17071_ (.A(_03271_),
    .X(_03368_));
 sky130_fd_sc_hd__nand2_1 _17072_ (.A(_03368_),
    .B(net3203),
    .Y(_03369_));
 sky130_fd_sc_hd__a22o_1 _17073_ (.A1(_03321_),
    .A2(_11136_),
    .B1(_03355_),
    .B2(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__inv_2 _17074_ (.A(_03370_),
    .Y(_00124_));
 sky130_fd_sc_hd__nand2_1 _17075_ (.A(_03368_),
    .B(net2992),
    .Y(_03371_));
 sky130_fd_sc_hd__a22o_1 _17076_ (.A1(_03321_),
    .A2(_02916_),
    .B1(_03355_),
    .B2(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__inv_2 _17077_ (.A(_03372_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _17078_ (.A(_03368_),
    .B(net2892),
    .Y(_03373_));
 sky130_fd_sc_hd__a22o_1 _17079_ (.A1(_03321_),
    .A2(_09425_),
    .B1(_03355_),
    .B2(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__inv_2 _17080_ (.A(net2893),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _17081_ (.A(_03368_),
    .B(net2857),
    .Y(_03375_));
 sky130_fd_sc_hd__a22o_1 _17082_ (.A1(_03321_),
    .A2(_02921_),
    .B1(_03355_),
    .B2(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__inv_2 _17083_ (.A(_03376_),
    .Y(_00127_));
 sky130_fd_sc_hd__nand2_1 _17084_ (.A(_03368_),
    .B(net2998),
    .Y(_03377_));
 sky130_fd_sc_hd__a22o_1 _17085_ (.A1(_03321_),
    .A2(net141),
    .B1(_03355_),
    .B2(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__inv_2 _17086_ (.A(_03378_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _17087_ (.A(_03368_),
    .B(net3011),
    .Y(_03379_));
 sky130_fd_sc_hd__a22o_1 _17088_ (.A1(_03321_),
    .A2(_09365_),
    .B1(_03355_),
    .B2(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__inv_2 _17089_ (.A(_03380_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_1 _17090_ (.A(_03368_),
    .B(net3329),
    .Y(_03381_));
 sky130_fd_sc_hd__a22o_1 _17091_ (.A1(_03321_),
    .A2(_10624_),
    .B1(_03355_),
    .B2(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__inv_2 _17092_ (.A(_03382_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _17093_ (.A(_03368_),
    .B(net3161),
    .Y(_03383_));
 sky130_fd_sc_hd__a22o_1 _17094_ (.A1(_03321_),
    .A2(_02928_),
    .B1(_03355_),
    .B2(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__inv_2 _17095_ (.A(_03384_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_1 _17096_ (.A(_03368_),
    .B(net3560),
    .Y(_03385_));
 sky130_fd_sc_hd__a22o_1 _17097_ (.A1(_03321_),
    .A2(net139),
    .B1(_03355_),
    .B2(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__inv_2 _17098_ (.A(_03386_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_1 _17099_ (.A(_03368_),
    .B(net3312),
    .Y(_03387_));
 sky130_fd_sc_hd__a22o_1 _17100_ (.A1(_03321_),
    .A2(net136),
    .B1(_03355_),
    .B2(_03387_),
    .X(_03388_));
 sky130_fd_sc_hd__inv_2 _17101_ (.A(_03388_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_1 _17102_ (.A(_03317_),
    .B(net3810),
    .Y(_03389_));
 sky130_fd_sc_hd__o2bb2a_1 _17103_ (.A1_N(_03389_),
    .A2_N(_03325_),
    .B1(_02992_),
    .B2(_03320_),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_1 _17104_ (.A(_03317_),
    .B(net3763),
    .Y(_03390_));
 sky130_fd_sc_hd__o2bb2a_1 _17105_ (.A1_N(_03390_),
    .A2_N(_03325_),
    .B1(_11316_),
    .B2(_03320_),
    .X(_00119_));
 sky130_fd_sc_hd__nand2_8 _17106_ (.A(_09509_),
    .B(_03163_),
    .Y(_03391_));
 sky130_fd_sc_hd__nor2_4 _17107_ (.A(_10469_),
    .B(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__nand2_4 _17108_ (.A(_03392_),
    .B(_10413_),
    .Y(_03393_));
 sky130_fd_sc_hd__buf_4 _17109_ (.A(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__buf_4 _17110_ (.A(_03393_),
    .X(_03395_));
 sky130_fd_sc_hd__nor2_1 _17111_ (.A(_11210_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__a31o_1 _17112_ (.A1(_03236_),
    .A2(net2463),
    .A3(_03394_),
    .B1(_03396_),
    .X(_00104_));
 sky130_fd_sc_hd__nor2_1 _17113_ (.A(_03170_),
    .B(_03395_),
    .Y(_03397_));
 sky130_fd_sc_hd__a31o_1 _17114_ (.A1(_03236_),
    .A2(net753),
    .A3(_03394_),
    .B1(_03397_),
    .X(_00105_));
 sky130_fd_sc_hd__buf_4 _17115_ (.A(_08776_),
    .X(_03398_));
 sky130_fd_sc_hd__buf_4 _17116_ (.A(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__nor2_1 _17117_ (.A(_03219_),
    .B(_03395_),
    .Y(_03400_));
 sky130_fd_sc_hd__a31o_1 _17118_ (.A1(_03399_),
    .A2(net683),
    .A3(_03394_),
    .B1(_03400_),
    .X(_00106_));
 sky130_fd_sc_hd__and3_1 _17119_ (.A(_03392_),
    .B(_11040_),
    .C(_03296_),
    .X(_03401_));
 sky130_fd_sc_hd__a31o_1 _17120_ (.A1(_03399_),
    .A2(net1556),
    .A3(_03394_),
    .B1(_03401_),
    .X(_00107_));
 sky130_fd_sc_hd__buf_4 _17121_ (.A(_10930_),
    .X(_03402_));
 sky130_fd_sc_hd__nand2_1 _17122_ (.A(_03402_),
    .B(net4005),
    .Y(_03403_));
 sky130_fd_sc_hd__and2_1 _17123_ (.A(_03392_),
    .B(_08778_),
    .X(_03404_));
 sky130_fd_sc_hd__buf_4 _17124_ (.A(_03404_),
    .X(_03405_));
 sky130_fd_sc_hd__a22o_1 _17125_ (.A1(_03395_),
    .A2(_03403_),
    .B1(_03405_),
    .B2(_09201_),
    .X(_03406_));
 sky130_fd_sc_hd__inv_2 _17126_ (.A(_03406_),
    .Y(_00108_));
 sky130_fd_sc_hd__and3_1 _17127_ (.A(_03392_),
    .B(_11391_),
    .C(_03296_),
    .X(_03407_));
 sky130_fd_sc_hd__a31o_1 _17128_ (.A1(_03399_),
    .A2(net1165),
    .A3(_03394_),
    .B1(_03407_),
    .X(_00109_));
 sky130_fd_sc_hd__nor2_1 _17129_ (.A(_10872_),
    .B(_03395_),
    .Y(_03408_));
 sky130_fd_sc_hd__a31o_1 _17130_ (.A1(_03399_),
    .A2(net1363),
    .A3(_03394_),
    .B1(_03408_),
    .X(_00110_));
 sky130_fd_sc_hd__and3_1 _17131_ (.A(_03392_),
    .B(_10874_),
    .C(_03296_),
    .X(_03409_));
 sky130_fd_sc_hd__a31o_1 _17132_ (.A1(_03399_),
    .A2(net2229),
    .A3(_03394_),
    .B1(_03409_),
    .X(_00111_));
 sky130_fd_sc_hd__nor2_1 _17133_ (.A(_10760_),
    .B(_03395_),
    .Y(_03410_));
 sky130_fd_sc_hd__a31o_1 _17134_ (.A1(_03399_),
    .A2(net1828),
    .A3(_03394_),
    .B1(_03410_),
    .X(_00096_));
 sky130_fd_sc_hd__nand2_1 _17135_ (.A(_03402_),
    .B(net4066),
    .Y(_03411_));
 sky130_fd_sc_hd__a22o_1 _17136_ (.A1(_03395_),
    .A2(_03411_),
    .B1(_03405_),
    .B2(_10313_),
    .X(_03412_));
 sky130_fd_sc_hd__inv_2 _17137_ (.A(_03412_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_1 _17138_ (.A(_03402_),
    .B(net3951),
    .Y(_03413_));
 sky130_fd_sc_hd__a22o_1 _17139_ (.A1(_03395_),
    .A2(_03413_),
    .B1(_03405_),
    .B2(_10316_),
    .X(_03414_));
 sky130_fd_sc_hd__inv_2 _17140_ (.A(_03414_),
    .Y(_00098_));
 sky130_fd_sc_hd__nor2_1 _17141_ (.A(_02904_),
    .B(_03395_),
    .Y(_03415_));
 sky130_fd_sc_hd__a31o_1 _17142_ (.A1(_03399_),
    .A2(net1241),
    .A3(_03394_),
    .B1(_03415_),
    .X(_00099_));
 sky130_fd_sc_hd__nor2_1 _17143_ (.A(_03020_),
    .B(_03395_),
    .Y(_03416_));
 sky130_fd_sc_hd__a31o_1 _17144_ (.A1(_03399_),
    .A2(net1868),
    .A3(_03394_),
    .B1(_03416_),
    .X(_00100_));
 sky130_fd_sc_hd__nand2_1 _17145_ (.A(_03402_),
    .B(net4166),
    .Y(_03417_));
 sky130_fd_sc_hd__a22o_1 _17146_ (.A1(_03393_),
    .A2(_03417_),
    .B1(_03405_),
    .B2(_09338_),
    .X(_03418_));
 sky130_fd_sc_hd__inv_2 _17147_ (.A(_03418_),
    .Y(_00101_));
 sky130_fd_sc_hd__and3_1 _17148_ (.A(_03392_),
    .B(_11291_),
    .C(_03296_),
    .X(_03419_));
 sky130_fd_sc_hd__a31o_1 _17149_ (.A1(_03399_),
    .A2(net1669),
    .A3(_03394_),
    .B1(_03419_),
    .X(_00102_));
 sky130_fd_sc_hd__nor2_1 _17150_ (.A(_03026_),
    .B(_03395_),
    .Y(_03420_));
 sky130_fd_sc_hd__a31o_1 _17151_ (.A1(_03399_),
    .A2(net1315),
    .A3(_03394_),
    .B1(_03420_),
    .X(_00103_));
 sky130_fd_sc_hd__nand2_1 _17152_ (.A(_03402_),
    .B(net4001),
    .Y(_03421_));
 sky130_fd_sc_hd__a22o_1 _17153_ (.A1(_03393_),
    .A2(_03421_),
    .B1(_03405_),
    .B2(_09415_),
    .X(_03422_));
 sky130_fd_sc_hd__inv_2 _17154_ (.A(_03422_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_1 _17155_ (.A(_03402_),
    .B(net4044),
    .Y(_03423_));
 sky130_fd_sc_hd__a22o_1 _17156_ (.A1(_03393_),
    .A2(_03423_),
    .B1(_03405_),
    .B2(_09249_),
    .X(_03424_));
 sky130_fd_sc_hd__inv_2 _17157_ (.A(_03424_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _17158_ (.A(_03402_),
    .B(net4042),
    .Y(_03425_));
 sky130_fd_sc_hd__a22o_1 _17159_ (.A1(_03393_),
    .A2(_03425_),
    .B1(_03405_),
    .B2(_09348_),
    .X(_03426_));
 sky130_fd_sc_hd__inv_2 _17160_ (.A(_03426_),
    .Y(_00082_));
 sky130_fd_sc_hd__and3_1 _17161_ (.A(_03392_),
    .B(_03032_),
    .C(_03296_),
    .X(_03427_));
 sky130_fd_sc_hd__a31o_1 _17162_ (.A1(_03399_),
    .A2(net907),
    .A3(_03394_),
    .B1(_03427_),
    .X(_00083_));
 sky130_fd_sc_hd__nand2_1 _17163_ (.A(_03402_),
    .B(net3997),
    .Y(_03428_));
 sky130_fd_sc_hd__a22o_1 _17164_ (.A1(_03393_),
    .A2(_03428_),
    .B1(_03405_),
    .B2(_09354_),
    .X(_03429_));
 sky130_fd_sc_hd__inv_2 _17165_ (.A(_03429_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _17166_ (.A(_03402_),
    .B(net4207),
    .Y(_03430_));
 sky130_fd_sc_hd__a22o_1 _17167_ (.A1(_03393_),
    .A2(_03430_),
    .B1(_03405_),
    .B2(_10331_),
    .X(_03431_));
 sky130_fd_sc_hd__inv_2 _17168_ (.A(_03431_),
    .Y(_00085_));
 sky130_fd_sc_hd__and3_1 _17169_ (.A(_03392_),
    .B(_03087_),
    .C(_03296_),
    .X(_03432_));
 sky130_fd_sc_hd__a31o_1 _17170_ (.A1(_03399_),
    .A2(net1151),
    .A3(_03394_),
    .B1(_03432_),
    .X(_00086_));
 sky130_fd_sc_hd__nand2_1 _17171_ (.A(_03402_),
    .B(net4059),
    .Y(_03433_));
 sky130_fd_sc_hd__a22o_1 _17172_ (.A1(_03393_),
    .A2(_03433_),
    .B1(_03405_),
    .B2(_10335_),
    .X(_03434_));
 sky130_fd_sc_hd__inv_2 _17173_ (.A(_03434_),
    .Y(_00087_));
 sky130_fd_sc_hd__and3_1 _17174_ (.A(_03392_),
    .B(_03196_),
    .C(_03296_),
    .X(_03435_));
 sky130_fd_sc_hd__a31o_1 _17175_ (.A1(_03399_),
    .A2(net1247),
    .A3(_03394_),
    .B1(_03435_),
    .X(_00072_));
 sky130_fd_sc_hd__nor2_1 _17176_ (.A(_10681_),
    .B(_03395_),
    .Y(_03436_));
 sky130_fd_sc_hd__a31o_1 _17177_ (.A1(_03399_),
    .A2(net995),
    .A3(_03395_),
    .B1(_03436_),
    .X(_00073_));
 sky130_fd_sc_hd__nand2_1 _17178_ (.A(_03402_),
    .B(net4074),
    .Y(_03437_));
 sky130_fd_sc_hd__a22o_1 _17179_ (.A1(_03393_),
    .A2(_03437_),
    .B1(_03405_),
    .B2(_09280_),
    .X(_03438_));
 sky130_fd_sc_hd__inv_2 _17180_ (.A(_03438_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(_03402_),
    .B(net4184),
    .Y(_03439_));
 sky130_fd_sc_hd__a22o_1 _17182_ (.A1(_03393_),
    .A2(_03439_),
    .B1(_03405_),
    .B2(_10342_),
    .X(_03440_));
 sky130_fd_sc_hd__inv_2 _17183_ (.A(_03440_),
    .Y(_00075_));
 sky130_fd_sc_hd__nand2_1 _17184_ (.A(_03402_),
    .B(net4163),
    .Y(_03441_));
 sky130_fd_sc_hd__a22o_1 _17185_ (.A1(_03393_),
    .A2(_03441_),
    .B1(_03405_),
    .B2(_09288_),
    .X(_03442_));
 sky130_fd_sc_hd__inv_2 _17186_ (.A(_03442_),
    .Y(_00076_));
 sky130_fd_sc_hd__and3_1 _17187_ (.A(_03392_),
    .B(_11426_),
    .C(_03296_),
    .X(_03443_));
 sky130_fd_sc_hd__a31o_1 _17188_ (.A1(_03399_),
    .A2(net1689),
    .A3(_03395_),
    .B1(_03443_),
    .X(_00077_));
 sky130_fd_sc_hd__nand2_1 _17189_ (.A(_09196_),
    .B(net2683),
    .Y(_03444_));
 sky130_fd_sc_hd__a22oi_1 _17190_ (.A1(_03392_),
    .A2(_10348_),
    .B1(_03394_),
    .B2(_03444_),
    .Y(_00078_));
 sky130_fd_sc_hd__nor2_1 _17191_ (.A(_09299_),
    .B(_03395_),
    .Y(_03445_));
 sky130_fd_sc_hd__a31o_1 _17192_ (.A1(_03399_),
    .A2(net897),
    .A3(_03395_),
    .B1(_03445_),
    .X(_00079_));
 sky130_fd_sc_hd__buf_4 _17193_ (.A(_03398_),
    .X(_03446_));
 sky130_fd_sc_hd__nor2_4 _17194_ (.A(_03391_),
    .B(_10292_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_4 _17195_ (.A(_03447_),
    .B(_09226_),
    .Y(_03448_));
 sky130_fd_sc_hd__buf_4 _17196_ (.A(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__buf_4 _17197_ (.A(_03448_),
    .X(_03450_));
 sky130_fd_sc_hd__nor2_1 _17198_ (.A(_11210_),
    .B(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__a31o_1 _17199_ (.A1(_03446_),
    .A2(net2467),
    .A3(_03449_),
    .B1(_03451_),
    .X(_00064_));
 sky130_fd_sc_hd__nor2_1 _17200_ (.A(_03170_),
    .B(_03450_),
    .Y(_03452_));
 sky130_fd_sc_hd__a31o_1 _17201_ (.A1(_03446_),
    .A2(net1443),
    .A3(_03449_),
    .B1(_03452_),
    .X(_00065_));
 sky130_fd_sc_hd__nor2_1 _17202_ (.A(_03219_),
    .B(_03450_),
    .Y(_03453_));
 sky130_fd_sc_hd__a31o_1 _17203_ (.A1(_03446_),
    .A2(net1319),
    .A3(_03449_),
    .B1(_03453_),
    .X(_00066_));
 sky130_fd_sc_hd__nand2_1 _17204_ (.A(_03402_),
    .B(net4069),
    .Y(_03454_));
 sky130_fd_sc_hd__inv_2 _17205_ (.A(_03391_),
    .Y(_03455_));
 sky130_fd_sc_hd__and3_1 _17206_ (.A(_10291_),
    .B(_03455_),
    .C(_08778_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_4 _17207_ (.A(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__a22o_1 _17208_ (.A1(_03448_),
    .A2(_03454_),
    .B1(_03457_),
    .B2(_09195_),
    .X(_03458_));
 sky130_fd_sc_hd__inv_2 _17209_ (.A(_03458_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_1 _17210_ (.A(_03402_),
    .B(net4254),
    .Y(_03459_));
 sky130_fd_sc_hd__a22o_1 _17211_ (.A1(_03448_),
    .A2(_03459_),
    .B1(_03457_),
    .B2(_09201_),
    .X(_03460_));
 sky130_fd_sc_hd__inv_2 _17212_ (.A(_03460_),
    .Y(_00068_));
 sky130_fd_sc_hd__and3_1 _17213_ (.A(_03447_),
    .B(_11391_),
    .C(_03296_),
    .X(_03461_));
 sky130_fd_sc_hd__a31o_1 _17214_ (.A1(_03446_),
    .A2(net1341),
    .A3(_03449_),
    .B1(_03461_),
    .X(_00069_));
 sky130_fd_sc_hd__nand2_1 _17215_ (.A(_03402_),
    .B(net4178),
    .Y(_03462_));
 sky130_fd_sc_hd__a22o_1 _17216_ (.A1(_03448_),
    .A2(_03462_),
    .B1(_03457_),
    .B2(_09398_),
    .X(_03463_));
 sky130_fd_sc_hd__inv_2 _17217_ (.A(_03463_),
    .Y(_00070_));
 sky130_fd_sc_hd__buf_4 _17218_ (.A(_10930_),
    .X(_03464_));
 sky130_fd_sc_hd__nand2_1 _17219_ (.A(_03464_),
    .B(net4003),
    .Y(_03465_));
 sky130_fd_sc_hd__a22o_1 _17220_ (.A1(_03448_),
    .A2(_03465_),
    .B1(_03457_),
    .B2(_09212_),
    .X(_03466_));
 sky130_fd_sc_hd__inv_2 _17221_ (.A(_03466_),
    .Y(_00071_));
 sky130_fd_sc_hd__buf_12 _17222_ (.A(_09215_),
    .X(_03467_));
 sky130_fd_sc_hd__nor2_1 _17223_ (.A(_03467_),
    .B(_03450_),
    .Y(_03468_));
 sky130_fd_sc_hd__a31o_1 _17224_ (.A1(_03446_),
    .A2(net507),
    .A3(_03449_),
    .B1(_03468_),
    .X(_00056_));
 sky130_fd_sc_hd__nand2_1 _17225_ (.A(_03464_),
    .B(net3949),
    .Y(_03469_));
 sky130_fd_sc_hd__a22o_1 _17226_ (.A1(_03448_),
    .A2(_03469_),
    .B1(_03457_),
    .B2(_10313_),
    .X(_03470_));
 sky130_fd_sc_hd__inv_2 _17227_ (.A(_03470_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand2_1 _17228_ (.A(_03464_),
    .B(net4006),
    .Y(_03471_));
 sky130_fd_sc_hd__a22o_1 _17229_ (.A1(_03448_),
    .A2(_03471_),
    .B1(_03457_),
    .B2(_10316_),
    .X(_03472_));
 sky130_fd_sc_hd__inv_2 _17230_ (.A(_03472_),
    .Y(_00058_));
 sky130_fd_sc_hd__nor2_1 _17231_ (.A(_02904_),
    .B(_03450_),
    .Y(_03473_));
 sky130_fd_sc_hd__a31o_1 _17232_ (.A1(_03446_),
    .A2(net1610),
    .A3(_03449_),
    .B1(_03473_),
    .X(_00059_));
 sky130_fd_sc_hd__nor2_1 _17233_ (.A(_03020_),
    .B(_03450_),
    .Y(_03474_));
 sky130_fd_sc_hd__a31o_1 _17234_ (.A1(_03446_),
    .A2(net743),
    .A3(_03449_),
    .B1(_03474_),
    .X(_00060_));
 sky130_fd_sc_hd__nor2_1 _17235_ (.A(_02845_),
    .B(_03450_),
    .Y(_03475_));
 sky130_fd_sc_hd__a31o_1 _17236_ (.A1(_03446_),
    .A2(net1229),
    .A3(_03449_),
    .B1(_03475_),
    .X(_00061_));
 sky130_fd_sc_hd__and3_1 _17237_ (.A(_03447_),
    .B(_11291_),
    .C(_03296_),
    .X(_03476_));
 sky130_fd_sc_hd__a31o_1 _17238_ (.A1(_03446_),
    .A2(net1135),
    .A3(_03449_),
    .B1(_03476_),
    .X(_00062_));
 sky130_fd_sc_hd__nand2_1 _17239_ (.A(_03464_),
    .B(net4053),
    .Y(_03477_));
 sky130_fd_sc_hd__a22o_1 _17240_ (.A1(_03448_),
    .A2(_03477_),
    .B1(_03457_),
    .B2(_09768_),
    .X(_03478_));
 sky130_fd_sc_hd__inv_2 _17241_ (.A(_03478_),
    .Y(_00063_));
 sky130_fd_sc_hd__nor2_1 _17242_ (.A(_03294_),
    .B(_03450_),
    .Y(_03479_));
 sky130_fd_sc_hd__a31o_1 _17243_ (.A1(_03446_),
    .A2(net625),
    .A3(_03449_),
    .B1(_03479_),
    .X(_00048_));
 sky130_fd_sc_hd__clkbuf_4 _17244_ (.A(_11219_),
    .X(_03480_));
 sky130_fd_sc_hd__and3_1 _17245_ (.A(_03447_),
    .B(_03029_),
    .C(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__a31o_1 _17246_ (.A1(_03446_),
    .A2(net2437),
    .A3(_03449_),
    .B1(_03481_),
    .X(_00049_));
 sky130_fd_sc_hd__buf_12 _17247_ (.A(_09252_),
    .X(_03482_));
 sky130_fd_sc_hd__nor2_1 _17248_ (.A(_03482_),
    .B(_03450_),
    .Y(_03483_));
 sky130_fd_sc_hd__a31o_1 _17249_ (.A1(_03446_),
    .A2(net2233),
    .A3(_03449_),
    .B1(_03483_),
    .X(_00050_));
 sky130_fd_sc_hd__nand2_1 _17250_ (.A(_03464_),
    .B(net4014),
    .Y(_03484_));
 sky130_fd_sc_hd__a22o_1 _17251_ (.A1(_03448_),
    .A2(_03484_),
    .B1(_03457_),
    .B2(_09256_),
    .X(_03485_));
 sky130_fd_sc_hd__inv_2 _17252_ (.A(_03485_),
    .Y(_00051_));
 sky130_fd_sc_hd__nor2_1 _17253_ (.A(_11010_),
    .B(_03450_),
    .Y(_03486_));
 sky130_fd_sc_hd__a31o_1 _17254_ (.A1(_03446_),
    .A2(net1277),
    .A3(_03449_),
    .B1(_03486_),
    .X(_00052_));
 sky130_fd_sc_hd__nand2_1 _17255_ (.A(_03464_),
    .B(net4204),
    .Y(_03487_));
 sky130_fd_sc_hd__a22o_1 _17256_ (.A1(_03448_),
    .A2(_03487_),
    .B1(_03457_),
    .B2(_10331_),
    .X(_03488_));
 sky130_fd_sc_hd__inv_2 _17257_ (.A(_03488_),
    .Y(_00053_));
 sky130_fd_sc_hd__and3_1 _17258_ (.A(_03447_),
    .B(_03087_),
    .C(_03480_),
    .X(_03489_));
 sky130_fd_sc_hd__a31o_1 _17259_ (.A1(_03446_),
    .A2(net2099),
    .A3(_03449_),
    .B1(_03489_),
    .X(_00054_));
 sky130_fd_sc_hd__nand2_1 _17260_ (.A(_03464_),
    .B(net3972),
    .Y(_03490_));
 sky130_fd_sc_hd__a22o_1 _17261_ (.A1(_03448_),
    .A2(_03490_),
    .B1(_03457_),
    .B2(_10335_),
    .X(_03491_));
 sky130_fd_sc_hd__inv_2 _17262_ (.A(_03491_),
    .Y(_00055_));
 sky130_fd_sc_hd__and3_1 _17263_ (.A(_03447_),
    .B(_03196_),
    .C(_03480_),
    .X(_03492_));
 sky130_fd_sc_hd__a31o_1 _17264_ (.A1(_03446_),
    .A2(net1857),
    .A3(_03449_),
    .B1(_03492_),
    .X(_00040_));
 sky130_fd_sc_hd__nor2_1 _17265_ (.A(_10681_),
    .B(_03450_),
    .Y(_03493_));
 sky130_fd_sc_hd__a31o_1 _17266_ (.A1(_03446_),
    .A2(net941),
    .A3(_03449_),
    .B1(_03493_),
    .X(_00041_));
 sky130_fd_sc_hd__nand2_1 _17267_ (.A(_03464_),
    .B(net3962),
    .Y(_03494_));
 sky130_fd_sc_hd__a22o_1 _17268_ (.A1(_03448_),
    .A2(_03494_),
    .B1(_03457_),
    .B2(_09280_),
    .X(_03495_));
 sky130_fd_sc_hd__inv_2 _17269_ (.A(_03495_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand2_1 _17270_ (.A(_03464_),
    .B(net3974),
    .Y(_03496_));
 sky130_fd_sc_hd__a22o_1 _17271_ (.A1(_03448_),
    .A2(_03496_),
    .B1(_03457_),
    .B2(_10342_),
    .X(_03497_));
 sky130_fd_sc_hd__inv_2 _17272_ (.A(_03497_),
    .Y(_00043_));
 sky130_fd_sc_hd__buf_4 _17273_ (.A(_03398_),
    .X(_03498_));
 sky130_fd_sc_hd__and3_1 _17274_ (.A(_03447_),
    .B(_10848_),
    .C(_03480_),
    .X(_03499_));
 sky130_fd_sc_hd__a31o_1 _17275_ (.A1(_03498_),
    .A2(net539),
    .A3(_03450_),
    .B1(_03499_),
    .X(_00044_));
 sky130_fd_sc_hd__and3_1 _17276_ (.A(_03447_),
    .B(_11426_),
    .C(_03480_),
    .X(_03500_));
 sky130_fd_sc_hd__a31o_1 _17277_ (.A1(_03498_),
    .A2(net1167),
    .A3(_03450_),
    .B1(_03500_),
    .X(_00045_));
 sky130_fd_sc_hd__nand2_1 _17278_ (.A(_03368_),
    .B(net3305),
    .Y(_03501_));
 sky130_fd_sc_hd__a22o_1 _17279_ (.A1(_09296_),
    .A2(_03447_),
    .B1(_03450_),
    .B2(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__inv_2 _17280_ (.A(net3306),
    .Y(_00046_));
 sky130_fd_sc_hd__nor2_1 _17281_ (.A(_09299_),
    .B(_03450_),
    .Y(_03503_));
 sky130_fd_sc_hd__a31o_1 _17282_ (.A1(_03498_),
    .A2(net1601),
    .A3(_03450_),
    .B1(_03503_),
    .X(_00047_));
 sky130_fd_sc_hd__nor2_4 _17283_ (.A(_03391_),
    .B(_10356_),
    .Y(_03504_));
 sky130_fd_sc_hd__nand2_4 _17284_ (.A(_03504_),
    .B(_09226_),
    .Y(_03505_));
 sky130_fd_sc_hd__buf_4 _17285_ (.A(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__buf_4 _17286_ (.A(_03505_),
    .X(_03507_));
 sky130_fd_sc_hd__nor2_1 _17287_ (.A(_11210_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__a31o_1 _17288_ (.A1(_03498_),
    .A2(net1902),
    .A3(_03506_),
    .B1(_03508_),
    .X(_00032_));
 sky130_fd_sc_hd__nor2_1 _17289_ (.A(_03170_),
    .B(_03507_),
    .Y(_03509_));
 sky130_fd_sc_hd__a31o_1 _17290_ (.A1(_03498_),
    .A2(net1159),
    .A3(_03506_),
    .B1(_03509_),
    .X(_00033_));
 sky130_fd_sc_hd__nor2_1 _17291_ (.A(_03219_),
    .B(_03507_),
    .Y(_03510_));
 sky130_fd_sc_hd__a31o_1 _17292_ (.A1(_03498_),
    .A2(net2379),
    .A3(_03506_),
    .B1(_03510_),
    .X(_00034_));
 sky130_fd_sc_hd__and3_1 _17293_ (.A(_03504_),
    .B(_11040_),
    .C(_03480_),
    .X(_03511_));
 sky130_fd_sc_hd__a31o_1 _17294_ (.A1(_03498_),
    .A2(net701),
    .A3(_03506_),
    .B1(_03511_),
    .X(_00035_));
 sky130_fd_sc_hd__and3_1 _17295_ (.A(_03504_),
    .B(_10586_),
    .C(_03480_),
    .X(_03512_));
 sky130_fd_sc_hd__a31o_1 _17296_ (.A1(_03498_),
    .A2(net763),
    .A3(_03506_),
    .B1(_03512_),
    .X(_00036_));
 sky130_fd_sc_hd__nand2_1 _17297_ (.A(_03464_),
    .B(net3947),
    .Y(_03513_));
 sky130_fd_sc_hd__and3_1 _17298_ (.A(_10355_),
    .B(_03455_),
    .C(_08778_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_4 _17299_ (.A(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__a22o_1 _17300_ (.A1(_03505_),
    .A2(_03513_),
    .B1(_03515_),
    .B2(_09205_),
    .X(_03516_));
 sky130_fd_sc_hd__inv_2 _17301_ (.A(_03516_),
    .Y(_00037_));
 sky130_fd_sc_hd__nor2_1 _17302_ (.A(_10872_),
    .B(_03507_),
    .Y(_03517_));
 sky130_fd_sc_hd__a31o_1 _17303_ (.A1(_03498_),
    .A2(net1543),
    .A3(_03506_),
    .B1(_03517_),
    .X(_00038_));
 sky130_fd_sc_hd__and3_1 _17304_ (.A(_03504_),
    .B(_10874_),
    .C(_03480_),
    .X(_03518_));
 sky130_fd_sc_hd__a31o_1 _17305_ (.A1(_03498_),
    .A2(net1757),
    .A3(_03506_),
    .B1(_03518_),
    .X(_00039_));
 sky130_fd_sc_hd__nor2_1 _17306_ (.A(_03467_),
    .B(_03507_),
    .Y(_03519_));
 sky130_fd_sc_hd__a31o_1 _17307_ (.A1(_03498_),
    .A2(net2328),
    .A3(_03506_),
    .B1(_03519_),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_1 _17308_ (.A(_03464_),
    .B(net3868),
    .Y(_03520_));
 sky130_fd_sc_hd__a22o_1 _17309_ (.A1(_03505_),
    .A2(_03520_),
    .B1(_03515_),
    .B2(_10313_),
    .X(_03521_));
 sky130_fd_sc_hd__inv_2 _17310_ (.A(_03521_),
    .Y(_00025_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(_03464_),
    .B(net4235),
    .Y(_03522_));
 sky130_fd_sc_hd__a22o_1 _17312_ (.A1(_03505_),
    .A2(_03522_),
    .B1(_03515_),
    .B2(_10316_),
    .X(_03523_));
 sky130_fd_sc_hd__inv_2 _17313_ (.A(_03523_),
    .Y(_00026_));
 sky130_fd_sc_hd__nor2_1 _17314_ (.A(_02904_),
    .B(_03507_),
    .Y(_03524_));
 sky130_fd_sc_hd__a31o_1 _17315_ (.A1(_03498_),
    .A2(net1570),
    .A3(_03506_),
    .B1(_03524_),
    .X(_00027_));
 sky130_fd_sc_hd__nor2_1 _17316_ (.A(_03020_),
    .B(_03507_),
    .Y(_03525_));
 sky130_fd_sc_hd__a31o_1 _17317_ (.A1(_03498_),
    .A2(net923),
    .A3(_03506_),
    .B1(_03525_),
    .X(_00028_));
 sky130_fd_sc_hd__nand2_1 _17318_ (.A(_03464_),
    .B(net3927),
    .Y(_03526_));
 sky130_fd_sc_hd__a22o_1 _17319_ (.A1(_03505_),
    .A2(_03526_),
    .B1(_03515_),
    .B2(_09338_),
    .X(_03527_));
 sky130_fd_sc_hd__inv_2 _17320_ (.A(_03527_),
    .Y(_00029_));
 sky130_fd_sc_hd__and3_1 _17321_ (.A(_03504_),
    .B(_11291_),
    .C(_03480_),
    .X(_03528_));
 sky130_fd_sc_hd__a31o_1 _17322_ (.A1(_03498_),
    .A2(net937),
    .A3(_03506_),
    .B1(_03528_),
    .X(_00030_));
 sky130_fd_sc_hd__nor2_1 _17323_ (.A(_03026_),
    .B(_03507_),
    .Y(_03529_));
 sky130_fd_sc_hd__a31o_1 _17324_ (.A1(_03498_),
    .A2(net867),
    .A3(_03506_),
    .B1(_03529_),
    .X(_00031_));
 sky130_fd_sc_hd__nor2_1 _17325_ (.A(_03294_),
    .B(_03507_),
    .Y(_03530_));
 sky130_fd_sc_hd__a31o_1 _17326_ (.A1(_03498_),
    .A2(net2422),
    .A3(_03506_),
    .B1(_03530_),
    .X(_00016_));
 sky130_fd_sc_hd__nand2_1 _17327_ (.A(_03464_),
    .B(net4140),
    .Y(_03531_));
 sky130_fd_sc_hd__a22o_1 _17328_ (.A1(_03505_),
    .A2(_03531_),
    .B1(_03515_),
    .B2(_09249_),
    .X(_03532_));
 sky130_fd_sc_hd__inv_2 _17329_ (.A(_03532_),
    .Y(_00017_));
 sky130_fd_sc_hd__buf_4 _17330_ (.A(_03398_),
    .X(_03533_));
 sky130_fd_sc_hd__nor2_1 _17331_ (.A(_03482_),
    .B(_03507_),
    .Y(_03534_));
 sky130_fd_sc_hd__a31o_1 _17332_ (.A1(_03533_),
    .A2(net2506),
    .A3(_03506_),
    .B1(_03534_),
    .X(_00018_));
 sky130_fd_sc_hd__and3_1 _17333_ (.A(_03504_),
    .B(_03032_),
    .C(_03480_),
    .X(_03535_));
 sky130_fd_sc_hd__a31o_1 _17334_ (.A1(_03533_),
    .A2(net769),
    .A3(_03506_),
    .B1(_03535_),
    .X(_00019_));
 sky130_fd_sc_hd__nand2_1 _17335_ (.A(_03464_),
    .B(net4282),
    .Y(_03536_));
 sky130_fd_sc_hd__a22o_1 _17336_ (.A1(_03505_),
    .A2(_03536_),
    .B1(_03515_),
    .B2(_09354_),
    .X(_03537_));
 sky130_fd_sc_hd__inv_2 _17337_ (.A(_03537_),
    .Y(_00020_));
 sky130_fd_sc_hd__nand2_1 _17338_ (.A(_03464_),
    .B(net3969),
    .Y(_03538_));
 sky130_fd_sc_hd__a22o_1 _17339_ (.A1(_03505_),
    .A2(_03538_),
    .B1(_03515_),
    .B2(_10331_),
    .X(_03539_));
 sky130_fd_sc_hd__inv_2 _17340_ (.A(_03539_),
    .Y(_00021_));
 sky130_fd_sc_hd__and3_1 _17341_ (.A(_03504_),
    .B(_03087_),
    .C(_03480_),
    .X(_03540_));
 sky130_fd_sc_hd__a31o_1 _17342_ (.A1(_03533_),
    .A2(net1303),
    .A3(_03506_),
    .B1(_03540_),
    .X(_00022_));
 sky130_fd_sc_hd__buf_4 _17343_ (.A(_08776_),
    .X(_03541_));
 sky130_fd_sc_hd__nand2_1 _17344_ (.A(_03541_),
    .B(net4088),
    .Y(_03542_));
 sky130_fd_sc_hd__a22o_1 _17345_ (.A1(_03505_),
    .A2(_03542_),
    .B1(_03515_),
    .B2(_10335_),
    .X(_03543_));
 sky130_fd_sc_hd__inv_2 _17346_ (.A(_03543_),
    .Y(_00023_));
 sky130_fd_sc_hd__and3_1 _17347_ (.A(_03504_),
    .B(_03196_),
    .C(_03480_),
    .X(_03544_));
 sky130_fd_sc_hd__a31o_1 _17348_ (.A1(_03533_),
    .A2(net723),
    .A3(_03507_),
    .B1(_03544_),
    .X(_00008_));
 sky130_fd_sc_hd__nor2_1 _17349_ (.A(_10681_),
    .B(_03507_),
    .Y(_03545_));
 sky130_fd_sc_hd__a31o_1 _17350_ (.A1(_03533_),
    .A2(net1928),
    .A3(_03507_),
    .B1(_03545_),
    .X(_00009_));
 sky130_fd_sc_hd__nand2_1 _17351_ (.A(_03541_),
    .B(net4250),
    .Y(_03546_));
 sky130_fd_sc_hd__a22o_1 _17352_ (.A1(_03505_),
    .A2(_03546_),
    .B1(_03515_),
    .B2(_09280_),
    .X(_03547_));
 sky130_fd_sc_hd__inv_2 _17353_ (.A(_03547_),
    .Y(_00010_));
 sky130_fd_sc_hd__nand2_1 _17354_ (.A(_03541_),
    .B(net4248),
    .Y(_03548_));
 sky130_fd_sc_hd__a22o_1 _17355_ (.A1(_03505_),
    .A2(_03548_),
    .B1(_03515_),
    .B2(_10342_),
    .X(_03549_));
 sky130_fd_sc_hd__inv_2 _17356_ (.A(_03549_),
    .Y(_00011_));
 sky130_fd_sc_hd__buf_8 _17357_ (.A(net77),
    .X(_03550_));
 sky130_fd_sc_hd__and3_1 _17358_ (.A(_03504_),
    .B(_03550_),
    .C(_03480_),
    .X(_03551_));
 sky130_fd_sc_hd__a31o_1 _17359_ (.A1(_03533_),
    .A2(net1583),
    .A3(_03507_),
    .B1(_03551_),
    .X(_00012_));
 sky130_fd_sc_hd__nand2_1 _17360_ (.A(_03541_),
    .B(net4073),
    .Y(_03552_));
 sky130_fd_sc_hd__a22o_1 _17361_ (.A1(_03505_),
    .A2(_03552_),
    .B1(_03515_),
    .B2(net136),
    .X(_03553_));
 sky130_fd_sc_hd__inv_2 _17362_ (.A(_03553_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_1 _17363_ (.A(_03368_),
    .B(net3621),
    .Y(_03554_));
 sky130_fd_sc_hd__a22o_1 _17364_ (.A1(_09296_),
    .A2(_03504_),
    .B1(_03507_),
    .B2(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__inv_2 _17365_ (.A(net3622),
    .Y(_00014_));
 sky130_fd_sc_hd__nand2_1 _17366_ (.A(_03368_),
    .B(net3398),
    .Y(_03556_));
 sky130_fd_sc_hd__a22o_1 _17367_ (.A1(_09440_),
    .A2(_03504_),
    .B1(_03507_),
    .B2(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__inv_2 _17368_ (.A(net3399),
    .Y(_00015_));
 sky130_fd_sc_hd__nor2_2 _17369_ (.A(_03391_),
    .B(_10411_),
    .Y(_03558_));
 sky130_fd_sc_hd__inv_2 _17370_ (.A(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__nor2_1 _17371_ (.A(_08728_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__inv_2 _17372_ (.A(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__buf_4 _17373_ (.A(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__buf_4 _17374_ (.A(_03561_),
    .X(_03563_));
 sky130_fd_sc_hd__nor2_1 _17375_ (.A(_11210_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__a31o_1 _17376_ (.A1(_03533_),
    .A2(net2249),
    .A3(_03562_),
    .B1(_03564_),
    .X(_02544_));
 sky130_fd_sc_hd__nor2_1 _17377_ (.A(_03170_),
    .B(_03563_),
    .Y(_03565_));
 sky130_fd_sc_hd__a31o_1 _17378_ (.A1(_03533_),
    .A2(net969),
    .A3(_03562_),
    .B1(_03565_),
    .X(_02545_));
 sky130_fd_sc_hd__nor2_1 _17379_ (.A(_03219_),
    .B(_03563_),
    .Y(_03566_));
 sky130_fd_sc_hd__a31o_1 _17380_ (.A1(_03533_),
    .A2(net1713),
    .A3(_03562_),
    .B1(_03566_),
    .X(_02546_));
 sky130_fd_sc_hd__and3_1 _17381_ (.A(_03558_),
    .B(_11040_),
    .C(_03480_),
    .X(_03567_));
 sky130_fd_sc_hd__a31o_1 _17382_ (.A1(_03562_),
    .A2(_03278_),
    .A3(net2399),
    .B1(_03567_),
    .X(_02547_));
 sky130_fd_sc_hd__and3_1 _17383_ (.A(_03558_),
    .B(_10586_),
    .C(_03480_),
    .X(_03568_));
 sky130_fd_sc_hd__a31o_1 _17384_ (.A1(_03562_),
    .A2(_03278_),
    .A3(net1081),
    .B1(_03568_),
    .X(_02548_));
 sky130_fd_sc_hd__and3_1 _17385_ (.A(_03558_),
    .B(_11391_),
    .C(_03480_),
    .X(_03569_));
 sky130_fd_sc_hd__a31o_1 _17386_ (.A1(_03562_),
    .A2(_03278_),
    .A3(net1900),
    .B1(_03569_),
    .X(_02549_));
 sky130_fd_sc_hd__nor2_8 _17387_ (.A(_08794_),
    .B(_03559_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand2_1 _17388_ (.A(_03368_),
    .B(net3327),
    .Y(_03571_));
 sky130_fd_sc_hd__a22o_1 _17389_ (.A1(_03570_),
    .A2(_11105_),
    .B1(_03563_),
    .B2(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__inv_2 _17390_ (.A(_03572_),
    .Y(_02550_));
 sky130_fd_sc_hd__nand2_1 _17391_ (.A(_03368_),
    .B(net3310),
    .Y(_03573_));
 sky130_fd_sc_hd__a22o_1 _17392_ (.A1(_03570_),
    .A2(_10591_),
    .B1(_03563_),
    .B2(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__inv_2 _17393_ (.A(_03574_),
    .Y(_02551_));
 sky130_fd_sc_hd__nand2_1 _17394_ (.A(_03368_),
    .B(net2790),
    .Y(_03575_));
 sky130_fd_sc_hd__a22o_1 _17395_ (.A1(_03570_),
    .A2(net135),
    .B1(_03563_),
    .B2(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__inv_2 _17396_ (.A(_03576_),
    .Y(_02536_));
 sky130_fd_sc_hd__buf_4 _17397_ (.A(_03271_),
    .X(_03577_));
 sky130_fd_sc_hd__nand2_1 _17398_ (.A(_03577_),
    .B(net3635),
    .Y(_03578_));
 sky130_fd_sc_hd__a22o_1 _17399_ (.A1(_03570_),
    .A2(_02899_),
    .B1(_03563_),
    .B2(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__inv_2 _17400_ (.A(_03579_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2_1 _17401_ (.A(_03577_),
    .B(net3241),
    .Y(_03580_));
 sky130_fd_sc_hd__a22o_1 _17402_ (.A1(_03570_),
    .A2(_02963_),
    .B1(_03563_),
    .B2(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__inv_2 _17403_ (.A(_03581_),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2_1 _17404_ (.A(_03577_),
    .B(net2981),
    .Y(_03582_));
 sky130_fd_sc_hd__a22o_1 _17405_ (.A1(_03570_),
    .A2(_09589_),
    .B1(_03563_),
    .B2(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__inv_2 _17406_ (.A(_03583_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor2_1 _17407_ (.A(_03020_),
    .B(_03563_),
    .Y(_03584_));
 sky130_fd_sc_hd__a31o_1 _17408_ (.A1(_03533_),
    .A2(net833),
    .A3(_03562_),
    .B1(_03584_),
    .X(_02540_));
 sky130_fd_sc_hd__nand2_1 _17409_ (.A(_03577_),
    .B(net3015),
    .Y(_03585_));
 sky130_fd_sc_hd__a22o_1 _17410_ (.A1(_03570_),
    .A2(_09338_),
    .B1(_03563_),
    .B2(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__inv_2 _17411_ (.A(_03586_),
    .Y(_02541_));
 sky130_fd_sc_hd__clkbuf_4 _17412_ (.A(_11219_),
    .X(_03587_));
 sky130_fd_sc_hd__and3_1 _17413_ (.A(_03558_),
    .B(_11291_),
    .C(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__a31o_1 _17414_ (.A1(_03562_),
    .A2(_03278_),
    .A3(net2208),
    .B1(_03588_),
    .X(_02542_));
 sky130_fd_sc_hd__nand2_1 _17415_ (.A(_03577_),
    .B(net2915),
    .Y(_03589_));
 sky130_fd_sc_hd__a22o_1 _17416_ (.A1(_03570_),
    .A2(_09768_),
    .B1(_03563_),
    .B2(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__inv_2 _17417_ (.A(_03590_),
    .Y(_02543_));
 sky130_fd_sc_hd__nor2_1 _17418_ (.A(_03294_),
    .B(_03563_),
    .Y(_03591_));
 sky130_fd_sc_hd__a31o_1 _17419_ (.A1(_03533_),
    .A2(net1639),
    .A3(_03562_),
    .B1(_03591_),
    .X(_02528_));
 sky130_fd_sc_hd__and3_1 _17420_ (.A(_03558_),
    .B(_03029_),
    .C(_03587_),
    .X(_03592_));
 sky130_fd_sc_hd__a31o_1 _17421_ (.A1(_03562_),
    .A2(_03278_),
    .A3(net2509),
    .B1(_03592_),
    .X(_02529_));
 sky130_fd_sc_hd__nor2_1 _17422_ (.A(_03482_),
    .B(_03563_),
    .Y(_03593_));
 sky130_fd_sc_hd__a31o_1 _17423_ (.A1(_03533_),
    .A2(net1079),
    .A3(_03562_),
    .B1(_03593_),
    .X(_02530_));
 sky130_fd_sc_hd__nand2_1 _17424_ (.A(_03577_),
    .B(net3712),
    .Y(_03594_));
 sky130_fd_sc_hd__a22o_1 _17425_ (.A1(_03570_),
    .A2(_09255_),
    .B1(_03561_),
    .B2(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__inv_2 _17426_ (.A(_03595_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_1 _17427_ (.A(_11010_),
    .B(_03563_),
    .Y(_03596_));
 sky130_fd_sc_hd__a31o_1 _17428_ (.A1(_03533_),
    .A2(net1291),
    .A3(_03562_),
    .B1(_03596_),
    .X(_02532_));
 sky130_fd_sc_hd__nand2_1 _17429_ (.A(_03577_),
    .B(net3409),
    .Y(_03597_));
 sky130_fd_sc_hd__a22o_1 _17430_ (.A1(_03570_),
    .A2(_02916_),
    .B1(_03561_),
    .B2(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__inv_2 _17431_ (.A(_03598_),
    .Y(_02533_));
 sky130_fd_sc_hd__nand2_1 _17432_ (.A(_03577_),
    .B(net2807),
    .Y(_03599_));
 sky130_fd_sc_hd__a22o_1 _17433_ (.A1(_03570_),
    .A2(_09425_),
    .B1(_03561_),
    .B2(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__inv_2 _17434_ (.A(_03600_),
    .Y(_02534_));
 sky130_fd_sc_hd__nand2_1 _17435_ (.A(_03577_),
    .B(net2843),
    .Y(_03601_));
 sky130_fd_sc_hd__a22o_1 _17436_ (.A1(_03570_),
    .A2(_02921_),
    .B1(_03561_),
    .B2(_03601_),
    .X(_03602_));
 sky130_fd_sc_hd__inv_2 _17437_ (.A(_03602_),
    .Y(_02535_));
 sky130_fd_sc_hd__nand2_1 _17438_ (.A(_03577_),
    .B(net3513),
    .Y(_03603_));
 sky130_fd_sc_hd__a22o_1 _17439_ (.A1(_03570_),
    .A2(net141),
    .B1(_03561_),
    .B2(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__inv_2 _17440_ (.A(_03604_),
    .Y(_02520_));
 sky130_fd_sc_hd__clkbuf_16 _17441_ (.A(_09276_),
    .X(_03605_));
 sky130_fd_sc_hd__nor2_1 _17442_ (.A(_03605_),
    .B(_03563_),
    .Y(_03606_));
 sky130_fd_sc_hd__a31o_1 _17443_ (.A1(_03533_),
    .A2(net1651),
    .A3(_03562_),
    .B1(_03606_),
    .X(_02521_));
 sky130_fd_sc_hd__and3_1 _17444_ (.A(_03558_),
    .B(_03199_),
    .C(_03587_),
    .X(_03607_));
 sky130_fd_sc_hd__a31o_1 _17445_ (.A1(_03562_),
    .A2(_03278_),
    .A3(net2630),
    .B1(_03607_),
    .X(_02522_));
 sky130_fd_sc_hd__nand2_1 _17446_ (.A(_03577_),
    .B(net3437),
    .Y(_03608_));
 sky130_fd_sc_hd__a22o_1 _17447_ (.A1(_03570_),
    .A2(_02928_),
    .B1(_03561_),
    .B2(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__inv_2 _17448_ (.A(_03609_),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _17449_ (.A(_03577_),
    .B(net3769),
    .Y(_03610_));
 sky130_fd_sc_hd__a22o_1 _17450_ (.A1(_03570_),
    .A2(net139),
    .B1(_03561_),
    .B2(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__inv_2 _17451_ (.A(_03611_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand2_1 _17452_ (.A(_03577_),
    .B(net3548),
    .Y(_03612_));
 sky130_fd_sc_hd__a22o_1 _17453_ (.A1(_03570_),
    .A2(net136),
    .B1(_03561_),
    .B2(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__inv_2 _17454_ (.A(_03613_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand2_1 _17455_ (.A(_03317_),
    .B(net3831),
    .Y(_03614_));
 sky130_fd_sc_hd__o2bb2a_1 _17456_ (.A1_N(_03614_),
    .A2_N(_03562_),
    .B1(_02992_),
    .B2(_03559_),
    .X(_02526_));
 sky130_fd_sc_hd__nand2_1 _17457_ (.A(_03317_),
    .B(net3902),
    .Y(_03615_));
 sky130_fd_sc_hd__o2bb2a_1 _17458_ (.A1_N(_03615_),
    .A2_N(_03562_),
    .B1(_11316_),
    .B2(_03559_),
    .X(_02527_));
 sky130_fd_sc_hd__nand2_8 _17459_ (.A(_09735_),
    .B(_03163_),
    .Y(_03616_));
 sky130_fd_sc_hd__nor2_4 _17460_ (.A(_10469_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__inv_2 _17461_ (.A(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__nor2_1 _17462_ (.A(_09304_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__inv_2 _17463_ (.A(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__buf_4 _17464_ (.A(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__buf_4 _17465_ (.A(_03620_),
    .X(_03622_));
 sky130_fd_sc_hd__nor2_1 _17466_ (.A(_11210_),
    .B(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__a31o_1 _17467_ (.A1(_03533_),
    .A2(net1767),
    .A3(_03621_),
    .B1(_03623_),
    .X(_02512_));
 sky130_fd_sc_hd__nor2_1 _17468_ (.A(_03170_),
    .B(_03622_),
    .Y(_03624_));
 sky130_fd_sc_hd__a31o_1 _17469_ (.A1(_03533_),
    .A2(net1686),
    .A3(_03621_),
    .B1(_03624_),
    .X(_02513_));
 sky130_fd_sc_hd__nor2_4 _17470_ (.A(_09190_),
    .B(_03618_),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_1 _17471_ (.A(_03577_),
    .B(net3264),
    .Y(_03626_));
 sky130_fd_sc_hd__a22o_1 _17472_ (.A1(_03625_),
    .A2(_09459_),
    .B1(_03622_),
    .B2(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__inv_2 _17473_ (.A(_03627_),
    .Y(_02514_));
 sky130_fd_sc_hd__and3_1 _17474_ (.A(_03617_),
    .B(_11040_),
    .C(_03587_),
    .X(_03628_));
 sky130_fd_sc_hd__a31o_1 _17475_ (.A1(_03621_),
    .A2(_03278_),
    .A3(net2443),
    .B1(_03628_),
    .X(_02515_));
 sky130_fd_sc_hd__buf_4 _17476_ (.A(_10645_),
    .X(_03629_));
 sky130_fd_sc_hd__and3_1 _17477_ (.A(_03617_),
    .B(_10586_),
    .C(_03587_),
    .X(_03630_));
 sky130_fd_sc_hd__a31o_1 _17478_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2236),
    .B1(_03630_),
    .X(_02516_));
 sky130_fd_sc_hd__and3_1 _17479_ (.A(_03617_),
    .B(_11391_),
    .C(_03587_),
    .X(_03631_));
 sky130_fd_sc_hd__a31o_1 _17480_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2425),
    .B1(_03631_),
    .X(_02517_));
 sky130_fd_sc_hd__buf_4 _17481_ (.A(_03398_),
    .X(_03632_));
 sky130_fd_sc_hd__nor2_1 _17482_ (.A(_09208_),
    .B(_03622_),
    .Y(_03633_));
 sky130_fd_sc_hd__a31o_1 _17483_ (.A1(_03632_),
    .A2(net2322),
    .A3(_03621_),
    .B1(_03633_),
    .X(_02518_));
 sky130_fd_sc_hd__and3_1 _17484_ (.A(_03617_),
    .B(_10874_),
    .C(_03587_),
    .X(_03634_));
 sky130_fd_sc_hd__a31o_1 _17485_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2485),
    .B1(_03634_),
    .X(_02519_));
 sky130_fd_sc_hd__nor2_1 _17486_ (.A(_03467_),
    .B(_03622_),
    .Y(_03635_));
 sky130_fd_sc_hd__a31o_1 _17487_ (.A1(_03632_),
    .A2(net1191),
    .A3(_03621_),
    .B1(_03635_),
    .X(_02504_));
 sky130_fd_sc_hd__nand2_1 _17488_ (.A(_03577_),
    .B(net3433),
    .Y(_03636_));
 sky130_fd_sc_hd__a22o_1 _17489_ (.A1(_03625_),
    .A2(_02899_),
    .B1(_03622_),
    .B2(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__inv_2 _17490_ (.A(_03637_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_1 _17491_ (.A(_03577_),
    .B(net3366),
    .Y(_03638_));
 sky130_fd_sc_hd__a22o_1 _17492_ (.A1(_03625_),
    .A2(_02963_),
    .B1(_03620_),
    .B2(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__inv_2 _17493_ (.A(_03639_),
    .Y(_02506_));
 sky130_fd_sc_hd__nor2_1 _17494_ (.A(_02904_),
    .B(_03622_),
    .Y(_03640_));
 sky130_fd_sc_hd__a31o_1 _17495_ (.A1(_03632_),
    .A2(net2021),
    .A3(_03622_),
    .B1(_03640_),
    .X(_02507_));
 sky130_fd_sc_hd__nor2_1 _17496_ (.A(_03020_),
    .B(_03622_),
    .Y(_03641_));
 sky130_fd_sc_hd__a31o_1 _17497_ (.A1(_03632_),
    .A2(net1616),
    .A3(_03622_),
    .B1(_03641_),
    .X(_02508_));
 sky130_fd_sc_hd__nor2_1 _17498_ (.A(_02845_),
    .B(_03622_),
    .Y(_03642_));
 sky130_fd_sc_hd__a31o_1 _17499_ (.A1(_03632_),
    .A2(net2228),
    .A3(_03622_),
    .B1(_03642_),
    .X(_02509_));
 sky130_fd_sc_hd__and3_1 _17500_ (.A(_03617_),
    .B(_11291_),
    .C(_03587_),
    .X(_03643_));
 sky130_fd_sc_hd__a31o_1 _17501_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net1749),
    .B1(_03643_),
    .X(_02510_));
 sky130_fd_sc_hd__clkbuf_8 _17502_ (.A(_03271_),
    .X(_03644_));
 sky130_fd_sc_hd__nand2_1 _17503_ (.A(_03644_),
    .B(net3244),
    .Y(_03645_));
 sky130_fd_sc_hd__a22o_1 _17504_ (.A1(_03625_),
    .A2(_09767_),
    .B1(_03620_),
    .B2(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__inv_2 _17505_ (.A(_03646_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2_1 _17506_ (.A(_03644_),
    .B(net3833),
    .Y(_03647_));
 sky130_fd_sc_hd__a22o_1 _17507_ (.A1(_03625_),
    .A2(net138),
    .B1(_03620_),
    .B2(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__inv_2 _17508_ (.A(_03648_),
    .Y(_02496_));
 sky130_fd_sc_hd__and3_1 _17509_ (.A(_03617_),
    .B(_03029_),
    .C(_03587_),
    .X(_03649_));
 sky130_fd_sc_hd__a31o_1 _17510_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2429),
    .B1(_03649_),
    .X(_02497_));
 sky130_fd_sc_hd__nor2_1 _17511_ (.A(_03482_),
    .B(_03622_),
    .Y(_03650_));
 sky130_fd_sc_hd__a31o_1 _17512_ (.A1(_03632_),
    .A2(net1936),
    .A3(_03622_),
    .B1(_03650_),
    .X(_02498_));
 sky130_fd_sc_hd__and3_1 _17513_ (.A(_03617_),
    .B(_03032_),
    .C(_03587_),
    .X(_03651_));
 sky130_fd_sc_hd__a31o_1 _17514_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2077),
    .B1(_03651_),
    .X(_02499_));
 sky130_fd_sc_hd__nand2_1 _17515_ (.A(_03644_),
    .B(net3040),
    .Y(_03652_));
 sky130_fd_sc_hd__a22o_1 _17516_ (.A1(_03625_),
    .A2(_11136_),
    .B1(_03620_),
    .B2(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__inv_2 _17517_ (.A(_03653_),
    .Y(_02500_));
 sky130_fd_sc_hd__nand2_1 _17518_ (.A(_03644_),
    .B(net3781),
    .Y(_03654_));
 sky130_fd_sc_hd__a22o_1 _17519_ (.A1(_03625_),
    .A2(_02916_),
    .B1(_03620_),
    .B2(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__inv_2 _17520_ (.A(_03655_),
    .Y(_02501_));
 sky130_fd_sc_hd__nand2_1 _17521_ (.A(_03644_),
    .B(net2852),
    .Y(_03656_));
 sky130_fd_sc_hd__a22o_1 _17522_ (.A1(_03625_),
    .A2(_09424_),
    .B1(_03620_),
    .B2(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__inv_2 _17523_ (.A(_03657_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(_03644_),
    .B(net2846),
    .Y(_03658_));
 sky130_fd_sc_hd__a22o_1 _17525_ (.A1(_03625_),
    .A2(_02921_),
    .B1(_03620_),
    .B2(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__inv_2 _17526_ (.A(_03659_),
    .Y(_02503_));
 sky130_fd_sc_hd__and3_1 _17527_ (.A(_03617_),
    .B(_03196_),
    .C(_03587_),
    .X(_03660_));
 sky130_fd_sc_hd__a31o_1 _17528_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2264),
    .B1(_03660_),
    .X(_02488_));
 sky130_fd_sc_hd__nor2_1 _17529_ (.A(_03605_),
    .B(_03622_),
    .Y(_03661_));
 sky130_fd_sc_hd__a31o_1 _17530_ (.A1(_03632_),
    .A2(net1999),
    .A3(_03622_),
    .B1(_03661_),
    .X(_02489_));
 sky130_fd_sc_hd__and3_1 _17531_ (.A(_03617_),
    .B(_03199_),
    .C(_03587_),
    .X(_03662_));
 sky130_fd_sc_hd__a31o_1 _17532_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2369),
    .B1(_03662_),
    .X(_02490_));
 sky130_fd_sc_hd__nand2_1 _17533_ (.A(_03644_),
    .B(net3849),
    .Y(_03663_));
 sky130_fd_sc_hd__a22o_1 _17534_ (.A1(_03625_),
    .A2(_02928_),
    .B1(_03620_),
    .B2(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__inv_2 _17535_ (.A(_03664_),
    .Y(_02491_));
 sky130_fd_sc_hd__and3_1 _17536_ (.A(_03617_),
    .B(_03550_),
    .C(_03587_),
    .X(_03665_));
 sky130_fd_sc_hd__a31o_1 _17537_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net1782),
    .B1(_03665_),
    .X(_02492_));
 sky130_fd_sc_hd__and3_1 _17538_ (.A(_03617_),
    .B(_11426_),
    .C(_03587_),
    .X(_03666_));
 sky130_fd_sc_hd__a31o_1 _17539_ (.A1(_03621_),
    .A2(_03629_),
    .A3(net2527),
    .B1(_03666_),
    .X(_02493_));
 sky130_fd_sc_hd__nand2_1 _17540_ (.A(_03317_),
    .B(net3628),
    .Y(_03667_));
 sky130_fd_sc_hd__o2bb2a_1 _17541_ (.A1_N(_03667_),
    .A2_N(_03621_),
    .B1(_02992_),
    .B2(_03618_),
    .X(_02494_));
 sky130_fd_sc_hd__nand2_1 _17542_ (.A(_08777_),
    .B(net2752),
    .Y(_03668_));
 sky130_fd_sc_hd__a32o_1 _17543_ (.A1(_03625_),
    .A2(_08791_),
    .A3(_09299_),
    .B1(_03620_),
    .B2(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__inv_2 _17544_ (.A(net2753),
    .Y(_02495_));
 sky130_fd_sc_hd__nor2_4 _17545_ (.A(_03616_),
    .B(_10292_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_4 _17546_ (.A(_03670_),
    .B(_10413_),
    .Y(_03671_));
 sky130_fd_sc_hd__buf_4 _17547_ (.A(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__buf_4 _17548_ (.A(_03671_),
    .X(_03673_));
 sky130_fd_sc_hd__nor2_1 _17549_ (.A(_11210_),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__a31o_1 _17550_ (.A1(_03632_),
    .A2(net2034),
    .A3(_03672_),
    .B1(_03674_),
    .X(_02480_));
 sky130_fd_sc_hd__nor2_1 _17551_ (.A(_03170_),
    .B(_03673_),
    .Y(_03675_));
 sky130_fd_sc_hd__a31o_1 _17552_ (.A1(_03632_),
    .A2(net979),
    .A3(_03672_),
    .B1(_03675_),
    .X(_02481_));
 sky130_fd_sc_hd__nand2_1 _17553_ (.A(_03541_),
    .B(net4019),
    .Y(_03676_));
 sky130_fd_sc_hd__inv_2 _17554_ (.A(_03616_),
    .Y(_03677_));
 sky130_fd_sc_hd__and3_1 _17555_ (.A(_10291_),
    .B(_03677_),
    .C(_08778_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_4 _17556_ (.A(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__a22o_1 _17557_ (.A1(_03673_),
    .A2(_03676_),
    .B1(_03679_),
    .B2(_09460_),
    .X(_03680_));
 sky130_fd_sc_hd__inv_2 _17558_ (.A(_03680_),
    .Y(_02482_));
 sky130_fd_sc_hd__and3_1 _17559_ (.A(_03670_),
    .B(net69),
    .C(_03587_),
    .X(_03681_));
 sky130_fd_sc_hd__a31o_1 _17560_ (.A1(_03632_),
    .A2(net1043),
    .A3(_03672_),
    .B1(_03681_),
    .X(_02483_));
 sky130_fd_sc_hd__nand2_1 _17561_ (.A(_03541_),
    .B(net4176),
    .Y(_03682_));
 sky130_fd_sc_hd__a22o_1 _17562_ (.A1(_03671_),
    .A2(_03682_),
    .B1(_03679_),
    .B2(_09201_),
    .X(_03683_));
 sky130_fd_sc_hd__inv_2 _17563_ (.A(_03683_),
    .Y(_02484_));
 sky130_fd_sc_hd__and3_1 _17564_ (.A(_03670_),
    .B(_11391_),
    .C(_03587_),
    .X(_03684_));
 sky130_fd_sc_hd__a31o_1 _17565_ (.A1(_03632_),
    .A2(net1327),
    .A3(_03672_),
    .B1(_03684_),
    .X(_02485_));
 sky130_fd_sc_hd__nor2_1 _17566_ (.A(_09208_),
    .B(_03673_),
    .Y(_03685_));
 sky130_fd_sc_hd__a31o_1 _17567_ (.A1(_03632_),
    .A2(net1251),
    .A3(_03672_),
    .B1(_03685_),
    .X(_02486_));
 sky130_fd_sc_hd__nand2_1 _17568_ (.A(_03541_),
    .B(net4164),
    .Y(_03686_));
 sky130_fd_sc_hd__a22o_1 _17569_ (.A1(_03671_),
    .A2(_03686_),
    .B1(_03679_),
    .B2(_09212_),
    .X(_03687_));
 sky130_fd_sc_hd__inv_2 _17570_ (.A(_03687_),
    .Y(_02487_));
 sky130_fd_sc_hd__nor2_1 _17571_ (.A(_03467_),
    .B(_03673_),
    .Y(_03688_));
 sky130_fd_sc_hd__a31o_1 _17572_ (.A1(_03632_),
    .A2(net2633),
    .A3(_03672_),
    .B1(_03688_),
    .X(_02472_));
 sky130_fd_sc_hd__nand2_1 _17573_ (.A(_03541_),
    .B(net4177),
    .Y(_03689_));
 sky130_fd_sc_hd__a22o_1 _17574_ (.A1(_03671_),
    .A2(_03689_),
    .B1(_03679_),
    .B2(_10313_),
    .X(_03690_));
 sky130_fd_sc_hd__inv_2 _17575_ (.A(_03690_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand2_1 _17576_ (.A(_03541_),
    .B(net4107),
    .Y(_03691_));
 sky130_fd_sc_hd__a22o_1 _17577_ (.A1(_03671_),
    .A2(_03691_),
    .B1(_03679_),
    .B2(_10316_),
    .X(_03692_));
 sky130_fd_sc_hd__inv_2 _17578_ (.A(_03692_),
    .Y(_02474_));
 sky130_fd_sc_hd__nor2_1 _17579_ (.A(_02904_),
    .B(_03673_),
    .Y(_03693_));
 sky130_fd_sc_hd__a31o_1 _17580_ (.A1(_03632_),
    .A2(net2417),
    .A3(_03672_),
    .B1(_03693_),
    .X(_02475_));
 sky130_fd_sc_hd__nor2_1 _17581_ (.A(_03020_),
    .B(_03673_),
    .Y(_03694_));
 sky130_fd_sc_hd__a31o_1 _17582_ (.A1(_03632_),
    .A2(net1077),
    .A3(_03672_),
    .B1(_03694_),
    .X(_02476_));
 sky130_fd_sc_hd__nor2_1 _17583_ (.A(_02845_),
    .B(_03673_),
    .Y(_03695_));
 sky130_fd_sc_hd__a31o_1 _17584_ (.A1(_03632_),
    .A2(net2180),
    .A3(_03672_),
    .B1(_03695_),
    .X(_02477_));
 sky130_fd_sc_hd__buf_4 _17585_ (.A(_03398_),
    .X(_03696_));
 sky130_fd_sc_hd__buf_4 _17586_ (.A(_11219_),
    .X(_03697_));
 sky130_fd_sc_hd__and3_1 _17587_ (.A(_03670_),
    .B(_11291_),
    .C(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__a31o_1 _17588_ (.A1(_03696_),
    .A2(net1193),
    .A3(_03672_),
    .B1(_03698_),
    .X(_02478_));
 sky130_fd_sc_hd__nor2_1 _17589_ (.A(_03026_),
    .B(_03673_),
    .Y(_03699_));
 sky130_fd_sc_hd__a31o_1 _17590_ (.A1(_03696_),
    .A2(net2319),
    .A3(_03672_),
    .B1(_03699_),
    .X(_02479_));
 sky130_fd_sc_hd__nand2_1 _17591_ (.A(_03541_),
    .B(net4269),
    .Y(_03700_));
 sky130_fd_sc_hd__a22o_1 _17592_ (.A1(_03671_),
    .A2(_03700_),
    .B1(_03679_),
    .B2(_09415_),
    .X(_03701_));
 sky130_fd_sc_hd__inv_2 _17593_ (.A(_03701_),
    .Y(_02456_));
 sky130_fd_sc_hd__and3_1 _17594_ (.A(_03670_),
    .B(_03029_),
    .C(_03697_),
    .X(_03702_));
 sky130_fd_sc_hd__a31o_1 _17595_ (.A1(_03696_),
    .A2(net2068),
    .A3(_03672_),
    .B1(_03702_),
    .X(_02457_));
 sky130_fd_sc_hd__nand2_1 _17596_ (.A(_03541_),
    .B(net4155),
    .Y(_03703_));
 sky130_fd_sc_hd__a22o_1 _17597_ (.A1(_03671_),
    .A2(_03703_),
    .B1(_03679_),
    .B2(_09348_),
    .X(_03704_));
 sky130_fd_sc_hd__inv_2 _17598_ (.A(_03704_),
    .Y(_02458_));
 sky130_fd_sc_hd__and3_1 _17599_ (.A(_03670_),
    .B(_03032_),
    .C(_03697_),
    .X(_03705_));
 sky130_fd_sc_hd__a31o_1 _17600_ (.A1(_03696_),
    .A2(net597),
    .A3(_03672_),
    .B1(_03705_),
    .X(_02459_));
 sky130_fd_sc_hd__nor2_1 _17601_ (.A(_09259_),
    .B(_03673_),
    .Y(_03706_));
 sky130_fd_sc_hd__a31o_1 _17602_ (.A1(_03696_),
    .A2(net1924),
    .A3(_03672_),
    .B1(_03706_),
    .X(_02460_));
 sky130_fd_sc_hd__nand2_1 _17603_ (.A(_03541_),
    .B(net4031),
    .Y(_03707_));
 sky130_fd_sc_hd__a22o_1 _17604_ (.A1(_03671_),
    .A2(_03707_),
    .B1(_03679_),
    .B2(_10331_),
    .X(_03708_));
 sky130_fd_sc_hd__inv_2 _17605_ (.A(_03708_),
    .Y(_02461_));
 sky130_fd_sc_hd__and3_1 _17606_ (.A(_03670_),
    .B(_03087_),
    .C(_03697_),
    .X(_03709_));
 sky130_fd_sc_hd__a31o_1 _17607_ (.A1(_03696_),
    .A2(net1888),
    .A3(_03672_),
    .B1(_03709_),
    .X(_02462_));
 sky130_fd_sc_hd__nand2_1 _17608_ (.A(_03541_),
    .B(net4104),
    .Y(_03710_));
 sky130_fd_sc_hd__a22o_1 _17609_ (.A1(_03671_),
    .A2(_03710_),
    .B1(_03679_),
    .B2(_10335_),
    .X(_03711_));
 sky130_fd_sc_hd__inv_2 _17610_ (.A(_03711_),
    .Y(_02463_));
 sky130_fd_sc_hd__nand2_1 _17611_ (.A(_03541_),
    .B(net4036),
    .Y(_03712_));
 sky130_fd_sc_hd__a22o_1 _17612_ (.A1(_03671_),
    .A2(_03712_),
    .B1(_03679_),
    .B2(_09495_),
    .X(_03713_));
 sky130_fd_sc_hd__inv_2 _17613_ (.A(_03713_),
    .Y(_02448_));
 sky130_fd_sc_hd__nor2_1 _17614_ (.A(_03605_),
    .B(_03673_),
    .Y(_03714_));
 sky130_fd_sc_hd__a31o_1 _17615_ (.A1(_03696_),
    .A2(net1688),
    .A3(_03672_),
    .B1(_03714_),
    .X(_02449_));
 sky130_fd_sc_hd__and3_1 _17616_ (.A(_03670_),
    .B(_03199_),
    .C(_03697_),
    .X(_03715_));
 sky130_fd_sc_hd__a31o_1 _17617_ (.A1(_03696_),
    .A2(net1801),
    .A3(_03673_),
    .B1(_03715_),
    .X(_02450_));
 sky130_fd_sc_hd__nand2_1 _17618_ (.A(_03541_),
    .B(net3924),
    .Y(_03716_));
 sky130_fd_sc_hd__a22o_1 _17619_ (.A1(_03671_),
    .A2(_03716_),
    .B1(_03679_),
    .B2(_10342_),
    .X(_03717_));
 sky130_fd_sc_hd__inv_2 _17620_ (.A(_03717_),
    .Y(_02451_));
 sky130_fd_sc_hd__and3_1 _17621_ (.A(_03670_),
    .B(_03550_),
    .C(_03697_),
    .X(_03718_));
 sky130_fd_sc_hd__a31o_1 _17622_ (.A1(_03696_),
    .A2(net1361),
    .A3(_03673_),
    .B1(_03718_),
    .X(_02452_));
 sky130_fd_sc_hd__and3_1 _17623_ (.A(_03670_),
    .B(_11426_),
    .C(_03697_),
    .X(_03719_));
 sky130_fd_sc_hd__a31o_1 _17624_ (.A1(_03696_),
    .A2(net1119),
    .A3(_03673_),
    .B1(_03719_),
    .X(_02453_));
 sky130_fd_sc_hd__nand2_1 _17625_ (.A(_03644_),
    .B(net3159),
    .Y(_03720_));
 sky130_fd_sc_hd__a22o_1 _17626_ (.A1(_09296_),
    .A2(_03670_),
    .B1(_03673_),
    .B2(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__inv_2 _17627_ (.A(_03721_),
    .Y(_02454_));
 sky130_fd_sc_hd__nand2_1 _17628_ (.A(_03644_),
    .B(net3185),
    .Y(_03722_));
 sky130_fd_sc_hd__a22o_1 _17629_ (.A1(_09440_),
    .A2(_03670_),
    .B1(_03673_),
    .B2(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__inv_2 _17630_ (.A(_03723_),
    .Y(_02455_));
 sky130_fd_sc_hd__nor2_4 _17631_ (.A(_03616_),
    .B(_10356_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2_4 _17632_ (.A(_03724_),
    .B(_09225_),
    .Y(_03725_));
 sky130_fd_sc_hd__buf_4 _17633_ (.A(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__nand2_1 _17634_ (.A(_03541_),
    .B(net4170),
    .Y(_03727_));
 sky130_fd_sc_hd__and3_1 _17635_ (.A(_10355_),
    .B(_03677_),
    .C(_08725_),
    .X(_03728_));
 sky130_fd_sc_hd__a22o_1 _17636_ (.A1(_03726_),
    .A2(_03727_),
    .B1(_09451_),
    .B2(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__inv_2 _17637_ (.A(net4171),
    .Y(_02440_));
 sky130_fd_sc_hd__buf_4 _17638_ (.A(_08776_),
    .X(_03730_));
 sky130_fd_sc_hd__nand2_1 _17639_ (.A(_03730_),
    .B(net3926),
    .Y(_03731_));
 sky130_fd_sc_hd__buf_4 _17640_ (.A(_03728_),
    .X(_03732_));
 sky130_fd_sc_hd__a22o_1 _17641_ (.A1(_03726_),
    .A2(_03731_),
    .B1(_03732_),
    .B2(_09315_),
    .X(_03733_));
 sky130_fd_sc_hd__inv_2 _17642_ (.A(_03733_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_1 _17643_ (.A(_03730_),
    .B(net3998),
    .Y(_03734_));
 sky130_fd_sc_hd__a22o_1 _17644_ (.A1(_03726_),
    .A2(_03734_),
    .B1(_03732_),
    .B2(_09460_),
    .X(_03735_));
 sky130_fd_sc_hd__inv_2 _17645_ (.A(_03735_),
    .Y(_02442_));
 sky130_fd_sc_hd__nand2_1 _17646_ (.A(_03730_),
    .B(net4100),
    .Y(_03736_));
 sky130_fd_sc_hd__a22o_1 _17647_ (.A1(_03726_),
    .A2(_03736_),
    .B1(_03732_),
    .B2(_09195_),
    .X(_03737_));
 sky130_fd_sc_hd__inv_2 _17648_ (.A(_03737_),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _17649_ (.A(_03730_),
    .B(net4057),
    .Y(_03738_));
 sky130_fd_sc_hd__a22o_1 _17650_ (.A1(_03726_),
    .A2(_03738_),
    .B1(_03732_),
    .B2(_09201_),
    .X(_03739_));
 sky130_fd_sc_hd__inv_2 _17651_ (.A(_03739_),
    .Y(_02444_));
 sky130_fd_sc_hd__nand2_1 _17652_ (.A(_03730_),
    .B(net3914),
    .Y(_03740_));
 sky130_fd_sc_hd__a22o_1 _17653_ (.A1(_03726_),
    .A2(_03740_),
    .B1(_03732_),
    .B2(_09205_),
    .X(_03741_));
 sky130_fd_sc_hd__inv_2 _17654_ (.A(_03741_),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _17655_ (.A(_03730_),
    .B(net4206),
    .Y(_03742_));
 sky130_fd_sc_hd__a22o_1 _17656_ (.A1(_03726_),
    .A2(_03742_),
    .B1(_03732_),
    .B2(_09398_),
    .X(_03743_));
 sky130_fd_sc_hd__inv_2 _17657_ (.A(_03743_),
    .Y(_02446_));
 sky130_fd_sc_hd__nand2_1 _17658_ (.A(_03730_),
    .B(net4135),
    .Y(_03744_));
 sky130_fd_sc_hd__a22o_1 _17659_ (.A1(_03726_),
    .A2(_03744_),
    .B1(_03732_),
    .B2(_09212_),
    .X(_03745_));
 sky130_fd_sc_hd__inv_2 _17660_ (.A(_03745_),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _17661_ (.A(_03730_),
    .B(net4256),
    .Y(_03746_));
 sky130_fd_sc_hd__a22o_1 _17662_ (.A1(_03726_),
    .A2(_03746_),
    .B1(_03732_),
    .B2(_09531_),
    .X(_03747_));
 sky130_fd_sc_hd__inv_2 _17663_ (.A(_03747_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_1 _17664_ (.A(_03730_),
    .B(net3925),
    .Y(_03748_));
 sky130_fd_sc_hd__a22o_1 _17665_ (.A1(_03726_),
    .A2(_03748_),
    .B1(_03732_),
    .B2(_10313_),
    .X(_03749_));
 sky130_fd_sc_hd__inv_2 _17666_ (.A(_03749_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_1 _17667_ (.A(_03730_),
    .B(net4030),
    .Y(_03750_));
 sky130_fd_sc_hd__a22o_1 _17668_ (.A1(_03725_),
    .A2(_03750_),
    .B1(_03732_),
    .B2(_10316_),
    .X(_03751_));
 sky130_fd_sc_hd__inv_2 _17669_ (.A(_03751_),
    .Y(_02434_));
 sky130_fd_sc_hd__buf_4 _17670_ (.A(_03725_),
    .X(_03752_));
 sky130_fd_sc_hd__nor2_1 _17671_ (.A(_02904_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__a31o_1 _17672_ (.A1(_03696_),
    .A2(net853),
    .A3(_03752_),
    .B1(_03753_),
    .X(_02435_));
 sky130_fd_sc_hd__nand2_1 _17673_ (.A(_03730_),
    .B(net3987),
    .Y(_03754_));
 sky130_fd_sc_hd__a22o_1 _17674_ (.A1(_03725_),
    .A2(_03754_),
    .B1(_03732_),
    .B2(_09593_),
    .X(_03755_));
 sky130_fd_sc_hd__inv_2 _17675_ (.A(_03755_),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _17676_ (.A(_02845_),
    .B(_03752_),
    .Y(_03756_));
 sky130_fd_sc_hd__a31o_1 _17677_ (.A1(_03696_),
    .A2(net899),
    .A3(_03752_),
    .B1(_03756_),
    .X(_02437_));
 sky130_fd_sc_hd__nand2_1 _17678_ (.A(_03730_),
    .B(net4040),
    .Y(_03757_));
 sky130_fd_sc_hd__a22o_1 _17679_ (.A1(_03725_),
    .A2(_03757_),
    .B1(_03732_),
    .B2(_09239_),
    .X(_03758_));
 sky130_fd_sc_hd__inv_2 _17680_ (.A(_03758_),
    .Y(_02438_));
 sky130_fd_sc_hd__nor2_1 _17681_ (.A(_03026_),
    .B(_03752_),
    .Y(_03759_));
 sky130_fd_sc_hd__a31o_1 _17682_ (.A1(_03696_),
    .A2(net1560),
    .A3(_03752_),
    .B1(_03759_),
    .X(_02439_));
 sky130_fd_sc_hd__nor2_1 _17683_ (.A(_03294_),
    .B(_03726_),
    .Y(_03760_));
 sky130_fd_sc_hd__a31o_1 _17684_ (.A1(_03696_),
    .A2(net1552),
    .A3(_03752_),
    .B1(_03760_),
    .X(_02424_));
 sky130_fd_sc_hd__and3_1 _17685_ (.A(_03724_),
    .B(_03029_),
    .C(_03697_),
    .X(_03761_));
 sky130_fd_sc_hd__a31o_1 _17686_ (.A1(_03696_),
    .A2(net2252),
    .A3(_03752_),
    .B1(_03761_),
    .X(_02425_));
 sky130_fd_sc_hd__nor2_1 _17687_ (.A(_03482_),
    .B(_03726_),
    .Y(_03762_));
 sky130_fd_sc_hd__a31o_1 _17688_ (.A1(_03696_),
    .A2(net2139),
    .A3(_03752_),
    .B1(_03762_),
    .X(_02426_));
 sky130_fd_sc_hd__buf_4 _17689_ (.A(_03398_),
    .X(_03763_));
 sky130_fd_sc_hd__and3_1 _17690_ (.A(_03724_),
    .B(_03032_),
    .C(_03697_),
    .X(_03764_));
 sky130_fd_sc_hd__a31o_1 _17691_ (.A1(_03763_),
    .A2(net841),
    .A3(_03752_),
    .B1(_03764_),
    .X(_02427_));
 sky130_fd_sc_hd__nor2_1 _17692_ (.A(_09259_),
    .B(_03726_),
    .Y(_03765_));
 sky130_fd_sc_hd__a31o_1 _17693_ (.A1(_03763_),
    .A2(net983),
    .A3(_03752_),
    .B1(_03765_),
    .X(_02428_));
 sky130_fd_sc_hd__nand2_1 _17694_ (.A(_03730_),
    .B(net4085),
    .Y(_03766_));
 sky130_fd_sc_hd__a22o_1 _17695_ (.A1(_03725_),
    .A2(_03766_),
    .B1(_03732_),
    .B2(_10331_),
    .X(_03767_));
 sky130_fd_sc_hd__inv_2 _17696_ (.A(_03767_),
    .Y(_02429_));
 sky130_fd_sc_hd__and3_1 _17697_ (.A(_03724_),
    .B(_03087_),
    .C(_03697_),
    .X(_03768_));
 sky130_fd_sc_hd__a31o_1 _17698_ (.A1(_03763_),
    .A2(net2410),
    .A3(_03752_),
    .B1(_03768_),
    .X(_02430_));
 sky130_fd_sc_hd__nand2_1 _17699_ (.A(_03730_),
    .B(net4024),
    .Y(_03769_));
 sky130_fd_sc_hd__a22o_1 _17700_ (.A1(_03725_),
    .A2(_03769_),
    .B1(_03732_),
    .B2(_10335_),
    .X(_03770_));
 sky130_fd_sc_hd__inv_2 _17701_ (.A(_03770_),
    .Y(_02431_));
 sky130_fd_sc_hd__and3_1 _17702_ (.A(_03724_),
    .B(_03196_),
    .C(_03697_),
    .X(_03771_));
 sky130_fd_sc_hd__a31o_1 _17703_ (.A1(_03763_),
    .A2(net1063),
    .A3(_03752_),
    .B1(_03771_),
    .X(_02416_));
 sky130_fd_sc_hd__nor2_1 _17704_ (.A(_03605_),
    .B(_03726_),
    .Y(_03772_));
 sky130_fd_sc_hd__a31o_1 _17705_ (.A1(_03763_),
    .A2(net821),
    .A3(_03752_),
    .B1(_03772_),
    .X(_02417_));
 sky130_fd_sc_hd__nand2_1 _17706_ (.A(_03730_),
    .B(net4075),
    .Y(_03773_));
 sky130_fd_sc_hd__a22o_1 _17707_ (.A1(_03725_),
    .A2(_03773_),
    .B1(_03732_),
    .B2(_09280_),
    .X(_03774_));
 sky130_fd_sc_hd__inv_2 _17708_ (.A(_03774_),
    .Y(_02418_));
 sky130_fd_sc_hd__nand2_1 _17709_ (.A(_03730_),
    .B(net4081),
    .Y(_03775_));
 sky130_fd_sc_hd__a22o_1 _17710_ (.A1(_03725_),
    .A2(_03775_),
    .B1(_03732_),
    .B2(_10342_),
    .X(_03776_));
 sky130_fd_sc_hd__inv_2 _17711_ (.A(_03776_),
    .Y(_02419_));
 sky130_fd_sc_hd__and3_1 _17712_ (.A(_03724_),
    .B(_03550_),
    .C(_03697_),
    .X(_03777_));
 sky130_fd_sc_hd__a31o_1 _17713_ (.A1(_03763_),
    .A2(net2427),
    .A3(_03752_),
    .B1(_03777_),
    .X(_02420_));
 sky130_fd_sc_hd__and3_1 _17714_ (.A(_03724_),
    .B(_11426_),
    .C(_03697_),
    .X(_03778_));
 sky130_fd_sc_hd__a31o_1 _17715_ (.A1(_03763_),
    .A2(net883),
    .A3(_03752_),
    .B1(_03778_),
    .X(_02421_));
 sky130_fd_sc_hd__nand2_1 _17716_ (.A(_03644_),
    .B(net3152),
    .Y(_03779_));
 sky130_fd_sc_hd__a22o_1 _17717_ (.A1(_09296_),
    .A2(_03724_),
    .B1(_03726_),
    .B2(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__inv_2 _17718_ (.A(_03780_),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _17719_ (.A(_03644_),
    .B(net3413),
    .Y(_03781_));
 sky130_fd_sc_hd__a22o_1 _17720_ (.A1(_09440_),
    .A2(_03724_),
    .B1(_03726_),
    .B2(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__inv_2 _17721_ (.A(_03782_),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_2 _17722_ (.A(_03616_),
    .B(_10411_),
    .Y(_03783_));
 sky130_fd_sc_hd__inv_2 _17723_ (.A(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__nor2_1 _17724_ (.A(_08727_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__clkinv_4 _17725_ (.A(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__buf_4 _17726_ (.A(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__buf_4 _17727_ (.A(_03786_),
    .X(_03788_));
 sky130_fd_sc_hd__nor2_1 _17728_ (.A(_09180_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__a31o_1 _17729_ (.A1(_03763_),
    .A2(net2416),
    .A3(_03787_),
    .B1(_03789_),
    .X(_02408_));
 sky130_fd_sc_hd__nor2_1 _17730_ (.A(_03170_),
    .B(_03788_),
    .Y(_03790_));
 sky130_fd_sc_hd__a31o_1 _17731_ (.A1(_03763_),
    .A2(net1743),
    .A3(_03787_),
    .B1(_03790_),
    .X(_02409_));
 sky130_fd_sc_hd__nor2_1 _17732_ (.A(_03219_),
    .B(_03788_),
    .Y(_03791_));
 sky130_fd_sc_hd__a31o_1 _17733_ (.A1(_03763_),
    .A2(net1221),
    .A3(_03787_),
    .B1(_03791_),
    .X(_02410_));
 sky130_fd_sc_hd__and3_1 _17734_ (.A(_03783_),
    .B(net69),
    .C(_03697_),
    .X(_03792_));
 sky130_fd_sc_hd__a31o_1 _17735_ (.A1(_03787_),
    .A2(_03629_),
    .A3(net2250),
    .B1(_03792_),
    .X(_02411_));
 sky130_fd_sc_hd__nor2_4 _17736_ (.A(_09190_),
    .B(_03784_),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_1 _17737_ (.A(_03644_),
    .B(net2870),
    .Y(_03794_));
 sky130_fd_sc_hd__a22o_1 _17738_ (.A1(_03793_),
    .A2(_11330_),
    .B1(_03788_),
    .B2(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__inv_2 _17739_ (.A(_03795_),
    .Y(_02412_));
 sky130_fd_sc_hd__and3_1 _17740_ (.A(_03783_),
    .B(_11391_),
    .C(_03697_),
    .X(_03796_));
 sky130_fd_sc_hd__a31o_1 _17741_ (.A1(_03787_),
    .A2(_03629_),
    .A3(net1511),
    .B1(_03796_),
    .X(_02413_));
 sky130_fd_sc_hd__nand2_1 _17742_ (.A(_03644_),
    .B(net3219),
    .Y(_03797_));
 sky130_fd_sc_hd__a22o_1 _17743_ (.A1(_03793_),
    .A2(_11105_),
    .B1(_03786_),
    .B2(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__inv_2 _17744_ (.A(_03798_),
    .Y(_02414_));
 sky130_fd_sc_hd__and3_1 _17745_ (.A(_03783_),
    .B(_10874_),
    .C(_03697_),
    .X(_03799_));
 sky130_fd_sc_hd__a31o_1 _17746_ (.A1(_03787_),
    .A2(_03629_),
    .A3(net1297),
    .B1(_03799_),
    .X(_02415_));
 sky130_fd_sc_hd__nand2_1 _17747_ (.A(_03644_),
    .B(net3631),
    .Y(_03800_));
 sky130_fd_sc_hd__a22o_1 _17748_ (.A1(_03793_),
    .A2(net135),
    .B1(_03786_),
    .B2(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__inv_2 _17749_ (.A(_03801_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand2_1 _17750_ (.A(_03644_),
    .B(net3165),
    .Y(_03802_));
 sky130_fd_sc_hd__a22o_1 _17751_ (.A1(_03793_),
    .A2(_02899_),
    .B1(_03786_),
    .B2(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__inv_2 _17752_ (.A(_03803_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand2_1 _17753_ (.A(_03644_),
    .B(net3250),
    .Y(_03804_));
 sky130_fd_sc_hd__a22o_1 _17754_ (.A1(_03793_),
    .A2(_02963_),
    .B1(_03786_),
    .B2(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__inv_2 _17755_ (.A(_03805_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_1 _17756_ (.A(_02904_),
    .B(_03788_),
    .Y(_03806_));
 sky130_fd_sc_hd__a31o_1 _17757_ (.A1(_03763_),
    .A2(net631),
    .A3(_03787_),
    .B1(_03806_),
    .X(_02403_));
 sky130_fd_sc_hd__nor2_1 _17758_ (.A(_03020_),
    .B(_03788_),
    .Y(_03807_));
 sky130_fd_sc_hd__a31o_1 _17759_ (.A1(_03763_),
    .A2(net2409),
    .A3(_03787_),
    .B1(_03807_),
    .X(_02404_));
 sky130_fd_sc_hd__nor2_1 _17760_ (.A(_02845_),
    .B(_03788_),
    .Y(_03808_));
 sky130_fd_sc_hd__a31o_1 _17761_ (.A1(_03763_),
    .A2(net609),
    .A3(_03787_),
    .B1(_03808_),
    .X(_02405_));
 sky130_fd_sc_hd__buf_4 _17762_ (.A(_11219_),
    .X(_03809_));
 sky130_fd_sc_hd__and3_1 _17763_ (.A(_03783_),
    .B(net64),
    .C(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__a31o_1 _17764_ (.A1(_03787_),
    .A2(_03629_),
    .A3(net1169),
    .B1(_03810_),
    .X(_02406_));
 sky130_fd_sc_hd__nor2_1 _17765_ (.A(_03026_),
    .B(_03788_),
    .Y(_03811_));
 sky130_fd_sc_hd__a31o_1 _17766_ (.A1(_03763_),
    .A2(net653),
    .A3(_03787_),
    .B1(_03811_),
    .X(_02407_));
 sky130_fd_sc_hd__nor2_1 _17767_ (.A(_03294_),
    .B(_03788_),
    .Y(_03812_));
 sky130_fd_sc_hd__a31o_1 _17768_ (.A1(_03763_),
    .A2(net947),
    .A3(_03788_),
    .B1(_03812_),
    .X(_02392_));
 sky130_fd_sc_hd__and3_1 _17769_ (.A(_03783_),
    .B(_03029_),
    .C(_03809_),
    .X(_03813_));
 sky130_fd_sc_hd__a31o_1 _17770_ (.A1(_03787_),
    .A2(_03629_),
    .A3(net1339),
    .B1(_03813_),
    .X(_02393_));
 sky130_fd_sc_hd__nor2_1 _17771_ (.A(_03482_),
    .B(_03788_),
    .Y(_03814_));
 sky130_fd_sc_hd__a31o_1 _17772_ (.A1(_03763_),
    .A2(net839),
    .A3(_03788_),
    .B1(_03814_),
    .X(_02394_));
 sky130_fd_sc_hd__buf_4 _17773_ (.A(_03271_),
    .X(_03815_));
 sky130_fd_sc_hd__nand2_1 _17774_ (.A(_03815_),
    .B(net3208),
    .Y(_03816_));
 sky130_fd_sc_hd__a22o_1 _17775_ (.A1(_03793_),
    .A2(_09255_),
    .B1(_03786_),
    .B2(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__inv_2 _17776_ (.A(_03817_),
    .Y(_02395_));
 sky130_fd_sc_hd__clkbuf_8 _17777_ (.A(_03398_),
    .X(_03818_));
 sky130_fd_sc_hd__nor2_1 _17778_ (.A(_09259_),
    .B(_03788_),
    .Y(_03819_));
 sky130_fd_sc_hd__a31o_1 _17779_ (.A1(_03818_),
    .A2(net879),
    .A3(_03788_),
    .B1(_03819_),
    .X(_02396_));
 sky130_fd_sc_hd__nand2_1 _17780_ (.A(_03815_),
    .B(net3350),
    .Y(_03820_));
 sky130_fd_sc_hd__a22o_1 _17781_ (.A1(_03793_),
    .A2(_02916_),
    .B1(_03786_),
    .B2(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__inv_2 _17782_ (.A(_03821_),
    .Y(_02397_));
 sky130_fd_sc_hd__and3_1 _17783_ (.A(_03783_),
    .B(_03087_),
    .C(_03809_),
    .X(_03822_));
 sky130_fd_sc_hd__a31o_1 _17784_ (.A1(_03787_),
    .A2(_03629_),
    .A3(net1554),
    .B1(_03822_),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_1 _17785_ (.A(_03815_),
    .B(net3605),
    .Y(_03823_));
 sky130_fd_sc_hd__a22o_1 _17786_ (.A1(_03793_),
    .A2(_02921_),
    .B1(_03786_),
    .B2(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__inv_2 _17787_ (.A(_03824_),
    .Y(_02399_));
 sky130_fd_sc_hd__nand2_1 _17788_ (.A(_03815_),
    .B(net3307),
    .Y(_03825_));
 sky130_fd_sc_hd__a22o_1 _17789_ (.A1(_03793_),
    .A2(net141),
    .B1(_03786_),
    .B2(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__inv_2 _17790_ (.A(_03826_),
    .Y(_02384_));
 sky130_fd_sc_hd__nor2_1 _17791_ (.A(_03605_),
    .B(_03788_),
    .Y(_03827_));
 sky130_fd_sc_hd__a31o_1 _17792_ (.A1(_03818_),
    .A2(net1333),
    .A3(_03788_),
    .B1(_03827_),
    .X(_02385_));
 sky130_fd_sc_hd__nand2_1 _17793_ (.A(_03815_),
    .B(net3407),
    .Y(_03828_));
 sky130_fd_sc_hd__a22o_1 _17794_ (.A1(_03793_),
    .A2(_10624_),
    .B1(_03786_),
    .B2(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__inv_2 _17795_ (.A(_03829_),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _17796_ (.A(_03815_),
    .B(net3345),
    .Y(_03830_));
 sky130_fd_sc_hd__a22o_1 _17797_ (.A1(_03793_),
    .A2(_02928_),
    .B1(_03786_),
    .B2(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__inv_2 _17798_ (.A(_03831_),
    .Y(_02387_));
 sky130_fd_sc_hd__nand2_1 _17799_ (.A(_03815_),
    .B(net3271),
    .Y(_03832_));
 sky130_fd_sc_hd__a22o_1 _17800_ (.A1(_03793_),
    .A2(net139),
    .B1(_03786_),
    .B2(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__inv_2 _17801_ (.A(_03833_),
    .Y(_02388_));
 sky130_fd_sc_hd__buf_8 _17802_ (.A(_09222_),
    .X(_03834_));
 sky130_fd_sc_hd__buf_4 _17803_ (.A(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__and3_1 _17804_ (.A(_03783_),
    .B(net78),
    .C(_03809_),
    .X(_03836_));
 sky130_fd_sc_hd__a31o_1 _17805_ (.A1(_03787_),
    .A2(_03835_),
    .A3(net2260),
    .B1(_03836_),
    .X(_02389_));
 sky130_fd_sc_hd__nand2_1 _17806_ (.A(_03317_),
    .B(net3818),
    .Y(_03837_));
 sky130_fd_sc_hd__o2bb2a_1 _17807_ (.A1_N(_03837_),
    .A2_N(_03787_),
    .B1(_02992_),
    .B2(_03784_),
    .X(_02390_));
 sky130_fd_sc_hd__nand2_1 _17808_ (.A(_03317_),
    .B(net3673),
    .Y(_03838_));
 sky130_fd_sc_hd__o2bb2a_1 _17809_ (.A1_N(_03838_),
    .A2_N(_03787_),
    .B1(_11316_),
    .B2(_03784_),
    .X(_02391_));
 sky130_fd_sc_hd__nand2_4 _17810_ (.A(_03163_),
    .B(_09982_),
    .Y(_03839_));
 sky130_fd_sc_hd__nor2_4 _17811_ (.A(_03839_),
    .B(_10469_),
    .Y(_03840_));
 sky130_fd_sc_hd__inv_2 _17812_ (.A(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__nor2_1 _17813_ (.A(_09625_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__inv_2 _17814_ (.A(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__buf_4 _17815_ (.A(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__buf_4 _17816_ (.A(_03843_),
    .X(_03845_));
 sky130_fd_sc_hd__nor2_1 _17817_ (.A(_09180_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__a31o_1 _17818_ (.A1(_03818_),
    .A2(net1115),
    .A3(_03844_),
    .B1(_03846_),
    .X(_02368_));
 sky130_fd_sc_hd__nor2_1 _17819_ (.A(_03170_),
    .B(_03845_),
    .Y(_03847_));
 sky130_fd_sc_hd__a31o_1 _17820_ (.A1(_03818_),
    .A2(net1137),
    .A3(_03844_),
    .B1(_03847_),
    .X(_02369_));
 sky130_fd_sc_hd__nor2_1 _17821_ (.A(_03219_),
    .B(_03845_),
    .Y(_03848_));
 sky130_fd_sc_hd__a31o_1 _17822_ (.A1(_03818_),
    .A2(net2098),
    .A3(_03844_),
    .B1(_03848_),
    .X(_02370_));
 sky130_fd_sc_hd__and3_1 _17823_ (.A(_03840_),
    .B(net69),
    .C(_03809_),
    .X(_03849_));
 sky130_fd_sc_hd__a31o_1 _17824_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net1423),
    .B1(_03849_),
    .X(_02371_));
 sky130_fd_sc_hd__and3_1 _17825_ (.A(_03840_),
    .B(_10586_),
    .C(_03809_),
    .X(_03850_));
 sky130_fd_sc_hd__a31o_1 _17826_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net2279),
    .B1(_03850_),
    .X(_02372_));
 sky130_fd_sc_hd__and3_1 _17827_ (.A(_03840_),
    .B(_11391_),
    .C(_03809_),
    .X(_03851_));
 sky130_fd_sc_hd__a31o_1 _17828_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net1345),
    .B1(_03851_),
    .X(_02373_));
 sky130_fd_sc_hd__nor2_4 _17829_ (.A(_08795_),
    .B(_03841_),
    .Y(_03852_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(_03815_),
    .B(net3632),
    .Y(_03853_));
 sky130_fd_sc_hd__a22o_1 _17831_ (.A1(_03852_),
    .A2(_11105_),
    .B1(_03845_),
    .B2(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__inv_2 _17832_ (.A(_03854_),
    .Y(_02374_));
 sky130_fd_sc_hd__nand2_1 _17833_ (.A(_03815_),
    .B(net3084),
    .Y(_03855_));
 sky130_fd_sc_hd__a22o_1 _17834_ (.A1(_03852_),
    .A2(_10591_),
    .B1(_03845_),
    .B2(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__inv_2 _17835_ (.A(_03856_),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2_1 _17836_ (.A(_03467_),
    .B(_03845_),
    .Y(_03857_));
 sky130_fd_sc_hd__a31o_1 _17837_ (.A1(_03818_),
    .A2(net767),
    .A3(_03845_),
    .B1(_03857_),
    .X(_02360_));
 sky130_fd_sc_hd__nand2_1 _17838_ (.A(_03815_),
    .B(net3494),
    .Y(_03858_));
 sky130_fd_sc_hd__a22o_1 _17839_ (.A1(_03852_),
    .A2(_02899_),
    .B1(_03845_),
    .B2(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__inv_2 _17840_ (.A(_03859_),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_1 _17841_ (.A(_03815_),
    .B(net3557),
    .Y(_03860_));
 sky130_fd_sc_hd__a22o_1 _17842_ (.A1(_03852_),
    .A2(_02963_),
    .B1(_03843_),
    .B2(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__inv_2 _17843_ (.A(_03861_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand2_1 _17844_ (.A(_03815_),
    .B(net3151),
    .Y(_03862_));
 sky130_fd_sc_hd__a22o_1 _17845_ (.A1(_03852_),
    .A2(_09589_),
    .B1(_03843_),
    .B2(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__inv_2 _17846_ (.A(_03863_),
    .Y(_02363_));
 sky130_fd_sc_hd__nor2_1 _17847_ (.A(_03020_),
    .B(_03845_),
    .Y(_03864_));
 sky130_fd_sc_hd__a31o_1 _17848_ (.A1(_03818_),
    .A2(net2009),
    .A3(_03845_),
    .B1(_03864_),
    .X(_02364_));
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(_02845_),
    .B(_03845_),
    .Y(_03865_));
 sky130_fd_sc_hd__a31o_1 _17850_ (.A1(_03818_),
    .A2(net1521),
    .A3(_03845_),
    .B1(_03865_),
    .X(_02365_));
 sky130_fd_sc_hd__and3_1 _17851_ (.A(_03840_),
    .B(net64),
    .C(_03809_),
    .X(_03866_));
 sky130_fd_sc_hd__a31o_1 _17852_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net2365),
    .B1(_03866_),
    .X(_02366_));
 sky130_fd_sc_hd__nand2_1 _17853_ (.A(_03815_),
    .B(net3786),
    .Y(_03867_));
 sky130_fd_sc_hd__a22o_1 _17854_ (.A1(_03852_),
    .A2(_09767_),
    .B1(_03843_),
    .B2(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__inv_2 _17855_ (.A(_03868_),
    .Y(_02367_));
 sky130_fd_sc_hd__nand2_1 _17856_ (.A(_03815_),
    .B(net3553),
    .Y(_03869_));
 sky130_fd_sc_hd__a22o_1 _17857_ (.A1(_03852_),
    .A2(net138),
    .B1(_03843_),
    .B2(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__inv_2 _17858_ (.A(_03870_),
    .Y(_02352_));
 sky130_fd_sc_hd__and3_1 _17859_ (.A(_03840_),
    .B(_03029_),
    .C(_03809_),
    .X(_03871_));
 sky130_fd_sc_hd__a31o_1 _17860_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net2166),
    .B1(_03871_),
    .X(_02353_));
 sky130_fd_sc_hd__nor2_1 _17861_ (.A(_03482_),
    .B(_03845_),
    .Y(_03872_));
 sky130_fd_sc_hd__a31o_1 _17862_ (.A1(_03818_),
    .A2(net1099),
    .A3(_03845_),
    .B1(_03872_),
    .X(_02354_));
 sky130_fd_sc_hd__and3_1 _17863_ (.A(_03840_),
    .B(_03032_),
    .C(_03809_),
    .X(_03873_));
 sky130_fd_sc_hd__a31o_1 _17864_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net2247),
    .B1(_03873_),
    .X(_02355_));
 sky130_fd_sc_hd__nand2_1 _17865_ (.A(_03815_),
    .B(net3439),
    .Y(_03874_));
 sky130_fd_sc_hd__a22o_1 _17866_ (.A1(_03852_),
    .A2(_11136_),
    .B1(_03843_),
    .B2(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__inv_2 _17867_ (.A(_03875_),
    .Y(_02356_));
 sky130_fd_sc_hd__nand2_1 _17868_ (.A(_03815_),
    .B(net3070),
    .Y(_03876_));
 sky130_fd_sc_hd__a22o_1 _17869_ (.A1(_03852_),
    .A2(_02916_),
    .B1(_03843_),
    .B2(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__inv_2 _17870_ (.A(_03877_),
    .Y(_02357_));
 sky130_fd_sc_hd__and3_1 _17871_ (.A(_03840_),
    .B(_03087_),
    .C(_03809_),
    .X(_03878_));
 sky130_fd_sc_hd__a31o_1 _17872_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net803),
    .B1(_03878_),
    .X(_02358_));
 sky130_fd_sc_hd__clkbuf_8 _17873_ (.A(_03271_),
    .X(_03879_));
 sky130_fd_sc_hd__nand2_1 _17874_ (.A(_03879_),
    .B(net2967),
    .Y(_03880_));
 sky130_fd_sc_hd__a22o_1 _17875_ (.A1(_03852_),
    .A2(_02921_),
    .B1(_03843_),
    .B2(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__inv_2 _17876_ (.A(_03881_),
    .Y(_02359_));
 sky130_fd_sc_hd__and3_1 _17877_ (.A(_03840_),
    .B(_03196_),
    .C(_03809_),
    .X(_03882_));
 sky130_fd_sc_hd__a31o_1 _17878_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net1281),
    .B1(_03882_),
    .X(_02344_));
 sky130_fd_sc_hd__nor2_1 _17879_ (.A(_03605_),
    .B(_03845_),
    .Y(_03883_));
 sky130_fd_sc_hd__a31o_1 _17880_ (.A1(_03818_),
    .A2(net2540),
    .A3(_03845_),
    .B1(_03883_),
    .X(_02345_));
 sky130_fd_sc_hd__and3_1 _17881_ (.A(_03840_),
    .B(_03199_),
    .C(_03809_),
    .X(_03884_));
 sky130_fd_sc_hd__a31o_1 _17882_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net1253),
    .B1(_03884_),
    .X(_02346_));
 sky130_fd_sc_hd__nand2_1 _17883_ (.A(_03879_),
    .B(net3056),
    .Y(_03885_));
 sky130_fd_sc_hd__a22o_1 _17884_ (.A1(_03852_),
    .A2(_02928_),
    .B1(_03843_),
    .B2(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__inv_2 _17885_ (.A(_03886_),
    .Y(_02347_));
 sky130_fd_sc_hd__and3_1 _17886_ (.A(_03840_),
    .B(_03550_),
    .C(_03809_),
    .X(_03887_));
 sky130_fd_sc_hd__a31o_1 _17887_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net1906),
    .B1(_03887_),
    .X(_02348_));
 sky130_fd_sc_hd__and3_1 _17888_ (.A(_03840_),
    .B(net78),
    .C(_03809_),
    .X(_03888_));
 sky130_fd_sc_hd__a31o_1 _17889_ (.A1(_03844_),
    .A2(_03835_),
    .A3(net1763),
    .B1(_03888_),
    .X(_02349_));
 sky130_fd_sc_hd__nand2_1 _17890_ (.A(_03317_),
    .B(net3107),
    .Y(_03889_));
 sky130_fd_sc_hd__o2bb2a_1 _17891_ (.A1_N(_03889_),
    .A2_N(_03844_),
    .B1(_02992_),
    .B2(_03841_),
    .X(_02350_));
 sky130_fd_sc_hd__nand2_1 _17892_ (.A(_03317_),
    .B(net3641),
    .Y(_03890_));
 sky130_fd_sc_hd__o2bb2a_1 _17893_ (.A1_N(_03890_),
    .A2_N(_03844_),
    .B1(_11316_),
    .B2(_03841_),
    .X(_02351_));
 sky130_fd_sc_hd__nor2_4 _17894_ (.A(_03839_),
    .B(_10292_),
    .Y(_03891_));
 sky130_fd_sc_hd__nand2_4 _17895_ (.A(_03891_),
    .B(_10413_),
    .Y(_03892_));
 sky130_fd_sc_hd__buf_4 _17896_ (.A(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__buf_4 _17897_ (.A(_03892_),
    .X(_03894_));
 sky130_fd_sc_hd__nor2_1 _17898_ (.A(_09180_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__a31o_1 _17899_ (.A1(_03818_),
    .A2(net2533),
    .A3(_03893_),
    .B1(_03895_),
    .X(_02336_));
 sky130_fd_sc_hd__buf_4 _17900_ (.A(_08776_),
    .X(_03896_));
 sky130_fd_sc_hd__nand2_1 _17901_ (.A(_03896_),
    .B(net3973),
    .Y(_03897_));
 sky130_fd_sc_hd__inv_2 _17902_ (.A(_03839_),
    .Y(_03898_));
 sky130_fd_sc_hd__and3_1 _17903_ (.A(_10291_),
    .B(_03898_),
    .C(_08725_),
    .X(_03899_));
 sky130_fd_sc_hd__clkbuf_4 _17904_ (.A(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__a22o_1 _17905_ (.A1(_03894_),
    .A2(_03897_),
    .B1(_03900_),
    .B2(_09315_),
    .X(_03901_));
 sky130_fd_sc_hd__inv_2 _17906_ (.A(_03901_),
    .Y(_02337_));
 sky130_fd_sc_hd__nand2_1 _17907_ (.A(_03896_),
    .B(net3978),
    .Y(_03902_));
 sky130_fd_sc_hd__a22o_1 _17908_ (.A1(_03894_),
    .A2(_03902_),
    .B1(_03900_),
    .B2(_09460_),
    .X(_03903_));
 sky130_fd_sc_hd__inv_2 _17909_ (.A(_03903_),
    .Y(_02338_));
 sky130_fd_sc_hd__and3_1 _17910_ (.A(_03891_),
    .B(net69),
    .C(_03809_),
    .X(_03904_));
 sky130_fd_sc_hd__a31o_1 _17911_ (.A1(_03818_),
    .A2(net2590),
    .A3(_03893_),
    .B1(_03904_),
    .X(_02339_));
 sky130_fd_sc_hd__buf_4 _17912_ (.A(_11219_),
    .X(_03905_));
 sky130_fd_sc_hd__and3_1 _17913_ (.A(_03891_),
    .B(_10586_),
    .C(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__a31o_1 _17914_ (.A1(_03818_),
    .A2(net2199),
    .A3(_03893_),
    .B1(_03906_),
    .X(_02340_));
 sky130_fd_sc_hd__nand2_1 _17915_ (.A(_03896_),
    .B(net3943),
    .Y(_03907_));
 sky130_fd_sc_hd__a22o_1 _17916_ (.A1(_03894_),
    .A2(_03907_),
    .B1(_03900_),
    .B2(_09205_),
    .X(_03908_));
 sky130_fd_sc_hd__inv_2 _17917_ (.A(_03908_),
    .Y(_02341_));
 sky130_fd_sc_hd__nor2_1 _17918_ (.A(_09208_),
    .B(_03894_),
    .Y(_03909_));
 sky130_fd_sc_hd__a31o_1 _17919_ (.A1(_03818_),
    .A2(net1347),
    .A3(_03893_),
    .B1(_03909_),
    .X(_02342_));
 sky130_fd_sc_hd__and3_1 _17920_ (.A(_03891_),
    .B(net74),
    .C(_03905_),
    .X(_03910_));
 sky130_fd_sc_hd__a31o_1 _17921_ (.A1(_03818_),
    .A2(net1171),
    .A3(_03893_),
    .B1(_03910_),
    .X(_02343_));
 sky130_fd_sc_hd__nor2_1 _17922_ (.A(_03467_),
    .B(_03894_),
    .Y(_03911_));
 sky130_fd_sc_hd__a31o_1 _17923_ (.A1(_03818_),
    .A2(net2639),
    .A3(_03893_),
    .B1(_03911_),
    .X(_02328_));
 sky130_fd_sc_hd__nand2_1 _17924_ (.A(_03896_),
    .B(net3964),
    .Y(_03912_));
 sky130_fd_sc_hd__a22o_1 _17925_ (.A1(_03894_),
    .A2(_03912_),
    .B1(_03900_),
    .B2(_09219_),
    .X(_03913_));
 sky130_fd_sc_hd__inv_2 _17926_ (.A(_03913_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _17927_ (.A(_03896_),
    .B(net4162),
    .Y(_03914_));
 sky130_fd_sc_hd__a22o_1 _17928_ (.A1(_03892_),
    .A2(_03914_),
    .B1(_03900_),
    .B2(_09332_),
    .X(_03915_));
 sky130_fd_sc_hd__inv_2 _17929_ (.A(_03915_),
    .Y(_02330_));
 sky130_fd_sc_hd__buf_4 _17930_ (.A(_03398_),
    .X(_03916_));
 sky130_fd_sc_hd__nor2_1 _17931_ (.A(_02904_),
    .B(_03894_),
    .Y(_03917_));
 sky130_fd_sc_hd__a31o_1 _17932_ (.A1(_03916_),
    .A2(net451),
    .A3(_03893_),
    .B1(_03917_),
    .X(_02331_));
 sky130_fd_sc_hd__nand2_1 _17933_ (.A(_03896_),
    .B(net3934),
    .Y(_03918_));
 sky130_fd_sc_hd__a22o_1 _17934_ (.A1(_03892_),
    .A2(_03918_),
    .B1(_03900_),
    .B2(_09593_),
    .X(_03919_));
 sky130_fd_sc_hd__inv_2 _17935_ (.A(_03919_),
    .Y(_02332_));
 sky130_fd_sc_hd__nor2_1 _17936_ (.A(_02845_),
    .B(_03894_),
    .Y(_03920_));
 sky130_fd_sc_hd__a31o_1 _17937_ (.A1(_03916_),
    .A2(net2626),
    .A3(_03893_),
    .B1(_03920_),
    .X(_02333_));
 sky130_fd_sc_hd__nand2_1 _17938_ (.A(_03896_),
    .B(net4064),
    .Y(_03921_));
 sky130_fd_sc_hd__a22o_1 _17939_ (.A1(_03892_),
    .A2(_03921_),
    .B1(_03900_),
    .B2(_09239_),
    .X(_03922_));
 sky130_fd_sc_hd__inv_2 _17940_ (.A(_03922_),
    .Y(_02334_));
 sky130_fd_sc_hd__nor2_1 _17941_ (.A(_03026_),
    .B(_03894_),
    .Y(_03923_));
 sky130_fd_sc_hd__a31o_1 _17942_ (.A1(_03916_),
    .A2(net2130),
    .A3(_03893_),
    .B1(_03923_),
    .X(_02335_));
 sky130_fd_sc_hd__nor2_1 _17943_ (.A(_03294_),
    .B(_03894_),
    .Y(_03924_));
 sky130_fd_sc_hd__a31o_1 _17944_ (.A1(_03916_),
    .A2(net2643),
    .A3(_03893_),
    .B1(_03924_),
    .X(_02320_));
 sky130_fd_sc_hd__and3_1 _17945_ (.A(_03891_),
    .B(_03029_),
    .C(_03905_),
    .X(_03925_));
 sky130_fd_sc_hd__a31o_1 _17946_ (.A1(_03916_),
    .A2(net2123),
    .A3(_03893_),
    .B1(_03925_),
    .X(_02321_));
 sky130_fd_sc_hd__nand2_1 _17947_ (.A(_03896_),
    .B(net4126),
    .Y(_03926_));
 sky130_fd_sc_hd__a22o_1 _17948_ (.A1(_03892_),
    .A2(_03926_),
    .B1(_03900_),
    .B2(_09348_),
    .X(_03927_));
 sky130_fd_sc_hd__inv_2 _17949_ (.A(_03927_),
    .Y(_02322_));
 sky130_fd_sc_hd__and3_1 _17950_ (.A(_03891_),
    .B(_03032_),
    .C(_03905_),
    .X(_03928_));
 sky130_fd_sc_hd__a31o_1 _17951_ (.A1(_03916_),
    .A2(net1323),
    .A3(_03893_),
    .B1(_03928_),
    .X(_02323_));
 sky130_fd_sc_hd__nand2_1 _17952_ (.A(_03896_),
    .B(net4029),
    .Y(_03929_));
 sky130_fd_sc_hd__a22o_1 _17953_ (.A1(_03892_),
    .A2(_03929_),
    .B1(_03900_),
    .B2(_09354_),
    .X(_03930_));
 sky130_fd_sc_hd__inv_2 _17954_ (.A(_03930_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_1 _17955_ (.A(_03896_),
    .B(net4149),
    .Y(_03931_));
 sky130_fd_sc_hd__a22o_1 _17956_ (.A1(_03892_),
    .A2(_03931_),
    .B1(_03900_),
    .B2(_09263_),
    .X(_03932_));
 sky130_fd_sc_hd__inv_2 _17957_ (.A(_03932_),
    .Y(_02325_));
 sky130_fd_sc_hd__and3_1 _17958_ (.A(_03891_),
    .B(_03087_),
    .C(_03905_),
    .X(_03933_));
 sky130_fd_sc_hd__a31o_1 _17959_ (.A1(_03916_),
    .A2(net1564),
    .A3(_03893_),
    .B1(_03933_),
    .X(_02326_));
 sky130_fd_sc_hd__nand2_1 _17960_ (.A(_03896_),
    .B(net4208),
    .Y(_03934_));
 sky130_fd_sc_hd__a22o_1 _17961_ (.A1(_03892_),
    .A2(_03934_),
    .B1(_03900_),
    .B2(_09269_),
    .X(_03935_));
 sky130_fd_sc_hd__inv_2 _17962_ (.A(_03935_),
    .Y(_02327_));
 sky130_fd_sc_hd__nand2_1 _17963_ (.A(_03896_),
    .B(net4093),
    .Y(_03936_));
 sky130_fd_sc_hd__a22o_1 _17964_ (.A1(_03892_),
    .A2(_03936_),
    .B1(_03900_),
    .B2(_09495_),
    .X(_03937_));
 sky130_fd_sc_hd__inv_2 _17965_ (.A(_03937_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _17966_ (.A(_03605_),
    .B(_03894_),
    .Y(_03938_));
 sky130_fd_sc_hd__a31o_1 _17967_ (.A1(_03916_),
    .A2(net2415),
    .A3(_03893_),
    .B1(_03938_),
    .X(_02313_));
 sky130_fd_sc_hd__and3_1 _17968_ (.A(_03891_),
    .B(_03199_),
    .C(_03905_),
    .X(_03939_));
 sky130_fd_sc_hd__a31o_1 _17969_ (.A1(_03916_),
    .A2(net2206),
    .A3(_03893_),
    .B1(_03939_),
    .X(_02314_));
 sky130_fd_sc_hd__nand2_1 _17970_ (.A(_03896_),
    .B(net4291),
    .Y(_03940_));
 sky130_fd_sc_hd__a22o_1 _17971_ (.A1(_03892_),
    .A2(_03940_),
    .B1(_03900_),
    .B2(_09284_),
    .X(_03941_));
 sky130_fd_sc_hd__inv_2 _17972_ (.A(_03941_),
    .Y(_02315_));
 sky130_fd_sc_hd__and3_1 _17973_ (.A(_03891_),
    .B(_03550_),
    .C(_03905_),
    .X(_03942_));
 sky130_fd_sc_hd__a31o_1 _17974_ (.A1(_03916_),
    .A2(net2608),
    .A3(_03893_),
    .B1(_03942_),
    .X(_02316_));
 sky130_fd_sc_hd__and3_1 _17975_ (.A(_03891_),
    .B(net78),
    .C(_03905_),
    .X(_03943_));
 sky130_fd_sc_hd__a31o_1 _17976_ (.A1(_03916_),
    .A2(net973),
    .A3(_03894_),
    .B1(_03943_),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_1 _17977_ (.A(_03879_),
    .B(net3253),
    .Y(_03944_));
 sky130_fd_sc_hd__a22o_1 _17978_ (.A1(_09296_),
    .A2(_03891_),
    .B1(_03894_),
    .B2(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__inv_2 _17979_ (.A(net3254),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_1 _17980_ (.A(_09299_),
    .B(_03894_),
    .Y(_03946_));
 sky130_fd_sc_hd__a31o_1 _17981_ (.A1(_03916_),
    .A2(net1501),
    .A3(_03894_),
    .B1(_03946_),
    .X(_02319_));
 sky130_fd_sc_hd__nor2_4 _17982_ (.A(_03839_),
    .B(_10356_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_4 _17983_ (.A(_03947_),
    .B(_09225_),
    .Y(_03948_));
 sky130_fd_sc_hd__buf_4 _17984_ (.A(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__nand2_1 _17985_ (.A(_03896_),
    .B(net3985),
    .Y(_03950_));
 sky130_fd_sc_hd__and3_1 _17986_ (.A(_10355_),
    .B(_03898_),
    .C(_08725_),
    .X(_03951_));
 sky130_fd_sc_hd__buf_4 _17987_ (.A(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__a22o_1 _17988_ (.A1(_03949_),
    .A2(_03950_),
    .B1(_09451_),
    .B2(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__inv_2 _17989_ (.A(_03953_),
    .Y(_02304_));
 sky130_fd_sc_hd__buf_4 _17990_ (.A(_03948_),
    .X(_03954_));
 sky130_fd_sc_hd__nor2_1 _17991_ (.A(_03170_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__a31o_1 _17992_ (.A1(_03916_),
    .A2(net599),
    .A3(_03954_),
    .B1(_03955_),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_1 _17993_ (.A(_03219_),
    .B(_03949_),
    .Y(_03956_));
 sky130_fd_sc_hd__a31o_1 _17994_ (.A1(_03916_),
    .A2(net831),
    .A3(_03954_),
    .B1(_03956_),
    .X(_02306_));
 sky130_fd_sc_hd__nand2_1 _17995_ (.A(_03896_),
    .B(net3936),
    .Y(_03957_));
 sky130_fd_sc_hd__a22o_1 _17996_ (.A1(_03949_),
    .A2(_03957_),
    .B1(_03952_),
    .B2(_09195_),
    .X(_03958_));
 sky130_fd_sc_hd__inv_2 _17997_ (.A(_03958_),
    .Y(_02307_));
 sky130_fd_sc_hd__and3_1 _17998_ (.A(_03947_),
    .B(_10586_),
    .C(_03905_),
    .X(_03959_));
 sky130_fd_sc_hd__a31o_1 _17999_ (.A1(_03916_),
    .A2(net781),
    .A3(_03954_),
    .B1(_03959_),
    .X(_02308_));
 sky130_fd_sc_hd__nand2_1 _18000_ (.A(_03896_),
    .B(net4167),
    .Y(_03960_));
 sky130_fd_sc_hd__a22o_1 _18001_ (.A1(_03949_),
    .A2(_03960_),
    .B1(_03952_),
    .B2(_09205_),
    .X(_03961_));
 sky130_fd_sc_hd__inv_2 _18002_ (.A(_03961_),
    .Y(_02309_));
 sky130_fd_sc_hd__nor2_1 _18003_ (.A(_09208_),
    .B(_03949_),
    .Y(_03962_));
 sky130_fd_sc_hd__a31o_1 _18004_ (.A1(_03916_),
    .A2(net1431),
    .A3(_03954_),
    .B1(_03962_),
    .X(_02310_));
 sky130_fd_sc_hd__buf_4 _18005_ (.A(_09164_),
    .X(_03963_));
 sky130_fd_sc_hd__and3_1 _18006_ (.A(_03947_),
    .B(net74),
    .C(_03905_),
    .X(_03964_));
 sky130_fd_sc_hd__a31o_1 _18007_ (.A1(_03963_),
    .A2(net1577),
    .A3(_03954_),
    .B1(_03964_),
    .X(_02311_));
 sky130_fd_sc_hd__nand2_1 _18008_ (.A(_10707_),
    .B(net4121),
    .Y(_03965_));
 sky130_fd_sc_hd__a22o_1 _18009_ (.A1(_03949_),
    .A2(_03965_),
    .B1(_03952_),
    .B2(_09531_),
    .X(_03966_));
 sky130_fd_sc_hd__inv_2 _18010_ (.A(_03966_),
    .Y(_02296_));
 sky130_fd_sc_hd__nand2_1 _18011_ (.A(_10707_),
    .B(net4052),
    .Y(_03967_));
 sky130_fd_sc_hd__a22o_1 _18012_ (.A1(_03949_),
    .A2(_03967_),
    .B1(_03952_),
    .B2(_09219_),
    .X(_03968_));
 sky130_fd_sc_hd__inv_2 _18013_ (.A(_03968_),
    .Y(_02297_));
 sky130_fd_sc_hd__nand2_1 _18014_ (.A(_10707_),
    .B(net4090),
    .Y(_03969_));
 sky130_fd_sc_hd__a22o_1 _18015_ (.A1(_03949_),
    .A2(_03969_),
    .B1(_03952_),
    .B2(_09332_),
    .X(_03970_));
 sky130_fd_sc_hd__inv_2 _18016_ (.A(_03970_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _18017_ (.A(_02904_),
    .B(_03949_),
    .Y(_03971_));
 sky130_fd_sc_hd__a31o_1 _18018_ (.A1(_03963_),
    .A2(net905),
    .A3(_03954_),
    .B1(_03971_),
    .X(_02299_));
 sky130_fd_sc_hd__nand2_1 _18019_ (.A(_10707_),
    .B(net3938),
    .Y(_03972_));
 sky130_fd_sc_hd__a22o_1 _18020_ (.A1(_03948_),
    .A2(_03972_),
    .B1(_03952_),
    .B2(_09593_),
    .X(_03973_));
 sky130_fd_sc_hd__inv_2 _18021_ (.A(_03973_),
    .Y(_02300_));
 sky130_fd_sc_hd__nand2_1 _18022_ (.A(_10707_),
    .B(net4220),
    .Y(_03974_));
 sky130_fd_sc_hd__a22o_1 _18023_ (.A1(_03948_),
    .A2(_03974_),
    .B1(_03952_),
    .B2(_09338_),
    .X(_03975_));
 sky130_fd_sc_hd__inv_2 _18024_ (.A(_03975_),
    .Y(_02301_));
 sky130_fd_sc_hd__and3_1 _18025_ (.A(_03947_),
    .B(net64),
    .C(_03905_),
    .X(_03976_));
 sky130_fd_sc_hd__a31o_1 _18026_ (.A1(_03963_),
    .A2(net913),
    .A3(_03954_),
    .B1(_03976_),
    .X(_02302_));
 sky130_fd_sc_hd__nor2_1 _18027_ (.A(_03026_),
    .B(_03949_),
    .Y(_03977_));
 sky130_fd_sc_hd__a31o_1 _18028_ (.A1(_03963_),
    .A2(net1343),
    .A3(_03954_),
    .B1(_03977_),
    .X(_02303_));
 sky130_fd_sc_hd__nor2_1 _18029_ (.A(_03294_),
    .B(_03949_),
    .Y(_03978_));
 sky130_fd_sc_hd__a31o_1 _18030_ (.A1(_03963_),
    .A2(net751),
    .A3(_03954_),
    .B1(_03978_),
    .X(_02280_));
 sky130_fd_sc_hd__nand2_1 _18031_ (.A(_10707_),
    .B(net4068),
    .Y(_03979_));
 sky130_fd_sc_hd__a22o_1 _18032_ (.A1(_03948_),
    .A2(_03979_),
    .B1(_03952_),
    .B2(_09249_),
    .X(_03980_));
 sky130_fd_sc_hd__inv_2 _18033_ (.A(_03980_),
    .Y(_02281_));
 sky130_fd_sc_hd__nor2_1 _18034_ (.A(_03482_),
    .B(_03949_),
    .Y(_03981_));
 sky130_fd_sc_hd__a31o_1 _18035_ (.A1(_03963_),
    .A2(net989),
    .A3(_03954_),
    .B1(_03981_),
    .X(_02282_));
 sky130_fd_sc_hd__and3_1 _18036_ (.A(_03947_),
    .B(_03032_),
    .C(_03905_),
    .X(_03982_));
 sky130_fd_sc_hd__a31o_1 _18037_ (.A1(_03963_),
    .A2(net649),
    .A3(_03954_),
    .B1(_03982_),
    .X(_02283_));
 sky130_fd_sc_hd__nor2_1 _18038_ (.A(_09259_),
    .B(_03949_),
    .Y(_03983_));
 sky130_fd_sc_hd__a31o_1 _18039_ (.A1(_03963_),
    .A2(net869),
    .A3(_03954_),
    .B1(_03983_),
    .X(_02284_));
 sky130_fd_sc_hd__nand2_1 _18040_ (.A(_10707_),
    .B(net4083),
    .Y(_03984_));
 sky130_fd_sc_hd__a22o_1 _18041_ (.A1(_03948_),
    .A2(_03984_),
    .B1(_03952_),
    .B2(_09263_),
    .X(_03985_));
 sky130_fd_sc_hd__inv_2 _18042_ (.A(_03985_),
    .Y(_02285_));
 sky130_fd_sc_hd__and3_1 _18043_ (.A(_03947_),
    .B(_03087_),
    .C(_03905_),
    .X(_03986_));
 sky130_fd_sc_hd__a31o_1 _18044_ (.A1(_03963_),
    .A2(net2220),
    .A3(_03954_),
    .B1(_03986_),
    .X(_02286_));
 sky130_fd_sc_hd__nand2_1 _18045_ (.A(_10707_),
    .B(net4284),
    .Y(_03987_));
 sky130_fd_sc_hd__a22o_1 _18046_ (.A1(_03948_),
    .A2(_03987_),
    .B1(_03952_),
    .B2(_09269_),
    .X(_03988_));
 sky130_fd_sc_hd__inv_2 _18047_ (.A(_03988_),
    .Y(_02287_));
 sky130_fd_sc_hd__and3_1 _18048_ (.A(_03947_),
    .B(_03196_),
    .C(_03905_),
    .X(_03989_));
 sky130_fd_sc_hd__a31o_1 _18049_ (.A1(_03963_),
    .A2(net675),
    .A3(_03954_),
    .B1(_03989_),
    .X(_02272_));
 sky130_fd_sc_hd__nor2_1 _18050_ (.A(_03605_),
    .B(_03949_),
    .Y(_03990_));
 sky130_fd_sc_hd__a31o_1 _18051_ (.A1(_03963_),
    .A2(net2358),
    .A3(_03954_),
    .B1(_03990_),
    .X(_02273_));
 sky130_fd_sc_hd__nand2_1 _18052_ (.A(_10707_),
    .B(net4046),
    .Y(_03991_));
 sky130_fd_sc_hd__a22o_1 _18053_ (.A1(_03948_),
    .A2(_03991_),
    .B1(_03952_),
    .B2(_09280_),
    .X(_03992_));
 sky130_fd_sc_hd__inv_2 _18054_ (.A(_03992_),
    .Y(_02274_));
 sky130_fd_sc_hd__nand2_1 _18055_ (.A(_10707_),
    .B(net4227),
    .Y(_03993_));
 sky130_fd_sc_hd__a22o_1 _18056_ (.A1(_03948_),
    .A2(_03993_),
    .B1(_03952_),
    .B2(_09284_),
    .X(_03994_));
 sky130_fd_sc_hd__inv_2 _18057_ (.A(_03994_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_1 _18058_ (.A(_10707_),
    .B(net4084),
    .Y(_03995_));
 sky130_fd_sc_hd__a22o_1 _18059_ (.A1(_03948_),
    .A2(_03995_),
    .B1(_03952_),
    .B2(_09288_),
    .X(_03996_));
 sky130_fd_sc_hd__inv_2 _18060_ (.A(_03996_),
    .Y(_02276_));
 sky130_fd_sc_hd__nand2_1 _18061_ (.A(_10707_),
    .B(net4102),
    .Y(_03997_));
 sky130_fd_sc_hd__a22o_1 _18062_ (.A1(_03948_),
    .A2(_03997_),
    .B1(_03952_),
    .B2(net136),
    .X(_03998_));
 sky130_fd_sc_hd__inv_2 _18063_ (.A(_03998_),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _18064_ (.A(_03879_),
    .B(net3415),
    .Y(_03999_));
 sky130_fd_sc_hd__a22o_1 _18065_ (.A1(_09296_),
    .A2(_03947_),
    .B1(_03949_),
    .B2(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__inv_2 _18066_ (.A(net3416),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_1 _18067_ (.A(_03879_),
    .B(net3231),
    .Y(_04001_));
 sky130_fd_sc_hd__a22o_1 _18068_ (.A1(_09440_),
    .A2(_03947_),
    .B1(_03949_),
    .B2(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__inv_2 _18069_ (.A(net3232),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_2 _18070_ (.A(_03839_),
    .B(_10411_),
    .Y(_04003_));
 sky130_fd_sc_hd__inv_2 _18071_ (.A(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__nor2_1 _18072_ (.A(_09625_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__inv_2 _18073_ (.A(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__buf_4 _18074_ (.A(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__buf_4 _18075_ (.A(_04006_),
    .X(_04008_));
 sky130_fd_sc_hd__nor2_1 _18076_ (.A(_09180_),
    .B(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__a31o_1 _18077_ (.A1(_03963_),
    .A2(net773),
    .A3(_04007_),
    .B1(_04009_),
    .X(_02264_));
 sky130_fd_sc_hd__nor2_8 _18078_ (.A(_08797_),
    .B(_04004_),
    .Y(_04010_));
 sky130_fd_sc_hd__nand2_1 _18079_ (.A(_03879_),
    .B(net3142),
    .Y(_04011_));
 sky130_fd_sc_hd__a22o_1 _18080_ (.A1(_04010_),
    .A2(_09314_),
    .B1(_04008_),
    .B2(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__inv_2 _18081_ (.A(_04012_),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(_03879_),
    .B(net3773),
    .Y(_04013_));
 sky130_fd_sc_hd__a22o_1 _18083_ (.A1(_04010_),
    .A2(_09459_),
    .B1(_04008_),
    .B2(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__inv_2 _18084_ (.A(_04014_),
    .Y(_02266_));
 sky130_fd_sc_hd__and3_1 _18085_ (.A(_04003_),
    .B(net69),
    .C(_03905_),
    .X(_04015_));
 sky130_fd_sc_hd__a31o_1 _18086_ (.A1(_04007_),
    .A2(_03835_),
    .A3(net2094),
    .B1(_04015_),
    .X(_02267_));
 sky130_fd_sc_hd__nand2_1 _18087_ (.A(_03879_),
    .B(net3218),
    .Y(_04016_));
 sky130_fd_sc_hd__a22o_1 _18088_ (.A1(_04010_),
    .A2(_11330_),
    .B1(_04008_),
    .B2(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__inv_2 _18089_ (.A(_04017_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand2_1 _18090_ (.A(_03879_),
    .B(net2862),
    .Y(_04018_));
 sky130_fd_sc_hd__a22o_1 _18091_ (.A1(_04010_),
    .A2(_10869_),
    .B1(_04008_),
    .B2(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__inv_2 _18092_ (.A(_04019_),
    .Y(_02269_));
 sky130_fd_sc_hd__nor2_1 _18093_ (.A(_09208_),
    .B(_04008_),
    .Y(_04020_));
 sky130_fd_sc_hd__a31o_1 _18094_ (.A1(_03963_),
    .A2(net1550),
    .A3(_04007_),
    .B1(_04020_),
    .X(_02270_));
 sky130_fd_sc_hd__and3_1 _18095_ (.A(_04003_),
    .B(net74),
    .C(_03905_),
    .X(_04021_));
 sky130_fd_sc_hd__a31o_1 _18096_ (.A1(_04007_),
    .A2(_03835_),
    .A3(net1934),
    .B1(_04021_),
    .X(_02271_));
 sky130_fd_sc_hd__nand2_1 _18097_ (.A(_03879_),
    .B(net3278),
    .Y(_04022_));
 sky130_fd_sc_hd__a22o_1 _18098_ (.A1(_04010_),
    .A2(_09530_),
    .B1(_04008_),
    .B2(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__inv_2 _18099_ (.A(_04023_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand2_1 _18100_ (.A(_03879_),
    .B(net3110),
    .Y(_04024_));
 sky130_fd_sc_hd__a22o_1 _18101_ (.A1(_04010_),
    .A2(_02899_),
    .B1(_04008_),
    .B2(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__inv_2 _18102_ (.A(_04025_),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_1 _18103_ (.A(_03879_),
    .B(net3032),
    .Y(_04026_));
 sky130_fd_sc_hd__a22o_1 _18104_ (.A1(_04010_),
    .A2(_02963_),
    .B1(_04008_),
    .B2(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__inv_2 _18105_ (.A(_04027_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _18106_ (.A(_02904_),
    .B(_04008_),
    .Y(_04028_));
 sky130_fd_sc_hd__a31o_1 _18107_ (.A1(_03963_),
    .A2(net1095),
    .A3(_04007_),
    .B1(_04028_),
    .X(_02259_));
 sky130_fd_sc_hd__nor2_1 _18108_ (.A(_03020_),
    .B(_04008_),
    .Y(_04029_));
 sky130_fd_sc_hd__a31o_1 _18109_ (.A1(_03963_),
    .A2(net959),
    .A3(_04007_),
    .B1(_04029_),
    .X(_02260_));
 sky130_fd_sc_hd__nor2_1 _18110_ (.A(_02845_),
    .B(_04008_),
    .Y(_04030_));
 sky130_fd_sc_hd__a31o_1 _18111_ (.A1(_03963_),
    .A2(net895),
    .A3(_04007_),
    .B1(_04030_),
    .X(_02261_));
 sky130_fd_sc_hd__nand2_1 _18112_ (.A(_03879_),
    .B(net3031),
    .Y(_04031_));
 sky130_fd_sc_hd__a22o_1 _18113_ (.A1(_04010_),
    .A2(_10202_),
    .B1(_04006_),
    .B2(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__inv_2 _18114_ (.A(_04032_),
    .Y(_02262_));
 sky130_fd_sc_hd__clkbuf_8 _18115_ (.A(_09164_),
    .X(_04033_));
 sky130_fd_sc_hd__nor2_1 _18116_ (.A(_03026_),
    .B(_04008_),
    .Y(_04034_));
 sky130_fd_sc_hd__a31o_1 _18117_ (.A1(_04033_),
    .A2(net1990),
    .A3(_04007_),
    .B1(_04034_),
    .X(_02263_));
 sky130_fd_sc_hd__nand2_1 _18118_ (.A(_03879_),
    .B(net3274),
    .Y(_04035_));
 sky130_fd_sc_hd__a22o_1 _18119_ (.A1(_04010_),
    .A2(net137),
    .B1(_04006_),
    .B2(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__inv_2 _18120_ (.A(_04036_),
    .Y(_02248_));
 sky130_fd_sc_hd__buf_4 _18121_ (.A(_11219_),
    .X(_04037_));
 sky130_fd_sc_hd__and3_1 _18122_ (.A(_04003_),
    .B(_03029_),
    .C(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__a31o_1 _18123_ (.A1(_04007_),
    .A2(_03835_),
    .A3(net2531),
    .B1(_04038_),
    .X(_02249_));
 sky130_fd_sc_hd__nor2_1 _18124_ (.A(_03482_),
    .B(_04008_),
    .Y(_04039_));
 sky130_fd_sc_hd__a31o_1 _18125_ (.A1(_04033_),
    .A2(net2385),
    .A3(_04007_),
    .B1(_04039_),
    .X(_02250_));
 sky130_fd_sc_hd__and3_1 _18126_ (.A(_04003_),
    .B(_03032_),
    .C(_04037_),
    .X(_04040_));
 sky130_fd_sc_hd__a31o_1 _18127_ (.A1(_04007_),
    .A2(_03835_),
    .A3(net2544),
    .B1(_04040_),
    .X(_02251_));
 sky130_fd_sc_hd__nor2_1 _18128_ (.A(_09259_),
    .B(_04008_),
    .Y(_04041_));
 sky130_fd_sc_hd__a31o_1 _18129_ (.A1(_04033_),
    .A2(net503),
    .A3(_04008_),
    .B1(_04041_),
    .X(_02252_));
 sky130_fd_sc_hd__nand2_1 _18130_ (.A(_03879_),
    .B(net2838),
    .Y(_04042_));
 sky130_fd_sc_hd__a22o_1 _18131_ (.A1(_04010_),
    .A2(_02916_),
    .B1(_04006_),
    .B2(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__inv_2 _18132_ (.A(_04043_),
    .Y(_02253_));
 sky130_fd_sc_hd__buf_4 _18133_ (.A(_03834_),
    .X(_04044_));
 sky130_fd_sc_hd__and3_1 _18134_ (.A(_04003_),
    .B(_03087_),
    .C(_04037_),
    .X(_04045_));
 sky130_fd_sc_hd__a31o_1 _18135_ (.A1(_04007_),
    .A2(_04044_),
    .A3(net2658),
    .B1(_04045_),
    .X(_02254_));
 sky130_fd_sc_hd__nand2_1 _18136_ (.A(_03879_),
    .B(net3187),
    .Y(_04046_));
 sky130_fd_sc_hd__a22o_1 _18137_ (.A1(_04010_),
    .A2(_02921_),
    .B1(_04006_),
    .B2(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__inv_2 _18138_ (.A(_04047_),
    .Y(_02255_));
 sky130_fd_sc_hd__clkbuf_8 _18139_ (.A(_03271_),
    .X(_04048_));
 sky130_fd_sc_hd__nand2_1 _18140_ (.A(_04048_),
    .B(net3368),
    .Y(_04049_));
 sky130_fd_sc_hd__a22o_1 _18141_ (.A1(_04010_),
    .A2(net141),
    .B1(_04006_),
    .B2(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__inv_2 _18142_ (.A(_04050_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_1 _18143_ (.A(_04048_),
    .B(net3364),
    .Y(_04051_));
 sky130_fd_sc_hd__a22o_1 _18144_ (.A1(_04010_),
    .A2(_09365_),
    .B1(_04006_),
    .B2(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__inv_2 _18145_ (.A(_04052_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _18146_ (.A(_04048_),
    .B(net3419),
    .Y(_04053_));
 sky130_fd_sc_hd__a22o_1 _18147_ (.A1(_04010_),
    .A2(_10624_),
    .B1(_04006_),
    .B2(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__inv_2 _18148_ (.A(_04054_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand2_1 _18149_ (.A(_04048_),
    .B(net3066),
    .Y(_04055_));
 sky130_fd_sc_hd__a22o_1 _18150_ (.A1(_04010_),
    .A2(_02928_),
    .B1(_04006_),
    .B2(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__inv_2 _18151_ (.A(_04056_),
    .Y(_02243_));
 sky130_fd_sc_hd__and3_1 _18152_ (.A(_04003_),
    .B(_03550_),
    .C(_04037_),
    .X(_04057_));
 sky130_fd_sc_hd__a31o_1 _18153_ (.A1(_04007_),
    .A2(_04044_),
    .A3(net1684),
    .B1(_04057_),
    .X(_02244_));
 sky130_fd_sc_hd__and3_1 _18154_ (.A(_04003_),
    .B(net78),
    .C(_04037_),
    .X(_04058_));
 sky130_fd_sc_hd__a31o_1 _18155_ (.A1(_04007_),
    .A2(_04044_),
    .A3(net2306),
    .B1(_04058_),
    .X(_02245_));
 sky130_fd_sc_hd__nand2_1 _18156_ (.A(_03317_),
    .B(net3784),
    .Y(_04059_));
 sky130_fd_sc_hd__o2bb2a_1 _18157_ (.A1_N(_04059_),
    .A2_N(_04007_),
    .B1(_02992_),
    .B2(_04004_),
    .X(_02246_));
 sky130_fd_sc_hd__nand2_1 _18158_ (.A(_03317_),
    .B(net3814),
    .Y(_04060_));
 sky130_fd_sc_hd__o2bb2a_1 _18159_ (.A1_N(_04060_),
    .A2_N(_04007_),
    .B1(_11316_),
    .B2(_04004_),
    .X(_02247_));
 sky130_fd_sc_hd__and3_4 _18160_ (.A(_09171_),
    .B(_09443_),
    .C(_09173_),
    .X(_04061_));
 sky130_fd_sc_hd__inv_2 _18161_ (.A(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__nor2_1 _18162_ (.A(_09304_),
    .B(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__clkinv_4 _18163_ (.A(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__buf_4 _18164_ (.A(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__buf_4 _18165_ (.A(_04064_),
    .X(_04066_));
 sky130_fd_sc_hd__nor2_1 _18166_ (.A(_09180_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a31o_1 _18167_ (.A1(_04033_),
    .A2(net2653),
    .A3(_04065_),
    .B1(_04067_),
    .X(_02232_));
 sky130_fd_sc_hd__nor2_4 _18168_ (.A(_08797_),
    .B(_04062_),
    .Y(_04068_));
 sky130_fd_sc_hd__nand2_1 _18169_ (.A(_04048_),
    .B(net3260),
    .Y(_04069_));
 sky130_fd_sc_hd__a22o_1 _18170_ (.A1(_04068_),
    .A2(_09314_),
    .B1(_04066_),
    .B2(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__inv_2 _18171_ (.A(_04070_),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_1 _18172_ (.A(_03219_),
    .B(_04066_),
    .Y(_04071_));
 sky130_fd_sc_hd__a31o_1 _18173_ (.A1(_04033_),
    .A2(net2652),
    .A3(_04065_),
    .B1(_04071_),
    .X(_02234_));
 sky130_fd_sc_hd__and3_1 _18174_ (.A(_04061_),
    .B(net69),
    .C(_04037_),
    .X(_04072_));
 sky130_fd_sc_hd__a31o_1 _18175_ (.A1(_04065_),
    .A2(_04044_),
    .A3(net2650),
    .B1(_04072_),
    .X(_02235_));
 sky130_fd_sc_hd__nand2_1 _18176_ (.A(_04048_),
    .B(net3341),
    .Y(_04073_));
 sky130_fd_sc_hd__a22o_1 _18177_ (.A1(_04068_),
    .A2(_11330_),
    .B1(_04066_),
    .B2(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__inv_2 _18178_ (.A(_04074_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand2_1 _18179_ (.A(_04048_),
    .B(net3579),
    .Y(_04075_));
 sky130_fd_sc_hd__a22o_1 _18180_ (.A1(_04068_),
    .A2(_10869_),
    .B1(_04066_),
    .B2(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__inv_2 _18181_ (.A(_04076_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_1 _18182_ (.A(_04048_),
    .B(net3817),
    .Y(_04077_));
 sky130_fd_sc_hd__a22o_1 _18183_ (.A1(_04068_),
    .A2(_11105_),
    .B1(_04066_),
    .B2(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__inv_2 _18184_ (.A(_04078_),
    .Y(_02238_));
 sky130_fd_sc_hd__nand2_1 _18185_ (.A(_04048_),
    .B(net2978),
    .Y(_04079_));
 sky130_fd_sc_hd__a22o_1 _18186_ (.A1(_04068_),
    .A2(_10591_),
    .B1(_04064_),
    .B2(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__inv_2 _18187_ (.A(_04080_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _18188_ (.A(_03467_),
    .B(_04066_),
    .Y(_04081_));
 sky130_fd_sc_hd__a31o_1 _18189_ (.A1(_04033_),
    .A2(net2108),
    .A3(_04065_),
    .B1(_04081_),
    .X(_02224_));
 sky130_fd_sc_hd__nand2_1 _18190_ (.A(_04048_),
    .B(net3147),
    .Y(_04082_));
 sky130_fd_sc_hd__a22o_1 _18191_ (.A1(_04068_),
    .A2(_02899_),
    .B1(_04064_),
    .B2(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__inv_2 _18192_ (.A(_04083_),
    .Y(_02225_));
 sky130_fd_sc_hd__nand2_1 _18193_ (.A(_04048_),
    .B(net3287),
    .Y(_04084_));
 sky130_fd_sc_hd__a22o_1 _18194_ (.A1(_04068_),
    .A2(_02963_),
    .B1(_04064_),
    .B2(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__inv_2 _18195_ (.A(_04085_),
    .Y(_02226_));
 sky130_fd_sc_hd__nor2_1 _18196_ (.A(_09229_),
    .B(_04066_),
    .Y(_04086_));
 sky130_fd_sc_hd__a31o_1 _18197_ (.A1(_04033_),
    .A2(net953),
    .A3(_04065_),
    .B1(_04086_),
    .X(_02227_));
 sky130_fd_sc_hd__nor2_1 _18198_ (.A(_03020_),
    .B(_04066_),
    .Y(_04087_));
 sky130_fd_sc_hd__a31o_1 _18199_ (.A1(_04033_),
    .A2(net1397),
    .A3(_04065_),
    .B1(_04087_),
    .X(_02228_));
 sky130_fd_sc_hd__nor2_1 _18200_ (.A(_02845_),
    .B(_04066_),
    .Y(_04088_));
 sky130_fd_sc_hd__a31o_1 _18201_ (.A1(_04033_),
    .A2(net1009),
    .A3(_04065_),
    .B1(_04088_),
    .X(_02229_));
 sky130_fd_sc_hd__and3_1 _18202_ (.A(_04061_),
    .B(net64),
    .C(_04037_),
    .X(_04089_));
 sky130_fd_sc_hd__a31o_1 _18203_ (.A1(_04065_),
    .A2(_04044_),
    .A3(net1495),
    .B1(_04089_),
    .X(_02230_));
 sky130_fd_sc_hd__nor2_1 _18204_ (.A(_03026_),
    .B(_04066_),
    .Y(_04090_));
 sky130_fd_sc_hd__a31o_1 _18205_ (.A1(_04033_),
    .A2(net1001),
    .A3(_04065_),
    .B1(_04090_),
    .X(_02231_));
 sky130_fd_sc_hd__nor2_1 _18206_ (.A(_03294_),
    .B(_04066_),
    .Y(_04091_));
 sky130_fd_sc_hd__a31o_1 _18207_ (.A1(_04033_),
    .A2(net2103),
    .A3(_04065_),
    .B1(_04091_),
    .X(_02216_));
 sky130_fd_sc_hd__nand2_1 _18208_ (.A(_04048_),
    .B(net3176),
    .Y(_04092_));
 sky130_fd_sc_hd__a22o_1 _18209_ (.A1(_04068_),
    .A2(_09249_),
    .B1(_04064_),
    .B2(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__inv_2 _18210_ (.A(_04093_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _18211_ (.A(_04048_),
    .B(net3025),
    .Y(_04094_));
 sky130_fd_sc_hd__a22o_1 _18212_ (.A1(_04068_),
    .A2(_09347_),
    .B1(_04064_),
    .B2(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__inv_2 _18213_ (.A(_04095_),
    .Y(_02218_));
 sky130_fd_sc_hd__and3_1 _18214_ (.A(_04061_),
    .B(_03032_),
    .C(_04037_),
    .X(_04096_));
 sky130_fd_sc_hd__a31o_1 _18215_ (.A1(_04065_),
    .A2(_04044_),
    .A3(net2240),
    .B1(_04096_),
    .X(_02219_));
 sky130_fd_sc_hd__nand2_1 _18216_ (.A(_04048_),
    .B(net3486),
    .Y(_04097_));
 sky130_fd_sc_hd__a22o_1 _18217_ (.A1(_04068_),
    .A2(_11136_),
    .B1(_04064_),
    .B2(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__inv_2 _18218_ (.A(_04098_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand2_1 _18219_ (.A(_04048_),
    .B(net3186),
    .Y(_04099_));
 sky130_fd_sc_hd__a22o_1 _18220_ (.A1(_04068_),
    .A2(_02916_),
    .B1(_04064_),
    .B2(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__inv_2 _18221_ (.A(_04100_),
    .Y(_02221_));
 sky130_fd_sc_hd__and3_1 _18222_ (.A(_04061_),
    .B(_03087_),
    .C(_04037_),
    .X(_04101_));
 sky130_fd_sc_hd__a31o_1 _18223_ (.A1(_04065_),
    .A2(_04044_),
    .A3(net1433),
    .B1(_04101_),
    .X(_02222_));
 sky130_fd_sc_hd__nand2_1 _18224_ (.A(_04048_),
    .B(net3356),
    .Y(_04102_));
 sky130_fd_sc_hd__a22o_1 _18225_ (.A1(_04068_),
    .A2(_02921_),
    .B1(_04064_),
    .B2(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__inv_2 _18226_ (.A(_04103_),
    .Y(_02223_));
 sky130_fd_sc_hd__and3_1 _18227_ (.A(_04061_),
    .B(_03196_),
    .C(_04037_),
    .X(_04104_));
 sky130_fd_sc_hd__a31o_1 _18228_ (.A1(_04065_),
    .A2(_04044_),
    .A3(net1955),
    .B1(_04104_),
    .X(_02208_));
 sky130_fd_sc_hd__nor2_1 _18229_ (.A(_03605_),
    .B(_04066_),
    .Y(_04105_));
 sky130_fd_sc_hd__a31o_1 _18230_ (.A1(_04033_),
    .A2(net1970),
    .A3(_04066_),
    .B1(_04105_),
    .X(_02209_));
 sky130_fd_sc_hd__buf_4 _18231_ (.A(_03271_),
    .X(_04106_));
 sky130_fd_sc_hd__nand2_1 _18232_ (.A(_04106_),
    .B(net3500),
    .Y(_04107_));
 sky130_fd_sc_hd__a22o_1 _18233_ (.A1(_04068_),
    .A2(_10624_),
    .B1(_04064_),
    .B2(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__inv_2 _18234_ (.A(_04108_),
    .Y(_02210_));
 sky130_fd_sc_hd__nand2_1 _18235_ (.A(_04106_),
    .B(net3596),
    .Y(_04109_));
 sky130_fd_sc_hd__a22o_1 _18236_ (.A1(_04068_),
    .A2(_02928_),
    .B1(_04064_),
    .B2(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__inv_2 _18237_ (.A(_04110_),
    .Y(_02211_));
 sky130_fd_sc_hd__and3_1 _18238_ (.A(_04061_),
    .B(_03550_),
    .C(_04037_),
    .X(_04111_));
 sky130_fd_sc_hd__a31o_1 _18239_ (.A1(_04065_),
    .A2(_04044_),
    .A3(net2254),
    .B1(_04111_),
    .X(_02212_));
 sky130_fd_sc_hd__and3_1 _18240_ (.A(_04061_),
    .B(net78),
    .C(_04037_),
    .X(_04112_));
 sky130_fd_sc_hd__a31o_1 _18241_ (.A1(_04065_),
    .A2(_04044_),
    .A3(net2291),
    .B1(_04112_),
    .X(_02213_));
 sky130_fd_sc_hd__nand2_1 _18242_ (.A(_03317_),
    .B(net3554),
    .Y(_04113_));
 sky130_fd_sc_hd__o2bb2a_1 _18243_ (.A1_N(_04113_),
    .A2_N(_04065_),
    .B1(_02992_),
    .B2(_04062_),
    .X(_02214_));
 sky130_fd_sc_hd__nor2_1 _18244_ (.A(_09299_),
    .B(_04066_),
    .Y(_04114_));
 sky130_fd_sc_hd__a31o_1 _18245_ (.A1(_04033_),
    .A2(net1883),
    .A3(_04066_),
    .B1(_04114_),
    .X(_02215_));
 sky130_fd_sc_hd__and3_4 _18246_ (.A(_09171_),
    .B(_09444_),
    .C(_09305_),
    .X(_04115_));
 sky130_fd_sc_hd__inv_2 _18247_ (.A(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__nor2_1 _18248_ (.A(_09304_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__inv_2 _18249_ (.A(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__buf_4 _18250_ (.A(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__buf_4 _18251_ (.A(_04118_),
    .X(_04120_));
 sky130_fd_sc_hd__nor2_1 _18252_ (.A(_09180_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__a31o_1 _18253_ (.A1(_04033_),
    .A2(net1093),
    .A3(_04119_),
    .B1(_04121_),
    .X(_02192_));
 sky130_fd_sc_hd__nor2_1 _18254_ (.A(_03170_),
    .B(_04120_),
    .Y(_04122_));
 sky130_fd_sc_hd__a31o_1 _18255_ (.A1(_04033_),
    .A2(net1101),
    .A3(_04119_),
    .B1(_04122_),
    .X(_02193_));
 sky130_fd_sc_hd__nor2_1 _18256_ (.A(_03219_),
    .B(_04120_),
    .Y(_04123_));
 sky130_fd_sc_hd__a31o_1 _18257_ (.A1(_04033_),
    .A2(net1997),
    .A3(_04119_),
    .B1(_04123_),
    .X(_02194_));
 sky130_fd_sc_hd__and3_1 _18258_ (.A(_04115_),
    .B(net69),
    .C(_04037_),
    .X(_04124_));
 sky130_fd_sc_hd__a31o_1 _18259_ (.A1(_04119_),
    .A2(_04044_),
    .A3(net2203),
    .B1(_04124_),
    .X(_02195_));
 sky130_fd_sc_hd__and3_1 _18260_ (.A(_04115_),
    .B(_10586_),
    .C(_04037_),
    .X(_04125_));
 sky130_fd_sc_hd__a31o_1 _18261_ (.A1(_04119_),
    .A2(_04044_),
    .A3(net2090),
    .B1(_04125_),
    .X(_02196_));
 sky130_fd_sc_hd__nor2_4 _18262_ (.A(_09190_),
    .B(_04116_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_1 _18263_ (.A(_04106_),
    .B(net3195),
    .Y(_04127_));
 sky130_fd_sc_hd__a22o_1 _18264_ (.A1(_04126_),
    .A2(_10869_),
    .B1(_04120_),
    .B2(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__inv_2 _18265_ (.A(_04128_),
    .Y(_02197_));
 sky130_fd_sc_hd__buf_4 _18266_ (.A(_09164_),
    .X(_04129_));
 sky130_fd_sc_hd__nor2_1 _18267_ (.A(_09208_),
    .B(_04120_),
    .Y(_04130_));
 sky130_fd_sc_hd__a31o_1 _18268_ (.A1(_04129_),
    .A2(net1535),
    .A3(_04119_),
    .B1(_04130_),
    .X(_02198_));
 sky130_fd_sc_hd__nand2_1 _18269_ (.A(_04106_),
    .B(net3093),
    .Y(_04131_));
 sky130_fd_sc_hd__a22o_1 _18270_ (.A1(_04126_),
    .A2(_10591_),
    .B1(_04120_),
    .B2(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__inv_2 _18271_ (.A(_04132_),
    .Y(_02199_));
 sky130_fd_sc_hd__nor2_1 _18272_ (.A(_03467_),
    .B(_04120_),
    .Y(_04133_));
 sky130_fd_sc_hd__a31o_1 _18273_ (.A1(_04129_),
    .A2(net2364),
    .A3(_04119_),
    .B1(_04133_),
    .X(_02184_));
 sky130_fd_sc_hd__nand2_1 _18274_ (.A(_04106_),
    .B(net3519),
    .Y(_04134_));
 sky130_fd_sc_hd__a22o_1 _18275_ (.A1(_04126_),
    .A2(_02899_),
    .B1(_04118_),
    .B2(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__inv_2 _18276_ (.A(_04135_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand2_1 _18277_ (.A(_04106_),
    .B(net3470),
    .Y(_04136_));
 sky130_fd_sc_hd__a22o_1 _18278_ (.A1(_04126_),
    .A2(_02963_),
    .B1(_04118_),
    .B2(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__inv_2 _18279_ (.A(_04137_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _18280_ (.A(_04106_),
    .B(net3424),
    .Y(_04138_));
 sky130_fd_sc_hd__a22o_1 _18281_ (.A1(_04126_),
    .A2(_09589_),
    .B1(_04118_),
    .B2(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__inv_2 _18282_ (.A(_04139_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _18283_ (.A(_09232_),
    .B(_04120_),
    .Y(_04140_));
 sky130_fd_sc_hd__a31o_1 _18284_ (.A1(_04129_),
    .A2(net2357),
    .A3(_04119_),
    .B1(_04140_),
    .X(_02188_));
 sky130_fd_sc_hd__nor2_1 _18285_ (.A(_09235_),
    .B(_04120_),
    .Y(_04141_));
 sky130_fd_sc_hd__a31o_1 _18286_ (.A1(_04129_),
    .A2(net1283),
    .A3(_04120_),
    .B1(_04141_),
    .X(_02189_));
 sky130_fd_sc_hd__nand2_1 _18287_ (.A(_04106_),
    .B(net3112),
    .Y(_04142_));
 sky130_fd_sc_hd__a22o_1 _18288_ (.A1(_04126_),
    .A2(_10202_),
    .B1(_04118_),
    .B2(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__inv_2 _18289_ (.A(_04143_),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _18290_ (.A(_04106_),
    .B(net3450),
    .Y(_04144_));
 sky130_fd_sc_hd__a22o_1 _18291_ (.A1(_04126_),
    .A2(_09767_),
    .B1(_04118_),
    .B2(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__inv_2 _18292_ (.A(_04145_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _18293_ (.A(_03294_),
    .B(_04120_),
    .Y(_04146_));
 sky130_fd_sc_hd__a31o_1 _18294_ (.A1(_04129_),
    .A2(net1808),
    .A3(_04120_),
    .B1(_04146_),
    .X(_02176_));
 sky130_fd_sc_hd__and3_1 _18295_ (.A(_04115_),
    .B(_03029_),
    .C(_04037_),
    .X(_04147_));
 sky130_fd_sc_hd__a31o_1 _18296_ (.A1(_04119_),
    .A2(_04044_),
    .A3(net2522),
    .B1(_04147_),
    .X(_02177_));
 sky130_fd_sc_hd__nor2_1 _18297_ (.A(_03482_),
    .B(_04120_),
    .Y(_04148_));
 sky130_fd_sc_hd__a31o_1 _18298_ (.A1(_04129_),
    .A2(net2329),
    .A3(_04120_),
    .B1(_04148_),
    .X(_02178_));
 sky130_fd_sc_hd__and3_1 _18299_ (.A(_04115_),
    .B(_03032_),
    .C(_04037_),
    .X(_04149_));
 sky130_fd_sc_hd__a31o_1 _18300_ (.A1(_04119_),
    .A2(_04044_),
    .A3(net2491),
    .B1(_04149_),
    .X(_02179_));
 sky130_fd_sc_hd__nand2_1 _18301_ (.A(_04106_),
    .B(net3466),
    .Y(_04150_));
 sky130_fd_sc_hd__a22o_1 _18302_ (.A1(_04126_),
    .A2(_11136_),
    .B1(_04118_),
    .B2(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__inv_2 _18303_ (.A(_04151_),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_1 _18304_ (.A(_04106_),
    .B(net3067),
    .Y(_04152_));
 sky130_fd_sc_hd__a22o_1 _18305_ (.A1(_04126_),
    .A2(_02916_),
    .B1(_04118_),
    .B2(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__inv_2 _18306_ (.A(_04153_),
    .Y(_02181_));
 sky130_fd_sc_hd__clkbuf_4 _18307_ (.A(_11219_),
    .X(_04154_));
 sky130_fd_sc_hd__and3_1 _18308_ (.A(_04115_),
    .B(net55),
    .C(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__a31o_1 _18309_ (.A1(_04119_),
    .A2(_04044_),
    .A3(net2201),
    .B1(_04155_),
    .X(_02182_));
 sky130_fd_sc_hd__nand2_1 _18310_ (.A(_04106_),
    .B(net3213),
    .Y(_04156_));
 sky130_fd_sc_hd__a22o_1 _18311_ (.A1(_04126_),
    .A2(_02921_),
    .B1(_04118_),
    .B2(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__inv_2 _18312_ (.A(_04157_),
    .Y(_02183_));
 sky130_fd_sc_hd__and3_1 _18313_ (.A(_04115_),
    .B(_03196_),
    .C(_04154_),
    .X(_04158_));
 sky130_fd_sc_hd__a31o_1 _18314_ (.A1(_04119_),
    .A2(_04044_),
    .A3(net2402),
    .B1(_04158_),
    .X(_02168_));
 sky130_fd_sc_hd__nor2_1 _18315_ (.A(_03605_),
    .B(_04120_),
    .Y(_04159_));
 sky130_fd_sc_hd__a31o_1 _18316_ (.A1(_04129_),
    .A2(net1041),
    .A3(_04120_),
    .B1(_04159_),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_1 _18317_ (.A(_04106_),
    .B(net3269),
    .Y(_04160_));
 sky130_fd_sc_hd__a22o_1 _18318_ (.A1(_04126_),
    .A2(_10624_),
    .B1(_04118_),
    .B2(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__inv_2 _18319_ (.A(_04161_),
    .Y(_02170_));
 sky130_fd_sc_hd__nand2_1 _18320_ (.A(_04106_),
    .B(net3456),
    .Y(_04162_));
 sky130_fd_sc_hd__a22o_1 _18321_ (.A1(_04126_),
    .A2(_02928_),
    .B1(_04118_),
    .B2(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__inv_2 _18322_ (.A(_04163_),
    .Y(_02171_));
 sky130_fd_sc_hd__buf_4 _18323_ (.A(_03834_),
    .X(_04164_));
 sky130_fd_sc_hd__and3_1 _18324_ (.A(_04115_),
    .B(_03550_),
    .C(_04154_),
    .X(_04165_));
 sky130_fd_sc_hd__a31o_1 _18325_ (.A1(_04119_),
    .A2(_04164_),
    .A3(net2386),
    .B1(_04165_),
    .X(_02172_));
 sky130_fd_sc_hd__nand2_1 _18326_ (.A(_03317_),
    .B(net3847),
    .Y(_04166_));
 sky130_fd_sc_hd__o2bb2a_1 _18327_ (.A1_N(_04166_),
    .A2_N(_04119_),
    .B1(_09294_),
    .B2(_04116_),
    .X(_02173_));
 sky130_fd_sc_hd__nand2_1 _18328_ (.A(_03317_),
    .B(net3705),
    .Y(_04167_));
 sky130_fd_sc_hd__o2bb2a_1 _18329_ (.A1_N(_04167_),
    .A2_N(_04119_),
    .B1(_02992_),
    .B2(_04116_),
    .X(_02174_));
 sky130_fd_sc_hd__nand2_1 _18330_ (.A(_03317_),
    .B(net3732),
    .Y(_04168_));
 sky130_fd_sc_hd__o2bb2a_1 _18331_ (.A1_N(_04168_),
    .A2_N(_04119_),
    .B1(_11316_),
    .B2(_04116_),
    .X(_02175_));
 sky130_fd_sc_hd__and3_4 _18332_ (.A(_09171_),
    .B(_09444_),
    .C(_09380_),
    .X(_04169_));
 sky130_fd_sc_hd__inv_2 _18333_ (.A(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__nor2_1 _18334_ (.A(_09625_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__inv_2 _18335_ (.A(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__buf_4 _18336_ (.A(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__buf_4 _18337_ (.A(_04172_),
    .X(_04174_));
 sky130_fd_sc_hd__nor2_1 _18338_ (.A(_09180_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__a31o_1 _18339_ (.A1(_04129_),
    .A2(net1541),
    .A3(_04173_),
    .B1(_04175_),
    .X(_02160_));
 sky130_fd_sc_hd__nor2_1 _18340_ (.A(_03170_),
    .B(_04174_),
    .Y(_04176_));
 sky130_fd_sc_hd__a31o_1 _18341_ (.A1(_04129_),
    .A2(net1643),
    .A3(_04173_),
    .B1(_04176_),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_4 _18342_ (.A(_08797_),
    .B(_04170_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_1 _18343_ (.A(_04106_),
    .B(net3177),
    .Y(_04178_));
 sky130_fd_sc_hd__a22o_1 _18344_ (.A1(_04177_),
    .A2(_09459_),
    .B1(_04174_),
    .B2(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__inv_2 _18345_ (.A(_04179_),
    .Y(_02162_));
 sky130_fd_sc_hd__and3_1 _18346_ (.A(_04169_),
    .B(net69),
    .C(_04154_),
    .X(_04180_));
 sky130_fd_sc_hd__a31o_1 _18347_ (.A1(_04173_),
    .A2(_04164_),
    .A3(net2178),
    .B1(_04180_),
    .X(_02163_));
 sky130_fd_sc_hd__nand2_1 _18348_ (.A(_04106_),
    .B(net3561),
    .Y(_04181_));
 sky130_fd_sc_hd__a22o_1 _18349_ (.A1(_04177_),
    .A2(_11330_),
    .B1(_04174_),
    .B2(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__inv_2 _18350_ (.A(_04182_),
    .Y(_02164_));
 sky130_fd_sc_hd__and3_1 _18351_ (.A(_04169_),
    .B(_11391_),
    .C(_04154_),
    .X(_04183_));
 sky130_fd_sc_hd__a31o_1 _18352_ (.A1(_04173_),
    .A2(_04164_),
    .A3(net1733),
    .B1(_04183_),
    .X(_02165_));
 sky130_fd_sc_hd__buf_4 _18353_ (.A(_08775_),
    .X(_04184_));
 sky130_fd_sc_hd__buf_4 _18354_ (.A(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__nand2_1 _18355_ (.A(_04185_),
    .B(net3386),
    .Y(_04186_));
 sky130_fd_sc_hd__a22o_1 _18356_ (.A1(_04177_),
    .A2(_11105_),
    .B1(_04174_),
    .B2(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__inv_2 _18357_ (.A(_04187_),
    .Y(_02166_));
 sky130_fd_sc_hd__and3_1 _18358_ (.A(_04169_),
    .B(net74),
    .C(_04154_),
    .X(_04188_));
 sky130_fd_sc_hd__a31o_1 _18359_ (.A1(_04173_),
    .A2(_04164_),
    .A3(net1562),
    .B1(_04188_),
    .X(_02167_));
 sky130_fd_sc_hd__nand2_1 _18360_ (.A(_04185_),
    .B(net3322),
    .Y(_04189_));
 sky130_fd_sc_hd__a22o_1 _18361_ (.A1(_04177_),
    .A2(net135),
    .B1(_04174_),
    .B2(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__inv_2 _18362_ (.A(_04190_),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_1 _18363_ (.A(_04185_),
    .B(net3680),
    .Y(_04191_));
 sky130_fd_sc_hd__a22o_1 _18364_ (.A1(_04177_),
    .A2(_02899_),
    .B1(_04174_),
    .B2(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__inv_2 _18365_ (.A(_04192_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_1 _18366_ (.A(_04185_),
    .B(net3377),
    .Y(_04193_));
 sky130_fd_sc_hd__a22o_1 _18367_ (.A1(_04177_),
    .A2(_02963_),
    .B1(_04174_),
    .B2(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__inv_2 _18368_ (.A(_04194_),
    .Y(_02154_));
 sky130_fd_sc_hd__nand2_1 _18369_ (.A(_04185_),
    .B(net3285),
    .Y(_04195_));
 sky130_fd_sc_hd__a22o_1 _18370_ (.A1(_04177_),
    .A2(_09588_),
    .B1(_04172_),
    .B2(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__inv_2 _18371_ (.A(_04196_),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _18372_ (.A(_09232_),
    .B(_04174_),
    .Y(_04197_));
 sky130_fd_sc_hd__a31o_1 _18373_ (.A1(_04129_),
    .A2(net2037),
    .A3(_04173_),
    .B1(_04197_),
    .X(_02156_));
 sky130_fd_sc_hd__nor2_1 _18374_ (.A(_09235_),
    .B(_04174_),
    .Y(_04198_));
 sky130_fd_sc_hd__a31o_1 _18375_ (.A1(_04129_),
    .A2(net1201),
    .A3(_04173_),
    .B1(_04198_),
    .X(_02157_));
 sky130_fd_sc_hd__and3_1 _18376_ (.A(_04169_),
    .B(net64),
    .C(_04154_),
    .X(_04199_));
 sky130_fd_sc_hd__a31o_1 _18377_ (.A1(_04173_),
    .A2(_04164_),
    .A3(net1761),
    .B1(_04199_),
    .X(_02158_));
 sky130_fd_sc_hd__nor2_1 _18378_ (.A(_03026_),
    .B(_04174_),
    .Y(_04200_));
 sky130_fd_sc_hd__a31o_1 _18379_ (.A1(_04129_),
    .A2(net661),
    .A3(_04173_),
    .B1(_04200_),
    .X(_02159_));
 sky130_fd_sc_hd__nor2_1 _18380_ (.A(_03294_),
    .B(_04174_),
    .Y(_04201_));
 sky130_fd_sc_hd__a31o_1 _18381_ (.A1(_04129_),
    .A2(net1985),
    .A3(_04173_),
    .B1(_04201_),
    .X(_02144_));
 sky130_fd_sc_hd__and3_1 _18382_ (.A(_04169_),
    .B(net82),
    .C(_04154_),
    .X(_04202_));
 sky130_fd_sc_hd__a31o_1 _18383_ (.A1(_04173_),
    .A2(_04164_),
    .A3(net2019),
    .B1(_04202_),
    .X(_02145_));
 sky130_fd_sc_hd__nor2_1 _18384_ (.A(_03482_),
    .B(_04174_),
    .Y(_04203_));
 sky130_fd_sc_hd__a31o_1 _18385_ (.A1(_04129_),
    .A2(net2036),
    .A3(_04174_),
    .B1(_04203_),
    .X(_02146_));
 sky130_fd_sc_hd__and3_1 _18386_ (.A(_04169_),
    .B(net52),
    .C(_04154_),
    .X(_04204_));
 sky130_fd_sc_hd__a31o_1 _18387_ (.A1(_04173_),
    .A2(_04164_),
    .A3(net1845),
    .B1(_04204_),
    .X(_02147_));
 sky130_fd_sc_hd__nor2_1 _18388_ (.A(_09259_),
    .B(_04174_),
    .Y(_04205_));
 sky130_fd_sc_hd__a31o_1 _18389_ (.A1(_04129_),
    .A2(net2431),
    .A3(_04174_),
    .B1(_04205_),
    .X(_02148_));
 sky130_fd_sc_hd__nand2_1 _18390_ (.A(_04185_),
    .B(net3759),
    .Y(_04206_));
 sky130_fd_sc_hd__a22o_1 _18391_ (.A1(_04177_),
    .A2(_02916_),
    .B1(_04172_),
    .B2(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__inv_2 _18392_ (.A(_04207_),
    .Y(_02149_));
 sky130_fd_sc_hd__and3_1 _18393_ (.A(_04169_),
    .B(net55),
    .C(_04154_),
    .X(_04208_));
 sky130_fd_sc_hd__a31o_1 _18394_ (.A1(_04173_),
    .A2(_04164_),
    .A3(net2243),
    .B1(_04208_),
    .X(_02150_));
 sky130_fd_sc_hd__nand2_1 _18395_ (.A(_04185_),
    .B(net3114),
    .Y(_04209_));
 sky130_fd_sc_hd__a22o_1 _18396_ (.A1(_04177_),
    .A2(_02921_),
    .B1(_04172_),
    .B2(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__inv_2 _18397_ (.A(_04210_),
    .Y(_02151_));
 sky130_fd_sc_hd__nand2_1 _18398_ (.A(_04185_),
    .B(net3420),
    .Y(_04211_));
 sky130_fd_sc_hd__a22o_1 _18399_ (.A1(_04177_),
    .A2(net141),
    .B1(_04172_),
    .B2(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__inv_2 _18400_ (.A(_04212_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _18401_ (.A(_04185_),
    .B(net3229),
    .Y(_04213_));
 sky130_fd_sc_hd__a22o_1 _18402_ (.A1(_04177_),
    .A2(_09365_),
    .B1(_04172_),
    .B2(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__inv_2 _18403_ (.A(_04214_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_1 _18404_ (.A(_04185_),
    .B(net3630),
    .Y(_04215_));
 sky130_fd_sc_hd__a22o_1 _18405_ (.A1(_04177_),
    .A2(_10624_),
    .B1(_04172_),
    .B2(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__inv_2 _18406_ (.A(_04216_),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2_1 _18407_ (.A(_04185_),
    .B(net3087),
    .Y(_04217_));
 sky130_fd_sc_hd__a22o_1 _18408_ (.A1(_04177_),
    .A2(_02928_),
    .B1(_04172_),
    .B2(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__inv_2 _18409_ (.A(_04218_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand2_1 _18410_ (.A(_04185_),
    .B(net3263),
    .Y(_04219_));
 sky130_fd_sc_hd__a22o_1 _18411_ (.A1(_04177_),
    .A2(_09287_),
    .B1(_04172_),
    .B2(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__inv_2 _18412_ (.A(_04220_),
    .Y(_02140_));
 sky130_fd_sc_hd__clkbuf_8 _18413_ (.A(_08800_),
    .X(_04221_));
 sky130_fd_sc_hd__nand2_1 _18414_ (.A(_04221_),
    .B(net3566),
    .Y(_04222_));
 sky130_fd_sc_hd__o2bb2a_1 _18415_ (.A1_N(_04222_),
    .A2_N(_04173_),
    .B1(_09294_),
    .B2(_04170_),
    .X(_02141_));
 sky130_fd_sc_hd__nand2_1 _18416_ (.A(_04221_),
    .B(net3738),
    .Y(_04223_));
 sky130_fd_sc_hd__o2bb2a_1 _18417_ (.A1_N(_04223_),
    .A2_N(_04173_),
    .B1(_02992_),
    .B2(_04170_),
    .X(_02142_));
 sky130_fd_sc_hd__nand2_1 _18418_ (.A(_04221_),
    .B(net3451),
    .Y(_04224_));
 sky130_fd_sc_hd__o2bb2a_1 _18419_ (.A1_N(_04224_),
    .A2_N(_04173_),
    .B1(_11316_),
    .B2(_04170_),
    .X(_02143_));
 sky130_fd_sc_hd__nor2_4 _18420_ (.A(_08736_),
    .B(_09446_),
    .Y(_04225_));
 sky130_fd_sc_hd__inv_2 _18421_ (.A(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__nor2_1 _18422_ (.A(_09304_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__clkinv_4 _18423_ (.A(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__buf_4 _18424_ (.A(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__buf_4 _18425_ (.A(_04228_),
    .X(_04230_));
 sky130_fd_sc_hd__nor2_1 _18426_ (.A(_09180_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__a31o_1 _18427_ (.A1(_04129_),
    .A2(net1249),
    .A3(_04229_),
    .B1(_04231_),
    .X(_02128_));
 sky130_fd_sc_hd__nor2_4 _18428_ (.A(_09190_),
    .B(_04226_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_1 _18429_ (.A(_04185_),
    .B(net3009),
    .Y(_04233_));
 sky130_fd_sc_hd__a22o_1 _18430_ (.A1(_04232_),
    .A2(_09314_),
    .B1(_04230_),
    .B2(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__inv_2 _18431_ (.A(_04234_),
    .Y(_02129_));
 sky130_fd_sc_hd__clkbuf_8 _18432_ (.A(_09164_),
    .X(_04235_));
 sky130_fd_sc_hd__nor2_1 _18433_ (.A(_03219_),
    .B(_04230_),
    .Y(_04236_));
 sky130_fd_sc_hd__a31o_1 _18434_ (.A1(_04235_),
    .A2(net1045),
    .A3(_04229_),
    .B1(_04236_),
    .X(_02130_));
 sky130_fd_sc_hd__nand2_1 _18435_ (.A(_04185_),
    .B(net3457),
    .Y(_04237_));
 sky130_fd_sc_hd__a22o_1 _18436_ (.A1(_04232_),
    .A2(_10983_),
    .B1(_04230_),
    .B2(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__inv_2 _18437_ (.A(_04238_),
    .Y(_02131_));
 sky130_fd_sc_hd__and3_1 _18438_ (.A(_04225_),
    .B(_10586_),
    .C(_04154_),
    .X(_04239_));
 sky130_fd_sc_hd__a31o_1 _18439_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net2559),
    .B1(_04239_),
    .X(_02132_));
 sky130_fd_sc_hd__and3_1 _18440_ (.A(_04225_),
    .B(net71),
    .C(_04154_),
    .X(_04240_));
 sky130_fd_sc_hd__a31o_1 _18441_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net2083),
    .B1(_04240_),
    .X(_02133_));
 sky130_fd_sc_hd__nor2_1 _18442_ (.A(_09208_),
    .B(_04230_),
    .Y(_04241_));
 sky130_fd_sc_hd__a31o_1 _18443_ (.A1(_04235_),
    .A2(net2404),
    .A3(_04229_),
    .B1(_04241_),
    .X(_02134_));
 sky130_fd_sc_hd__nand2_1 _18444_ (.A(_04185_),
    .B(net3249),
    .Y(_04242_));
 sky130_fd_sc_hd__a22o_1 _18445_ (.A1(_04232_),
    .A2(_10591_),
    .B1(_04228_),
    .B2(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__inv_2 _18446_ (.A(_04243_),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _18447_ (.A(_04185_),
    .B(net3410),
    .Y(_04244_));
 sky130_fd_sc_hd__a22o_1 _18448_ (.A1(_04232_),
    .A2(net135),
    .B1(_04228_),
    .B2(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__inv_2 _18449_ (.A(_04245_),
    .Y(_02120_));
 sky130_fd_sc_hd__buf_4 _18450_ (.A(_04184_),
    .X(_04246_));
 sky130_fd_sc_hd__nand2_1 _18451_ (.A(_04246_),
    .B(net3555),
    .Y(_04247_));
 sky130_fd_sc_hd__a22o_1 _18452_ (.A1(_04232_),
    .A2(_02899_),
    .B1(_04228_),
    .B2(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__inv_2 _18453_ (.A(_04248_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _18454_ (.A(_04246_),
    .B(net3402),
    .Y(_04249_));
 sky130_fd_sc_hd__a22o_1 _18455_ (.A1(_04232_),
    .A2(_02963_),
    .B1(_04228_),
    .B2(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__inv_2 _18456_ (.A(_04250_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _18457_ (.A(_09229_),
    .B(_04230_),
    .Y(_04251_));
 sky130_fd_sc_hd__a31o_1 _18458_ (.A1(_04235_),
    .A2(net1321),
    .A3(_04229_),
    .B1(_04251_),
    .X(_02123_));
 sky130_fd_sc_hd__nor2_1 _18459_ (.A(_09232_),
    .B(_04230_),
    .Y(_04252_));
 sky130_fd_sc_hd__a31o_1 _18460_ (.A1(_04235_),
    .A2(net1177),
    .A3(_04229_),
    .B1(_04252_),
    .X(_02124_));
 sky130_fd_sc_hd__nor2_1 _18461_ (.A(_09235_),
    .B(_04230_),
    .Y(_04253_));
 sky130_fd_sc_hd__a31o_1 _18462_ (.A1(_04235_),
    .A2(net1383),
    .A3(_04229_),
    .B1(_04253_),
    .X(_02125_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(_04246_),
    .B(net3054),
    .Y(_04254_));
 sky130_fd_sc_hd__a22o_1 _18464_ (.A1(_04232_),
    .A2(_10202_),
    .B1(_04228_),
    .B2(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__inv_2 _18465_ (.A(_04255_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor2_1 _18466_ (.A(_03026_),
    .B(_04230_),
    .Y(_04256_));
 sky130_fd_sc_hd__a31o_1 _18467_ (.A1(_04235_),
    .A2(net1263),
    .A3(_04230_),
    .B1(_04256_),
    .X(_02127_));
 sky130_fd_sc_hd__nand2_1 _18468_ (.A(_04246_),
    .B(net3504),
    .Y(_04257_));
 sky130_fd_sc_hd__a22o_1 _18469_ (.A1(_04232_),
    .A2(net138),
    .B1(_04228_),
    .B2(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__inv_2 _18470_ (.A(_04258_),
    .Y(_02104_));
 sky130_fd_sc_hd__and3_1 _18471_ (.A(_04225_),
    .B(net82),
    .C(_04154_),
    .X(_04259_));
 sky130_fd_sc_hd__a31o_1 _18472_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net2270),
    .B1(_04259_),
    .X(_02105_));
 sky130_fd_sc_hd__nor2_1 _18473_ (.A(_03482_),
    .B(_04230_),
    .Y(_04260_));
 sky130_fd_sc_hd__a31o_1 _18474_ (.A1(_04235_),
    .A2(net2562),
    .A3(_04230_),
    .B1(_04260_),
    .X(_02106_));
 sky130_fd_sc_hd__and3_1 _18475_ (.A(_04225_),
    .B(net52),
    .C(_04154_),
    .X(_04261_));
 sky130_fd_sc_hd__a31o_1 _18476_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net1917),
    .B1(_04261_),
    .X(_02107_));
 sky130_fd_sc_hd__nor2_1 _18477_ (.A(_09259_),
    .B(_04230_),
    .Y(_04262_));
 sky130_fd_sc_hd__a31o_1 _18478_ (.A1(_04235_),
    .A2(net1015),
    .A3(_04230_),
    .B1(_04262_),
    .X(_02108_));
 sky130_fd_sc_hd__nand2_1 _18479_ (.A(_04246_),
    .B(net3104),
    .Y(_04263_));
 sky130_fd_sc_hd__a22o_1 _18480_ (.A1(_04232_),
    .A2(_02916_),
    .B1(_04228_),
    .B2(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__inv_2 _18481_ (.A(_04264_),
    .Y(_02109_));
 sky130_fd_sc_hd__and3_1 _18482_ (.A(_04225_),
    .B(net55),
    .C(_04154_),
    .X(_04265_));
 sky130_fd_sc_hd__a31o_1 _18483_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net2304),
    .B1(_04265_),
    .X(_02110_));
 sky130_fd_sc_hd__nand2_1 _18484_ (.A(_04246_),
    .B(net2979),
    .Y(_04266_));
 sky130_fd_sc_hd__a22o_1 _18485_ (.A1(_04232_),
    .A2(_02921_),
    .B1(_04228_),
    .B2(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__inv_2 _18486_ (.A(_04267_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_04246_),
    .B(net3240),
    .Y(_04268_));
 sky130_fd_sc_hd__a22o_1 _18488_ (.A1(_04232_),
    .A2(net141),
    .B1(_04228_),
    .B2(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__inv_2 _18489_ (.A(_04269_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_1 _18490_ (.A(_03605_),
    .B(_04230_),
    .Y(_04270_));
 sky130_fd_sc_hd__a31o_1 _18491_ (.A1(_04235_),
    .A2(net2359),
    .A3(_04230_),
    .B1(_04270_),
    .X(_02097_));
 sky130_fd_sc_hd__and3_1 _18492_ (.A(_04225_),
    .B(_03199_),
    .C(_04154_),
    .X(_04271_));
 sky130_fd_sc_hd__a31o_1 _18493_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net2215),
    .B1(_04271_),
    .X(_02098_));
 sky130_fd_sc_hd__nand2_1 _18494_ (.A(_04246_),
    .B(net3098),
    .Y(_04272_));
 sky130_fd_sc_hd__a22o_1 _18495_ (.A1(_04232_),
    .A2(_02928_),
    .B1(_04228_),
    .B2(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__inv_2 _18496_ (.A(_04273_),
    .Y(_02099_));
 sky130_fd_sc_hd__buf_4 _18497_ (.A(_09226_),
    .X(_04274_));
 sky130_fd_sc_hd__and3_1 _18498_ (.A(_04225_),
    .B(_03550_),
    .C(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__a31o_1 _18499_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net2238),
    .B1(_04275_),
    .X(_02100_));
 sky130_fd_sc_hd__and3_1 _18500_ (.A(_04225_),
    .B(net78),
    .C(_04274_),
    .X(_04276_));
 sky130_fd_sc_hd__a31o_1 _18501_ (.A1(_04229_),
    .A2(_04164_),
    .A3(net1964),
    .B1(_04276_),
    .X(_02101_));
 sky130_fd_sc_hd__nand2_1 _18502_ (.A(_04221_),
    .B(net3765),
    .Y(_04277_));
 sky130_fd_sc_hd__o2bb2a_1 _18503_ (.A1_N(_04277_),
    .A2_N(_04229_),
    .B1(_02992_),
    .B2(_04226_),
    .X(_02102_));
 sky130_fd_sc_hd__nand2_1 _18504_ (.A(_04221_),
    .B(net3748),
    .Y(_04278_));
 sky130_fd_sc_hd__o2bb2a_1 _18505_ (.A1_N(_04278_),
    .A2_N(_04229_),
    .B1(_11316_),
    .B2(_04226_),
    .X(_02103_));
 sky130_fd_sc_hd__nor2_1 _18506_ (.A(_08736_),
    .B(_09512_),
    .Y(_04279_));
 sky130_fd_sc_hd__inv_2 _18507_ (.A(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__nor2_4 _18508_ (.A(_08794_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__buf_4 _18509_ (.A(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__nor2_1 _18510_ (.A(_09166_),
    .B(_04280_),
    .Y(_04283_));
 sky130_fd_sc_hd__inv_2 _18511_ (.A(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__buf_4 _18512_ (.A(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__nand2_1 _18513_ (.A(_04246_),
    .B(net3065),
    .Y(_04286_));
 sky130_fd_sc_hd__a22o_1 _18514_ (.A1(_04282_),
    .A2(_10239_),
    .B1(_04285_),
    .B2(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__inv_2 _18515_ (.A(_04287_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2_1 _18516_ (.A(_04246_),
    .B(net3101),
    .Y(_04288_));
 sky130_fd_sc_hd__a22o_1 _18517_ (.A1(_04282_),
    .A2(_09314_),
    .B1(_04285_),
    .B2(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__inv_2 _18518_ (.A(_04289_),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_1 _18519_ (.A(_04246_),
    .B(net3295),
    .Y(_04290_));
 sky130_fd_sc_hd__a22o_1 _18520_ (.A1(_04282_),
    .A2(_09459_),
    .B1(_04285_),
    .B2(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__inv_2 _18521_ (.A(_04291_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(_04246_),
    .B(net3256),
    .Y(_04292_));
 sky130_fd_sc_hd__a22o_1 _18523_ (.A1(_04282_),
    .A2(_10983_),
    .B1(_04285_),
    .B2(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__inv_2 _18524_ (.A(_04293_),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2_1 _18525_ (.A(_04246_),
    .B(net2882),
    .Y(_04294_));
 sky130_fd_sc_hd__a22o_1 _18526_ (.A1(_04282_),
    .A2(_11330_),
    .B1(_04285_),
    .B2(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__inv_2 _18527_ (.A(_04295_),
    .Y(_02092_));
 sky130_fd_sc_hd__nand2_1 _18528_ (.A(_04246_),
    .B(net3028),
    .Y(_04296_));
 sky130_fd_sc_hd__a22o_1 _18529_ (.A1(_04282_),
    .A2(_09204_),
    .B1(_04285_),
    .B2(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__inv_2 _18530_ (.A(_04297_),
    .Y(_02093_));
 sky130_fd_sc_hd__nand2_1 _18531_ (.A(_04246_),
    .B(net3521),
    .Y(_04298_));
 sky130_fd_sc_hd__a22o_1 _18532_ (.A1(_04282_),
    .A2(_11105_),
    .B1(_04285_),
    .B2(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__inv_2 _18533_ (.A(_04299_),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_1 _18534_ (.A(_04246_),
    .B(net3380),
    .Y(_04300_));
 sky130_fd_sc_hd__a22o_1 _18535_ (.A1(_04282_),
    .A2(_09211_),
    .B1(_04285_),
    .B2(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__inv_2 _18536_ (.A(_04301_),
    .Y(_02095_));
 sky130_fd_sc_hd__buf_4 _18537_ (.A(_04184_),
    .X(_04302_));
 sky130_fd_sc_hd__nand2_1 _18538_ (.A(_04302_),
    .B(net2993),
    .Y(_04303_));
 sky130_fd_sc_hd__a22o_1 _18539_ (.A1(_04282_),
    .A2(_09530_),
    .B1(_04285_),
    .B2(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__inv_2 _18540_ (.A(_04304_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _18541_ (.A(_04302_),
    .B(net3150),
    .Y(_04305_));
 sky130_fd_sc_hd__a22o_1 _18542_ (.A1(_04282_),
    .A2(_02899_),
    .B1(_04285_),
    .B2(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__inv_2 _18543_ (.A(_04306_),
    .Y(_02081_));
 sky130_fd_sc_hd__nand2_1 _18544_ (.A(_04302_),
    .B(net2965),
    .Y(_04307_));
 sky130_fd_sc_hd__a22o_1 _18545_ (.A1(_04282_),
    .A2(_02963_),
    .B1(_04285_),
    .B2(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__inv_2 _18546_ (.A(_04308_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _18547_ (.A(_04302_),
    .B(net2861),
    .Y(_04309_));
 sky130_fd_sc_hd__a22o_1 _18548_ (.A1(_04282_),
    .A2(_09588_),
    .B1(_04285_),
    .B2(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__inv_2 _18549_ (.A(_04310_),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _18550_ (.A(_04302_),
    .B(net3004),
    .Y(_04311_));
 sky130_fd_sc_hd__a22o_1 _18551_ (.A1(_04282_),
    .A2(_09592_),
    .B1(_04285_),
    .B2(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__inv_2 _18552_ (.A(_04312_),
    .Y(_02084_));
 sky130_fd_sc_hd__buf_4 _18553_ (.A(_04284_),
    .X(_04313_));
 sky130_fd_sc_hd__nand2_1 _18554_ (.A(_04302_),
    .B(net3071),
    .Y(_04314_));
 sky130_fd_sc_hd__a22o_1 _18555_ (.A1(_04282_),
    .A2(_09338_),
    .B1(_04313_),
    .B2(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__inv_2 _18556_ (.A(_04315_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_1 _18557_ (.A(_04302_),
    .B(net3183),
    .Y(_04316_));
 sky130_fd_sc_hd__a22o_1 _18558_ (.A1(_04282_),
    .A2(_10202_),
    .B1(_04313_),
    .B2(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__inv_2 _18559_ (.A(_04317_),
    .Y(_02086_));
 sky130_fd_sc_hd__nand2_1 _18560_ (.A(_04302_),
    .B(net3175),
    .Y(_04318_));
 sky130_fd_sc_hd__a22o_1 _18561_ (.A1(_04282_),
    .A2(_09767_),
    .B1(_04313_),
    .B2(_04318_),
    .X(_04319_));
 sky130_fd_sc_hd__inv_2 _18562_ (.A(_04319_),
    .Y(_02087_));
 sky130_fd_sc_hd__nand2_1 _18563_ (.A(_04302_),
    .B(net3284),
    .Y(_04320_));
 sky130_fd_sc_hd__a22o_1 _18564_ (.A1(_04281_),
    .A2(net137),
    .B1(_04313_),
    .B2(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__inv_2 _18565_ (.A(_04321_),
    .Y(_02072_));
 sky130_fd_sc_hd__nand2_1 _18566_ (.A(_04302_),
    .B(net3090),
    .Y(_04322_));
 sky130_fd_sc_hd__a22o_1 _18567_ (.A1(_04281_),
    .A2(_09248_),
    .B1(_04313_),
    .B2(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__inv_2 _18568_ (.A(_04323_),
    .Y(_02073_));
 sky130_fd_sc_hd__nand2_1 _18569_ (.A(_04302_),
    .B(net3144),
    .Y(_04324_));
 sky130_fd_sc_hd__a22o_1 _18570_ (.A1(_04281_),
    .A2(_09347_),
    .B1(_04313_),
    .B2(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__inv_2 _18571_ (.A(_04325_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2_1 _18572_ (.A(_04302_),
    .B(net3438),
    .Y(_04326_));
 sky130_fd_sc_hd__a22o_1 _18573_ (.A1(_04281_),
    .A2(_09255_),
    .B1(_04313_),
    .B2(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__inv_2 _18574_ (.A(_04327_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_1 _18575_ (.A(_04302_),
    .B(net3205),
    .Y(_04328_));
 sky130_fd_sc_hd__a22o_1 _18576_ (.A1(_04281_),
    .A2(_11136_),
    .B1(_04313_),
    .B2(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__inv_2 _18577_ (.A(_04329_),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_1 _18578_ (.A(_04302_),
    .B(net3473),
    .Y(_04330_));
 sky130_fd_sc_hd__a22o_1 _18579_ (.A1(_04281_),
    .A2(_02916_),
    .B1(_04313_),
    .B2(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__inv_2 _18580_ (.A(_04331_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_1 _18581_ (.A(_04302_),
    .B(net3220),
    .Y(_04332_));
 sky130_fd_sc_hd__a22o_1 _18582_ (.A1(_04281_),
    .A2(_09424_),
    .B1(_04313_),
    .B2(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__inv_2 _18583_ (.A(_04333_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand2_1 _18584_ (.A(_04302_),
    .B(net2997),
    .Y(_04334_));
 sky130_fd_sc_hd__a22o_1 _18585_ (.A1(_04281_),
    .A2(_02921_),
    .B1(_04313_),
    .B2(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__inv_2 _18586_ (.A(_04335_),
    .Y(_02079_));
 sky130_fd_sc_hd__buf_4 _18587_ (.A(_04184_),
    .X(_04336_));
 sky130_fd_sc_hd__nand2_1 _18588_ (.A(_04336_),
    .B(net2804),
    .Y(_04337_));
 sky130_fd_sc_hd__a22o_1 _18589_ (.A1(_04281_),
    .A2(_09494_),
    .B1(_04313_),
    .B2(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__inv_2 _18590_ (.A(_04338_),
    .Y(_02064_));
 sky130_fd_sc_hd__nand2_1 _18591_ (.A(_04336_),
    .B(net3222),
    .Y(_04339_));
 sky130_fd_sc_hd__a22o_1 _18592_ (.A1(_04281_),
    .A2(_09365_),
    .B1(_04313_),
    .B2(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__inv_2 _18593_ (.A(_04340_),
    .Y(_02065_));
 sky130_fd_sc_hd__nand2_1 _18594_ (.A(_04336_),
    .B(net3202),
    .Y(_04341_));
 sky130_fd_sc_hd__a22o_1 _18595_ (.A1(_04281_),
    .A2(_10624_),
    .B1(_04313_),
    .B2(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__inv_2 _18596_ (.A(_04342_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _18597_ (.A(_04336_),
    .B(net3010),
    .Y(_04343_));
 sky130_fd_sc_hd__a22o_1 _18598_ (.A1(_04281_),
    .A2(_02928_),
    .B1(_04313_),
    .B2(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__inv_2 _18599_ (.A(_04344_),
    .Y(_02067_));
 sky130_fd_sc_hd__nand2_1 _18600_ (.A(_04336_),
    .B(net3370),
    .Y(_04345_));
 sky130_fd_sc_hd__a22o_1 _18601_ (.A1(_04281_),
    .A2(_09287_),
    .B1(_04313_),
    .B2(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__inv_2 _18602_ (.A(_04346_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _18603_ (.A(_04221_),
    .B(net3512),
    .Y(_04347_));
 sky130_fd_sc_hd__o2bb2a_1 _18604_ (.A1_N(_04347_),
    .A2_N(_04285_),
    .B1(_09294_),
    .B2(_04280_),
    .X(_02069_));
 sky130_fd_sc_hd__nand2_1 _18605_ (.A(_04221_),
    .B(net3662),
    .Y(_04348_));
 sky130_fd_sc_hd__o2bb2a_1 _18606_ (.A1_N(_04348_),
    .A2_N(_04285_),
    .B1(_02992_),
    .B2(_04280_),
    .X(_02070_));
 sky130_fd_sc_hd__nand2_1 _18607_ (.A(_04221_),
    .B(net3449),
    .Y(_04349_));
 sky130_fd_sc_hd__o2bb2a_1 _18608_ (.A1_N(_04349_),
    .A2_N(_04285_),
    .B1(_11316_),
    .B2(_04280_),
    .X(_02071_));
 sky130_fd_sc_hd__and3_4 _18609_ (.A(_09511_),
    .B(_09444_),
    .C(_09305_),
    .X(_04350_));
 sky130_fd_sc_hd__inv_2 _18610_ (.A(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__nor2_1 _18611_ (.A(_08728_),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__inv_2 _18612_ (.A(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__buf_4 _18613_ (.A(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__nor2_1 _18614_ (.A(_09180_),
    .B(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__a31o_1 _18615_ (.A1(_04235_),
    .A2(net1367),
    .A3(_04354_),
    .B1(_04355_),
    .X(_02056_));
 sky130_fd_sc_hd__nor2_1 _18616_ (.A(_08797_),
    .B(_04351_),
    .Y(_04356_));
 sky130_fd_sc_hd__buf_4 _18617_ (.A(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__buf_4 _18618_ (.A(_04353_),
    .X(_04358_));
 sky130_fd_sc_hd__nand2_1 _18619_ (.A(_04336_),
    .B(net2955),
    .Y(_04359_));
 sky130_fd_sc_hd__a22o_1 _18620_ (.A1(_04357_),
    .A2(_09314_),
    .B1(_04358_),
    .B2(_04359_),
    .X(_04360_));
 sky130_fd_sc_hd__inv_2 _18621_ (.A(_04360_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_1 _18622_ (.A(_04336_),
    .B(net3153),
    .Y(_04361_));
 sky130_fd_sc_hd__a22o_1 _18623_ (.A1(_04357_),
    .A2(_09459_),
    .B1(_04358_),
    .B2(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__inv_2 _18624_ (.A(_04362_),
    .Y(_02058_));
 sky130_fd_sc_hd__nand2_1 _18625_ (.A(_04336_),
    .B(net3698),
    .Y(_04363_));
 sky130_fd_sc_hd__a22o_1 _18626_ (.A1(_04357_),
    .A2(_10983_),
    .B1(_04358_),
    .B2(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__inv_2 _18627_ (.A(_04364_),
    .Y(_02059_));
 sky130_fd_sc_hd__buf_4 _18628_ (.A(_03834_),
    .X(_04365_));
 sky130_fd_sc_hd__and3_1 _18629_ (.A(_04350_),
    .B(_10586_),
    .C(_04274_),
    .X(_04366_));
 sky130_fd_sc_hd__a31o_1 _18630_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net2432),
    .B1(_04366_),
    .X(_02060_));
 sky130_fd_sc_hd__and3_1 _18631_ (.A(_04350_),
    .B(net71),
    .C(_04274_),
    .X(_04367_));
 sky130_fd_sc_hd__a31o_1 _18632_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net1085),
    .B1(_04367_),
    .X(_02061_));
 sky130_fd_sc_hd__nor2_1 _18633_ (.A(_09208_),
    .B(_04358_),
    .Y(_04368_));
 sky130_fd_sc_hd__a31o_1 _18634_ (.A1(_04235_),
    .A2(net1499),
    .A3(_04354_),
    .B1(_04368_),
    .X(_02062_));
 sky130_fd_sc_hd__and3_1 _18635_ (.A(_04350_),
    .B(net74),
    .C(_04274_),
    .X(_04369_));
 sky130_fd_sc_hd__a31o_1 _18636_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net1389),
    .B1(_04369_),
    .X(_02063_));
 sky130_fd_sc_hd__nand2_1 _18637_ (.A(_04336_),
    .B(net3141),
    .Y(_04370_));
 sky130_fd_sc_hd__a22o_1 _18638_ (.A1(_04357_),
    .A2(net135),
    .B1(_04358_),
    .B2(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__inv_2 _18639_ (.A(_04371_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand2_1 _18640_ (.A(_04336_),
    .B(net3426),
    .Y(_04372_));
 sky130_fd_sc_hd__a22o_1 _18641_ (.A1(_04357_),
    .A2(_09218_),
    .B1(_04358_),
    .B2(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__inv_2 _18642_ (.A(_04373_),
    .Y(_02049_));
 sky130_fd_sc_hd__nand2_1 _18643_ (.A(_04336_),
    .B(net3333),
    .Y(_04374_));
 sky130_fd_sc_hd__a22o_1 _18644_ (.A1(_04357_),
    .A2(_02963_),
    .B1(_04358_),
    .B2(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__inv_2 _18645_ (.A(_04375_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _18646_ (.A(_04336_),
    .B(net2895),
    .Y(_04376_));
 sky130_fd_sc_hd__a22o_1 _18647_ (.A1(_04357_),
    .A2(_09588_),
    .B1(_04358_),
    .B2(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__inv_2 _18648_ (.A(_04377_),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _18649_ (.A(_04336_),
    .B(net3051),
    .Y(_04378_));
 sky130_fd_sc_hd__a22o_1 _18650_ (.A1(_04357_),
    .A2(_09592_),
    .B1(_04358_),
    .B2(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__inv_2 _18651_ (.A(_04379_),
    .Y(_02052_));
 sky130_fd_sc_hd__nor2_1 _18652_ (.A(_09235_),
    .B(_04358_),
    .Y(_04380_));
 sky130_fd_sc_hd__a31o_1 _18653_ (.A1(_04235_),
    .A2(net819),
    .A3(_04354_),
    .B1(_04380_),
    .X(_02053_));
 sky130_fd_sc_hd__and3_1 _18654_ (.A(_04350_),
    .B(net64),
    .C(_04274_),
    .X(_04381_));
 sky130_fd_sc_hd__a31o_1 _18655_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net1071),
    .B1(_04381_),
    .X(_02054_));
 sky130_fd_sc_hd__nor2_1 _18656_ (.A(_09242_),
    .B(_04358_),
    .Y(_04382_));
 sky130_fd_sc_hd__a31o_1 _18657_ (.A1(_04235_),
    .A2(net1117),
    .A3(_04354_),
    .B1(_04382_),
    .X(_02055_));
 sky130_fd_sc_hd__nand2_1 _18658_ (.A(_04336_),
    .B(net3371),
    .Y(_04383_));
 sky130_fd_sc_hd__a22o_1 _18659_ (.A1(_04357_),
    .A2(net138),
    .B1(_04358_),
    .B2(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__inv_2 _18660_ (.A(_04384_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _18661_ (.A(_04336_),
    .B(net2974),
    .Y(_04385_));
 sky130_fd_sc_hd__a22o_1 _18662_ (.A1(_04357_),
    .A2(_09248_),
    .B1(_04358_),
    .B2(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__inv_2 _18663_ (.A(_04386_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _18664_ (.A(_04336_),
    .B(net2946),
    .Y(_04387_));
 sky130_fd_sc_hd__a22o_1 _18665_ (.A1(_04357_),
    .A2(_09347_),
    .B1(_04358_),
    .B2(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__inv_2 _18666_ (.A(_04388_),
    .Y(_02042_));
 sky130_fd_sc_hd__clkbuf_8 _18667_ (.A(_04184_),
    .X(_04389_));
 sky130_fd_sc_hd__nand2_1 _18668_ (.A(_04389_),
    .B(net2864),
    .Y(_04390_));
 sky130_fd_sc_hd__a22o_1 _18669_ (.A1(_04357_),
    .A2(_09255_),
    .B1(_04358_),
    .B2(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__inv_2 _18670_ (.A(_04391_),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _18671_ (.A(_04389_),
    .B(net2856),
    .Y(_04392_));
 sky130_fd_sc_hd__a22o_1 _18672_ (.A1(_04357_),
    .A2(_11136_),
    .B1(_04353_),
    .B2(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__inv_2 _18673_ (.A(_04393_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand2_1 _18674_ (.A(_04389_),
    .B(net3373),
    .Y(_04394_));
 sky130_fd_sc_hd__a22o_1 _18675_ (.A1(_04357_),
    .A2(net145),
    .B1(_04353_),
    .B2(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__inv_2 _18676_ (.A(_04395_),
    .Y(_02045_));
 sky130_fd_sc_hd__and3_1 _18677_ (.A(_04350_),
    .B(net55),
    .C(_04274_),
    .X(_04396_));
 sky130_fd_sc_hd__a31o_1 _18678_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net1269),
    .B1(_04396_),
    .X(_02046_));
 sky130_fd_sc_hd__nand2_1 _18679_ (.A(_04389_),
    .B(net2987),
    .Y(_04397_));
 sky130_fd_sc_hd__a22o_1 _18680_ (.A1(_04357_),
    .A2(net144),
    .B1(_04353_),
    .B2(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__inv_2 _18681_ (.A(_04398_),
    .Y(_02047_));
 sky130_fd_sc_hd__and3_1 _18682_ (.A(_04350_),
    .B(_03196_),
    .C(_04274_),
    .X(_04399_));
 sky130_fd_sc_hd__a31o_1 _18683_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net499),
    .B1(_04399_),
    .X(_02032_));
 sky130_fd_sc_hd__nor2_1 _18684_ (.A(_03605_),
    .B(_04358_),
    .Y(_04400_));
 sky130_fd_sc_hd__a31o_1 _18685_ (.A1(_04235_),
    .A2(net2651),
    .A3(_04354_),
    .B1(_04400_),
    .X(_02033_));
 sky130_fd_sc_hd__and3_1 _18686_ (.A(_04350_),
    .B(_03199_),
    .C(_04274_),
    .X(_04401_));
 sky130_fd_sc_hd__a31o_1 _18687_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net1329),
    .B1(_04401_),
    .X(_02034_));
 sky130_fd_sc_hd__nand2_1 _18688_ (.A(_04389_),
    .B(net3703),
    .Y(_04402_));
 sky130_fd_sc_hd__a22o_1 _18689_ (.A1(_04357_),
    .A2(net140),
    .B1(_04353_),
    .B2(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__inv_2 _18690_ (.A(_04403_),
    .Y(_02035_));
 sky130_fd_sc_hd__and3_1 _18691_ (.A(_04350_),
    .B(_03550_),
    .C(_04274_),
    .X(_04404_));
 sky130_fd_sc_hd__a31o_1 _18692_ (.A1(_04354_),
    .A2(_04365_),
    .A3(net1477),
    .B1(_04404_),
    .X(_02036_));
 sky130_fd_sc_hd__nand2_1 _18693_ (.A(_04221_),
    .B(net3799),
    .Y(_04405_));
 sky130_fd_sc_hd__o2bb2a_1 _18694_ (.A1_N(_04405_),
    .A2_N(_04354_),
    .B1(_09294_),
    .B2(_04351_),
    .X(_02037_));
 sky130_fd_sc_hd__nand2_1 _18695_ (.A(_04221_),
    .B(net3995),
    .Y(_04406_));
 sky130_fd_sc_hd__o2bb2a_1 _18696_ (.A1_N(_04406_),
    .A2_N(_04354_),
    .B1(_02992_),
    .B2(_04351_),
    .X(_02038_));
 sky130_fd_sc_hd__nand2_1 _18697_ (.A(_08777_),
    .B(net2878),
    .Y(_04407_));
 sky130_fd_sc_hd__a32o_1 _18698_ (.A1(_04356_),
    .A2(_08791_),
    .A3(_09299_),
    .B1(_04353_),
    .B2(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__inv_2 _18699_ (.A(net2879),
    .Y(_02039_));
 sky130_fd_sc_hd__and3_4 _18700_ (.A(_09511_),
    .B(_09444_),
    .C(_09380_),
    .X(_04409_));
 sky130_fd_sc_hd__inv_2 _18701_ (.A(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nor2_1 _18702_ (.A(_09304_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__inv_2 _18703_ (.A(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__buf_4 _18704_ (.A(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__buf_4 _18705_ (.A(_04412_),
    .X(_04414_));
 sky130_fd_sc_hd__nor2_1 _18706_ (.A(_09180_),
    .B(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__a31o_1 _18707_ (.A1(_04235_),
    .A2(net1533),
    .A3(_04413_),
    .B1(_04415_),
    .X(_02016_));
 sky130_fd_sc_hd__nor2_1 _18708_ (.A(_03170_),
    .B(_04414_),
    .Y(_04416_));
 sky130_fd_sc_hd__a31o_1 _18709_ (.A1(_04235_),
    .A2(net1215),
    .A3(_04413_),
    .B1(_04416_),
    .X(_02017_));
 sky130_fd_sc_hd__clkbuf_8 _18710_ (.A(_09164_),
    .X(_04417_));
 sky130_fd_sc_hd__nor2_1 _18711_ (.A(_03219_),
    .B(_04414_),
    .Y(_04418_));
 sky130_fd_sc_hd__a31o_1 _18712_ (.A1(_04417_),
    .A2(net795),
    .A3(_04413_),
    .B1(_04418_),
    .X(_02018_));
 sky130_fd_sc_hd__and3_1 _18713_ (.A(_04409_),
    .B(net69),
    .C(_04274_),
    .X(_04419_));
 sky130_fd_sc_hd__a31o_1 _18714_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net1890),
    .B1(_04419_),
    .X(_02019_));
 sky130_fd_sc_hd__nor2_4 _18715_ (.A(_08795_),
    .B(_04410_),
    .Y(_04420_));
 sky130_fd_sc_hd__nand2_1 _18716_ (.A(_04389_),
    .B(net2930),
    .Y(_04421_));
 sky130_fd_sc_hd__a22o_1 _18717_ (.A1(_04420_),
    .A2(_11330_),
    .B1(_04414_),
    .B2(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__inv_2 _18718_ (.A(_04422_),
    .Y(_02020_));
 sky130_fd_sc_hd__and3_1 _18719_ (.A(_04409_),
    .B(net71),
    .C(_04274_),
    .X(_04423_));
 sky130_fd_sc_hd__a31o_1 _18720_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net2148),
    .B1(_04423_),
    .X(_02021_));
 sky130_fd_sc_hd__nor2_1 _18721_ (.A(_09208_),
    .B(_04414_),
    .Y(_04424_));
 sky130_fd_sc_hd__a31o_1 _18722_ (.A1(_04417_),
    .A2(net1197),
    .A3(_04413_),
    .B1(_04424_),
    .X(_02022_));
 sky130_fd_sc_hd__and3_1 _18723_ (.A(_04409_),
    .B(net74),
    .C(_04274_),
    .X(_04425_));
 sky130_fd_sc_hd__a31o_1 _18724_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net2348),
    .B1(_04425_),
    .X(_02023_));
 sky130_fd_sc_hd__nor2_1 _18725_ (.A(_03467_),
    .B(_04414_),
    .Y(_04426_));
 sky130_fd_sc_hd__a31o_1 _18726_ (.A1(_04417_),
    .A2(net2464),
    .A3(_04414_),
    .B1(_04426_),
    .X(_02008_));
 sky130_fd_sc_hd__nand2_1 _18727_ (.A(_04389_),
    .B(net2948),
    .Y(_04427_));
 sky130_fd_sc_hd__a22o_1 _18728_ (.A1(_04420_),
    .A2(_09218_),
    .B1(_04414_),
    .B2(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__inv_2 _18729_ (.A(_04428_),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _18730_ (.A(_04389_),
    .B(net3711),
    .Y(_04429_));
 sky130_fd_sc_hd__a22o_1 _18731_ (.A1(_04420_),
    .A2(net143),
    .B1(_04412_),
    .B2(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__inv_2 _18732_ (.A(_04430_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _18733_ (.A(_04389_),
    .B(net2988),
    .Y(_04431_));
 sky130_fd_sc_hd__a22o_1 _18734_ (.A1(_04420_),
    .A2(_09588_),
    .B1(_04412_),
    .B2(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__inv_2 _18735_ (.A(_04432_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _18736_ (.A(_04389_),
    .B(net3397),
    .Y(_04433_));
 sky130_fd_sc_hd__a22o_1 _18737_ (.A1(_04420_),
    .A2(_09592_),
    .B1(_04412_),
    .B2(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__inv_2 _18738_ (.A(_04434_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_1 _18739_ (.A(_09235_),
    .B(_04414_),
    .Y(_04435_));
 sky130_fd_sc_hd__a31o_1 _18740_ (.A1(_04417_),
    .A2(net881),
    .A3(_04414_),
    .B1(_04435_),
    .X(_02013_));
 sky130_fd_sc_hd__and3_1 _18741_ (.A(_04409_),
    .B(net64),
    .C(_04274_),
    .X(_04436_));
 sky130_fd_sc_hd__a31o_1 _18742_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net1399),
    .B1(_04436_),
    .X(_02014_));
 sky130_fd_sc_hd__nor2_1 _18743_ (.A(_09242_),
    .B(_04414_),
    .Y(_04437_));
 sky130_fd_sc_hd__a31o_1 _18744_ (.A1(_04417_),
    .A2(net855),
    .A3(_04414_),
    .B1(_04437_),
    .X(_02015_));
 sky130_fd_sc_hd__nand2_1 _18745_ (.A(_04389_),
    .B(net3559),
    .Y(_04438_));
 sky130_fd_sc_hd__a22o_1 _18746_ (.A1(_04420_),
    .A2(_09414_),
    .B1(_04412_),
    .B2(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__inv_2 _18747_ (.A(_04439_),
    .Y(_02000_));
 sky130_fd_sc_hd__and3_1 _18748_ (.A(_04409_),
    .B(net82),
    .C(_04274_),
    .X(_04440_));
 sky130_fd_sc_hd__a31o_1 _18749_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net2256),
    .B1(_04440_),
    .X(_02001_));
 sky130_fd_sc_hd__nor2_1 _18750_ (.A(_03482_),
    .B(_04414_),
    .Y(_04441_));
 sky130_fd_sc_hd__a31o_1 _18751_ (.A1(_04417_),
    .A2(net655),
    .A3(_04414_),
    .B1(_04441_),
    .X(_02002_));
 sky130_fd_sc_hd__and3_1 _18752_ (.A(_04409_),
    .B(net52),
    .C(_04274_),
    .X(_04442_));
 sky130_fd_sc_hd__a31o_1 _18753_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net1753),
    .B1(_04442_),
    .X(_02003_));
 sky130_fd_sc_hd__nor2_1 _18754_ (.A(_09259_),
    .B(_04414_),
    .Y(_04443_));
 sky130_fd_sc_hd__a31o_1 _18755_ (.A1(_04417_),
    .A2(net777),
    .A3(_04414_),
    .B1(_04443_),
    .X(_02004_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(_04389_),
    .B(net3688),
    .Y(_04444_));
 sky130_fd_sc_hd__a22o_1 _18757_ (.A1(_04420_),
    .A2(_09262_),
    .B1(_04412_),
    .B2(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__inv_2 _18758_ (.A(_04445_),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _18759_ (.A(_04389_),
    .B(net2823),
    .Y(_04446_));
 sky130_fd_sc_hd__a22o_1 _18760_ (.A1(_04420_),
    .A2(_09424_),
    .B1(_04412_),
    .B2(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__inv_2 _18761_ (.A(_04447_),
    .Y(_02006_));
 sky130_fd_sc_hd__nand2_1 _18762_ (.A(_04389_),
    .B(net3654),
    .Y(_04448_));
 sky130_fd_sc_hd__a22o_1 _18763_ (.A1(_04420_),
    .A2(_09268_),
    .B1(_04412_),
    .B2(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__inv_2 _18764_ (.A(_04449_),
    .Y(_02007_));
 sky130_fd_sc_hd__buf_4 _18765_ (.A(_09226_),
    .X(_04450_));
 sky130_fd_sc_hd__and3_1 _18766_ (.A(_04409_),
    .B(_03196_),
    .C(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__a31o_1 _18767_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net1407),
    .B1(_04451_),
    .X(_01992_));
 sky130_fd_sc_hd__nand2_1 _18768_ (.A(_04389_),
    .B(net2973),
    .Y(_04452_));
 sky130_fd_sc_hd__a22o_1 _18769_ (.A1(_04420_),
    .A2(_09365_),
    .B1(_04412_),
    .B2(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__inv_2 _18770_ (.A(_04453_),
    .Y(_01993_));
 sky130_fd_sc_hd__and3_1 _18771_ (.A(_04409_),
    .B(_03199_),
    .C(_04450_),
    .X(_04454_));
 sky130_fd_sc_hd__a31o_1 _18772_ (.A1(_04413_),
    .A2(_04365_),
    .A3(net1491),
    .B1(_04454_),
    .X(_01994_));
 sky130_fd_sc_hd__nand2_1 _18773_ (.A(_04389_),
    .B(net3719),
    .Y(_04455_));
 sky130_fd_sc_hd__a22o_1 _18774_ (.A1(_04420_),
    .A2(net140),
    .B1(_04412_),
    .B2(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__inv_2 _18775_ (.A(_04456_),
    .Y(_01995_));
 sky130_fd_sc_hd__clkbuf_8 _18776_ (.A(_03834_),
    .X(_04457_));
 sky130_fd_sc_hd__and3_1 _18777_ (.A(_04409_),
    .B(_03550_),
    .C(_04450_),
    .X(_04458_));
 sky130_fd_sc_hd__a31o_1 _18778_ (.A1(_04413_),
    .A2(_04457_),
    .A3(net2325),
    .B1(_04458_),
    .X(_01996_));
 sky130_fd_sc_hd__nand2_1 _18779_ (.A(_04221_),
    .B(net3886),
    .Y(_04459_));
 sky130_fd_sc_hd__o2bb2a_1 _18780_ (.A1_N(_04459_),
    .A2_N(_04413_),
    .B1(_09293_),
    .B2(_04410_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _18781_ (.A(_04221_),
    .B(net3639),
    .Y(_04460_));
 sky130_fd_sc_hd__o2bb2a_1 _18782_ (.A1_N(_04460_),
    .A2_N(_04413_),
    .B1(_09297_),
    .B2(_04410_),
    .X(_01998_));
 sky130_fd_sc_hd__nand2_1 _18783_ (.A(_04221_),
    .B(net3598),
    .Y(_04461_));
 sky130_fd_sc_hd__o2bb2a_1 _18784_ (.A1_N(_04461_),
    .A2_N(_04413_),
    .B1(_11316_),
    .B2(_04410_),
    .X(_01999_));
 sky130_fd_sc_hd__nor2_2 _18785_ (.A(_08736_),
    .B(_09677_),
    .Y(_04462_));
 sky130_fd_sc_hd__inv_2 _18786_ (.A(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__nor2_2 _18787_ (.A(_08794_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__buf_4 _18788_ (.A(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__nor2_1 _18789_ (.A(_08728_),
    .B(_04463_),
    .Y(_04466_));
 sky130_fd_sc_hd__inv_2 _18790_ (.A(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__buf_4 _18791_ (.A(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__buf_4 _18792_ (.A(_04184_),
    .X(_04469_));
 sky130_fd_sc_hd__nand2_1 _18793_ (.A(_04469_),
    .B(net2796),
    .Y(_04470_));
 sky130_fd_sc_hd__a22o_1 _18794_ (.A1(_04465_),
    .A2(_10239_),
    .B1(_04468_),
    .B2(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__inv_2 _18795_ (.A(_04471_),
    .Y(_01984_));
 sky130_fd_sc_hd__buf_4 _18796_ (.A(_04467_),
    .X(_04472_));
 sky130_fd_sc_hd__nor2_1 _18797_ (.A(_03170_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__a31o_1 _18798_ (.A1(_04417_),
    .A2(net1271),
    .A3(_04472_),
    .B1(_04473_),
    .X(_01985_));
 sky130_fd_sc_hd__nor2_1 _18799_ (.A(_03219_),
    .B(_04472_),
    .Y(_04474_));
 sky130_fd_sc_hd__a31o_1 _18800_ (.A1(_04417_),
    .A2(net1647),
    .A3(_04472_),
    .B1(_04474_),
    .X(_01986_));
 sky130_fd_sc_hd__nand2_1 _18801_ (.A(_04469_),
    .B(net2881),
    .Y(_04475_));
 sky130_fd_sc_hd__a22o_1 _18802_ (.A1(_04465_),
    .A2(_10983_),
    .B1(_04468_),
    .B2(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__inv_2 _18803_ (.A(_04476_),
    .Y(_01987_));
 sky130_fd_sc_hd__nand2_1 _18804_ (.A(_04469_),
    .B(net3576),
    .Y(_04477_));
 sky130_fd_sc_hd__a22o_1 _18805_ (.A1(_04465_),
    .A2(_11330_),
    .B1(_04468_),
    .B2(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__inv_2 _18806_ (.A(_04478_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand2_1 _18807_ (.A(_04469_),
    .B(net3357),
    .Y(_04479_));
 sky130_fd_sc_hd__a22o_1 _18808_ (.A1(_04465_),
    .A2(_09204_),
    .B1(_04468_),
    .B2(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__inv_2 _18809_ (.A(_04480_),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_1 _18810_ (.A(_04469_),
    .B(net3050),
    .Y(_04481_));
 sky130_fd_sc_hd__a22o_1 _18811_ (.A1(_04465_),
    .A2(_11105_),
    .B1(_04468_),
    .B2(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__inv_2 _18812_ (.A(_04482_),
    .Y(_01990_));
 sky130_fd_sc_hd__nand2_1 _18813_ (.A(_04469_),
    .B(net3454),
    .Y(_04483_));
 sky130_fd_sc_hd__a22o_1 _18814_ (.A1(_04465_),
    .A2(_09211_),
    .B1(_04468_),
    .B2(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__inv_2 _18815_ (.A(_04484_),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_1 _18816_ (.A(_03467_),
    .B(_04472_),
    .Y(_04485_));
 sky130_fd_sc_hd__a31o_1 _18817_ (.A1(_04417_),
    .A2(net1097),
    .A3(_04472_),
    .B1(_04485_),
    .X(_01976_));
 sky130_fd_sc_hd__nand2_1 _18818_ (.A(_04469_),
    .B(net2966),
    .Y(_04486_));
 sky130_fd_sc_hd__a22o_1 _18819_ (.A1(_04465_),
    .A2(_09218_),
    .B1(_04468_),
    .B2(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__inv_2 _18820_ (.A(_04487_),
    .Y(_01977_));
 sky130_fd_sc_hd__nand2_1 _18821_ (.A(_04469_),
    .B(net3046),
    .Y(_04488_));
 sky130_fd_sc_hd__a22o_1 _18822_ (.A1(_04465_),
    .A2(net143),
    .B1(_04468_),
    .B2(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__inv_2 _18823_ (.A(_04489_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _18824_ (.A(_09229_),
    .B(_04472_),
    .Y(_04490_));
 sky130_fd_sc_hd__a31o_1 _18825_ (.A1(_04417_),
    .A2(net1822),
    .A3(_04472_),
    .B1(_04490_),
    .X(_01979_));
 sky130_fd_sc_hd__nand2_1 _18826_ (.A(_04469_),
    .B(net3289),
    .Y(_04491_));
 sky130_fd_sc_hd__a22o_1 _18827_ (.A1(_04465_),
    .A2(_09592_),
    .B1(_04468_),
    .B2(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__inv_2 _18828_ (.A(_04492_),
    .Y(_01980_));
 sky130_fd_sc_hd__nand2_1 _18829_ (.A(_04469_),
    .B(net3510),
    .Y(_04493_));
 sky130_fd_sc_hd__a22o_1 _18830_ (.A1(_04465_),
    .A2(_09337_),
    .B1(_04468_),
    .B2(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__inv_2 _18831_ (.A(_04494_),
    .Y(_01981_));
 sky130_fd_sc_hd__and3_1 _18832_ (.A(_04462_),
    .B(net64),
    .C(_04450_),
    .X(_04495_));
 sky130_fd_sc_hd__a31o_1 _18833_ (.A1(_04472_),
    .A2(_04457_),
    .A3(net2337),
    .B1(_04495_),
    .X(_01982_));
 sky130_fd_sc_hd__nand2_1 _18834_ (.A(_04469_),
    .B(net3686),
    .Y(_04496_));
 sky130_fd_sc_hd__a22o_1 _18835_ (.A1(_04465_),
    .A2(_09767_),
    .B1(_04468_),
    .B2(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__inv_2 _18836_ (.A(_04497_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _18837_ (.A(_03294_),
    .B(_04468_),
    .Y(_04498_));
 sky130_fd_sc_hd__a31o_1 _18838_ (.A1(_04417_),
    .A2(net875),
    .A3(_04472_),
    .B1(_04498_),
    .X(_01968_));
 sky130_fd_sc_hd__nand2_1 _18839_ (.A(_04469_),
    .B(net3535),
    .Y(_04499_));
 sky130_fd_sc_hd__a22o_1 _18840_ (.A1(_04465_),
    .A2(_09248_),
    .B1(_04468_),
    .B2(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__inv_2 _18841_ (.A(_04500_),
    .Y(_01969_));
 sky130_fd_sc_hd__nand2_1 _18842_ (.A(_04469_),
    .B(net3154),
    .Y(_04501_));
 sky130_fd_sc_hd__a22o_1 _18843_ (.A1(_04465_),
    .A2(_09347_),
    .B1(_04468_),
    .B2(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__inv_2 _18844_ (.A(_04502_),
    .Y(_01970_));
 sky130_fd_sc_hd__and3_1 _18845_ (.A(_04462_),
    .B(net52),
    .C(_04450_),
    .X(_04503_));
 sky130_fd_sc_hd__a31o_1 _18846_ (.A1(_04472_),
    .A2(_04457_),
    .A3(net1309),
    .B1(_04503_),
    .X(_01971_));
 sky130_fd_sc_hd__nand2_1 _18847_ (.A(_04469_),
    .B(net3503),
    .Y(_04504_));
 sky130_fd_sc_hd__a22o_1 _18848_ (.A1(_04465_),
    .A2(_11136_),
    .B1(_04468_),
    .B2(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__inv_2 _18849_ (.A(_04505_),
    .Y(_01972_));
 sky130_fd_sc_hd__nand2_1 _18850_ (.A(_04469_),
    .B(net3430),
    .Y(_04506_));
 sky130_fd_sc_hd__a22o_1 _18851_ (.A1(_04465_),
    .A2(_09262_),
    .B1(_04467_),
    .B2(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__inv_2 _18852_ (.A(_04507_),
    .Y(_01973_));
 sky130_fd_sc_hd__nand2_1 _18853_ (.A(_04469_),
    .B(net3482),
    .Y(_04508_));
 sky130_fd_sc_hd__a22o_1 _18854_ (.A1(_04465_),
    .A2(_09424_),
    .B1(_04467_),
    .B2(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__inv_2 _18855_ (.A(_04509_),
    .Y(_01974_));
 sky130_fd_sc_hd__buf_4 _18856_ (.A(_04184_),
    .X(_04510_));
 sky130_fd_sc_hd__nand2_1 _18857_ (.A(_04510_),
    .B(net3105),
    .Y(_04511_));
 sky130_fd_sc_hd__a22o_1 _18858_ (.A1(_04464_),
    .A2(_09268_),
    .B1(_04467_),
    .B2(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__inv_2 _18859_ (.A(_04512_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _18860_ (.A(_04510_),
    .B(net3558),
    .Y(_04513_));
 sky130_fd_sc_hd__a22o_1 _18861_ (.A1(_04464_),
    .A2(_09494_),
    .B1(_04467_),
    .B2(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__inv_2 _18862_ (.A(_04514_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2_1 _18863_ (.A(_03605_),
    .B(_04468_),
    .Y(_04515_));
 sky130_fd_sc_hd__a31o_1 _18864_ (.A1(_04417_),
    .A2(net2635),
    .A3(_04472_),
    .B1(_04515_),
    .X(_01961_));
 sky130_fd_sc_hd__and3_1 _18865_ (.A(_04462_),
    .B(_03199_),
    .C(_04450_),
    .X(_04516_));
 sky130_fd_sc_hd__a31o_1 _18866_ (.A1(_04472_),
    .A2(_04457_),
    .A3(net2602),
    .B1(_04516_),
    .X(_01962_));
 sky130_fd_sc_hd__nand2_1 _18867_ (.A(_04510_),
    .B(net3522),
    .Y(_04517_));
 sky130_fd_sc_hd__a22o_1 _18868_ (.A1(_04464_),
    .A2(net140),
    .B1(_04467_),
    .B2(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__inv_2 _18869_ (.A(_04518_),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_1 _18870_ (.A(_04510_),
    .B(net2934),
    .Y(_04519_));
 sky130_fd_sc_hd__a22o_1 _18871_ (.A1(_04464_),
    .A2(_09287_),
    .B1(_04467_),
    .B2(_04519_),
    .X(_04520_));
 sky130_fd_sc_hd__inv_2 _18872_ (.A(_04520_),
    .Y(_01964_));
 sky130_fd_sc_hd__and3_1 _18873_ (.A(_04462_),
    .B(net78),
    .C(_04450_),
    .X(_04521_));
 sky130_fd_sc_hd__a31o_1 _18874_ (.A1(_04472_),
    .A2(_04457_),
    .A3(net1589),
    .B1(_04521_),
    .X(_01965_));
 sky130_fd_sc_hd__nand2_1 _18875_ (.A(_04221_),
    .B(net3823),
    .Y(_04522_));
 sky130_fd_sc_hd__o2bb2a_1 _18876_ (.A1_N(_04522_),
    .A2_N(_04472_),
    .B1(_09297_),
    .B2(_04463_),
    .X(_01966_));
 sky130_fd_sc_hd__nand2_1 _18877_ (.A(_04221_),
    .B(net3829),
    .Y(_04523_));
 sky130_fd_sc_hd__o2bb2a_1 _18878_ (.A1_N(_04523_),
    .A2_N(_04472_),
    .B1(_09441_),
    .B2(_04463_),
    .X(_01967_));
 sky130_fd_sc_hd__nor2_2 _18879_ (.A(_08736_),
    .B(_09738_),
    .Y(_04524_));
 sky130_fd_sc_hd__inv_2 _18880_ (.A(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2_1 _18881_ (.A(_09166_),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__clkinv_4 _18882_ (.A(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__buf_4 _18883_ (.A(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__buf_4 _18884_ (.A(_04527_),
    .X(_04529_));
 sky130_fd_sc_hd__nor2_1 _18885_ (.A(_09180_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__a31o_1 _18886_ (.A1(_04417_),
    .A2(net2479),
    .A3(_04528_),
    .B1(_04530_),
    .X(_01952_));
 sky130_fd_sc_hd__nor2_4 _18887_ (.A(_09190_),
    .B(_04525_),
    .Y(_04531_));
 sky130_fd_sc_hd__nand2_1 _18888_ (.A(_04510_),
    .B(net3811),
    .Y(_04532_));
 sky130_fd_sc_hd__a22o_1 _18889_ (.A1(_04531_),
    .A2(_09314_),
    .B1(_04527_),
    .B2(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__inv_2 _18890_ (.A(_04533_),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _18891_ (.A(_03219_),
    .B(_04529_),
    .Y(_04534_));
 sky130_fd_sc_hd__a31o_1 _18892_ (.A1(_04417_),
    .A2(net613),
    .A3(_04528_),
    .B1(_04534_),
    .X(_01954_));
 sky130_fd_sc_hd__nand2_1 _18893_ (.A(_04510_),
    .B(net3798),
    .Y(_04535_));
 sky130_fd_sc_hd__a22o_1 _18894_ (.A1(_04531_),
    .A2(_10983_),
    .B1(_04527_),
    .B2(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__inv_2 _18895_ (.A(_04536_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _18896_ (.A(_04510_),
    .B(net3891),
    .Y(_04537_));
 sky130_fd_sc_hd__a22o_1 _18897_ (.A1(_04531_),
    .A2(_11330_),
    .B1(_04527_),
    .B2(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__inv_2 _18898_ (.A(_04538_),
    .Y(_01956_));
 sky130_fd_sc_hd__and3_1 _18899_ (.A(_04524_),
    .B(net71),
    .C(_04450_),
    .X(_04539_));
 sky130_fd_sc_hd__a31o_1 _18900_ (.A1(_04528_),
    .A2(_04457_),
    .A3(net2601),
    .B1(_04539_),
    .X(_01957_));
 sky130_fd_sc_hd__nor2_1 _18901_ (.A(_09208_),
    .B(_04529_),
    .Y(_04540_));
 sky130_fd_sc_hd__a31o_1 _18902_ (.A1(_04417_),
    .A2(net2350),
    .A3(_04528_),
    .B1(_04540_),
    .X(_01958_));
 sky130_fd_sc_hd__and3_1 _18903_ (.A(_04524_),
    .B(net74),
    .C(_04450_),
    .X(_04541_));
 sky130_fd_sc_hd__a31o_1 _18904_ (.A1(_04528_),
    .A2(_04457_),
    .A3(net2577),
    .B1(_04541_),
    .X(_01959_));
 sky130_fd_sc_hd__buf_4 _18905_ (.A(_09164_),
    .X(_04542_));
 sky130_fd_sc_hd__nor2_1 _18906_ (.A(_03467_),
    .B(_04529_),
    .Y(_04543_));
 sky130_fd_sc_hd__a31o_1 _18907_ (.A1(_04542_),
    .A2(net497),
    .A3(_04528_),
    .B1(_04543_),
    .X(_01864_));
 sky130_fd_sc_hd__nand2_1 _18908_ (.A(_04510_),
    .B(net3384),
    .Y(_04544_));
 sky130_fd_sc_hd__a22o_1 _18909_ (.A1(_04531_),
    .A2(net146),
    .B1(_04527_),
    .B2(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__inv_2 _18910_ (.A(_04545_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _18911_ (.A(_04510_),
    .B(net2950),
    .Y(_04546_));
 sky130_fd_sc_hd__a22o_1 _18912_ (.A1(_04531_),
    .A2(net143),
    .B1(_04527_),
    .B2(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__inv_2 _18913_ (.A(_04547_),
    .Y(_01866_));
 sky130_fd_sc_hd__nor2_1 _18914_ (.A(_09229_),
    .B(_04529_),
    .Y(_04548_));
 sky130_fd_sc_hd__a31o_1 _18915_ (.A1(_04542_),
    .A2(net1109),
    .A3(_04528_),
    .B1(_04548_),
    .X(_01867_));
 sky130_fd_sc_hd__nor2_1 _18916_ (.A(_09232_),
    .B(_04529_),
    .Y(_04549_));
 sky130_fd_sc_hd__a31o_1 _18917_ (.A1(_04542_),
    .A2(net2176),
    .A3(_04528_),
    .B1(_04549_),
    .X(_01868_));
 sky130_fd_sc_hd__nor2_1 _18918_ (.A(_09235_),
    .B(_04529_),
    .Y(_04550_));
 sky130_fd_sc_hd__a31o_1 _18919_ (.A1(_04542_),
    .A2(net1351),
    .A3(_04528_),
    .B1(_04550_),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_1 _18920_ (.A(_04510_),
    .B(net3729),
    .Y(_04551_));
 sky130_fd_sc_hd__a22o_1 _18921_ (.A1(_04531_),
    .A2(_09238_),
    .B1(_04527_),
    .B2(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__inv_2 _18922_ (.A(_04552_),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _18923_ (.A(_04510_),
    .B(net3379),
    .Y(_04553_));
 sky130_fd_sc_hd__a22o_1 _18924_ (.A1(_04531_),
    .A2(_09767_),
    .B1(_04527_),
    .B2(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__inv_2 _18925_ (.A(_04554_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _18926_ (.A(_03294_),
    .B(_04529_),
    .Y(_04555_));
 sky130_fd_sc_hd__a31o_1 _18927_ (.A1(_04542_),
    .A2(net1429),
    .A3(_04528_),
    .B1(_04555_),
    .X(_01768_));
 sky130_fd_sc_hd__nand2_1 _18928_ (.A(_04510_),
    .B(net3016),
    .Y(_04556_));
 sky130_fd_sc_hd__a22o_1 _18929_ (.A1(_04531_),
    .A2(_09248_),
    .B1(_04527_),
    .B2(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__inv_2 _18930_ (.A(_04557_),
    .Y(_01769_));
 sky130_fd_sc_hd__nor2_1 _18931_ (.A(_03482_),
    .B(_04529_),
    .Y(_04558_));
 sky130_fd_sc_hd__a31o_1 _18932_ (.A1(_04542_),
    .A2(net2082),
    .A3(_04529_),
    .B1(_04558_),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_1 _18933_ (.A(_04510_),
    .B(net3069),
    .Y(_04559_));
 sky130_fd_sc_hd__a22o_1 _18934_ (.A1(_04531_),
    .A2(_09255_),
    .B1(_04527_),
    .B2(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__inv_2 _18935_ (.A(_04560_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _18936_ (.A(_09259_),
    .B(_04529_),
    .Y(_04561_));
 sky130_fd_sc_hd__a31o_1 _18937_ (.A1(_04542_),
    .A2(net799),
    .A3(_04529_),
    .B1(_04561_),
    .X(_01772_));
 sky130_fd_sc_hd__nand2_1 _18938_ (.A(_04510_),
    .B(net2940),
    .Y(_04562_));
 sky130_fd_sc_hd__a22o_1 _18939_ (.A1(_04531_),
    .A2(net145),
    .B1(_04527_),
    .B2(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__inv_2 _18940_ (.A(_04563_),
    .Y(_01773_));
 sky130_fd_sc_hd__and3_1 _18941_ (.A(_04524_),
    .B(net55),
    .C(_04450_),
    .X(_04564_));
 sky130_fd_sc_hd__a31o_1 _18942_ (.A1(_04528_),
    .A2(_04457_),
    .A3(net1373),
    .B1(_04564_),
    .X(_01774_));
 sky130_fd_sc_hd__nand2_1 _18943_ (.A(_04510_),
    .B(net3082),
    .Y(_04565_));
 sky130_fd_sc_hd__a22o_1 _18944_ (.A1(_04531_),
    .A2(net144),
    .B1(_04527_),
    .B2(_04565_),
    .X(_04566_));
 sky130_fd_sc_hd__inv_2 _18945_ (.A(_04566_),
    .Y(_01775_));
 sky130_fd_sc_hd__and3_1 _18946_ (.A(_04524_),
    .B(_03196_),
    .C(_04450_),
    .X(_04567_));
 sky130_fd_sc_hd__a31o_1 _18947_ (.A1(_04528_),
    .A2(_04457_),
    .A3(net615),
    .B1(_04567_),
    .X(_01680_));
 sky130_fd_sc_hd__nor2_1 _18948_ (.A(_03605_),
    .B(_04529_),
    .Y(_04568_));
 sky130_fd_sc_hd__a31o_1 _18949_ (.A1(_04542_),
    .A2(net2461),
    .A3(_04529_),
    .B1(_04568_),
    .X(_01681_));
 sky130_fd_sc_hd__and3_1 _18950_ (.A(_04524_),
    .B(_03199_),
    .C(_04450_),
    .X(_04569_));
 sky130_fd_sc_hd__a31o_1 _18951_ (.A1(_04528_),
    .A2(_04457_),
    .A3(net1780),
    .B1(_04569_),
    .X(_01682_));
 sky130_fd_sc_hd__nand2_1 _18952_ (.A(_04510_),
    .B(net3196),
    .Y(_04570_));
 sky130_fd_sc_hd__a22o_1 _18953_ (.A1(_04531_),
    .A2(net140),
    .B1(_04527_),
    .B2(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__inv_2 _18954_ (.A(_04571_),
    .Y(_01683_));
 sky130_fd_sc_hd__and3_1 _18955_ (.A(_04524_),
    .B(_03550_),
    .C(_04450_),
    .X(_04572_));
 sky130_fd_sc_hd__a31o_1 _18956_ (.A1(_04528_),
    .A2(_04457_),
    .A3(net1463),
    .B1(_04572_),
    .X(_01684_));
 sky130_fd_sc_hd__and3_1 _18957_ (.A(_04524_),
    .B(net78),
    .C(_04450_),
    .X(_04573_));
 sky130_fd_sc_hd__a31o_1 _18958_ (.A1(_04528_),
    .A2(_04457_),
    .A3(net1671),
    .B1(_04573_),
    .X(_01685_));
 sky130_fd_sc_hd__nand2_1 _18959_ (.A(_04221_),
    .B(net3620),
    .Y(_04574_));
 sky130_fd_sc_hd__o2bb2a_1 _18960_ (.A1_N(_04574_),
    .A2_N(_04528_),
    .B1(_09297_),
    .B2(_04525_),
    .X(_01686_));
 sky130_fd_sc_hd__nor2_1 _18961_ (.A(_09299_),
    .B(_04529_),
    .Y(_04575_));
 sky130_fd_sc_hd__a31o_1 _18962_ (.A1(_04542_),
    .A2(net1645),
    .A3(_04529_),
    .B1(_04575_),
    .X(_01687_));
 sky130_fd_sc_hd__and3_4 _18963_ (.A(_09737_),
    .B(_09444_),
    .C(_09305_),
    .X(_04576_));
 sky130_fd_sc_hd__inv_2 _18964_ (.A(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__nor2_1 _18965_ (.A(_09166_),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__clkinv_4 _18966_ (.A(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__buf_4 _18967_ (.A(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__buf_4 _18968_ (.A(_04579_),
    .X(_04581_));
 sky130_fd_sc_hd__nor2_1 _18969_ (.A(_09180_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__a31o_1 _18970_ (.A1(_04542_),
    .A2(net2115),
    .A3(_04580_),
    .B1(_04582_),
    .X(_01592_));
 sky130_fd_sc_hd__nor2_1 _18971_ (.A(_03170_),
    .B(_04581_),
    .Y(_04583_));
 sky130_fd_sc_hd__a31o_1 _18972_ (.A1(_04542_),
    .A2(net2709),
    .A3(_04580_),
    .B1(_04583_),
    .X(_01593_));
 sky130_fd_sc_hd__nor2_1 _18973_ (.A(_03219_),
    .B(_04581_),
    .Y(_04584_));
 sky130_fd_sc_hd__a31o_1 _18974_ (.A1(_04542_),
    .A2(net2710),
    .A3(_04580_),
    .B1(_04584_),
    .X(_01594_));
 sky130_fd_sc_hd__nor2_4 _18975_ (.A(_08797_),
    .B(_04577_),
    .Y(_04585_));
 sky130_fd_sc_hd__buf_4 _18976_ (.A(_04184_),
    .X(_04586_));
 sky130_fd_sc_hd__nand2_1 _18977_ (.A(_04586_),
    .B(net4275),
    .Y(_04587_));
 sky130_fd_sc_hd__a22o_1 _18978_ (.A1(_04585_),
    .A2(_10983_),
    .B1(_04581_),
    .B2(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__inv_2 _18979_ (.A(_04588_),
    .Y(_01595_));
 sky130_fd_sc_hd__and3_1 _18980_ (.A(_04576_),
    .B(_10586_),
    .C(_04450_),
    .X(_04589_));
 sky130_fd_sc_hd__a31o_1 _18981_ (.A1(_04580_),
    .A2(_04457_),
    .A3(net2563),
    .B1(_04589_),
    .X(_01596_));
 sky130_fd_sc_hd__and3_1 _18982_ (.A(_04576_),
    .B(net71),
    .C(_04450_),
    .X(_04590_));
 sky130_fd_sc_hd__a31o_1 _18983_ (.A1(_04580_),
    .A2(_04457_),
    .A3(net2605),
    .B1(_04590_),
    .X(_01597_));
 sky130_fd_sc_hd__nor2_1 _18984_ (.A(_09208_),
    .B(_04581_),
    .Y(_04591_));
 sky130_fd_sc_hd__a31o_1 _18985_ (.A1(_04542_),
    .A2(net1680),
    .A3(_04580_),
    .B1(_04591_),
    .X(_01598_));
 sky130_fd_sc_hd__nand2_1 _18986_ (.A(_04586_),
    .B(net3841),
    .Y(_04592_));
 sky130_fd_sc_hd__a22o_1 _18987_ (.A1(_04585_),
    .A2(_09211_),
    .B1(_04581_),
    .B2(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__inv_2 _18988_ (.A(_04593_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand2_1 _18989_ (.A(_04586_),
    .B(net3774),
    .Y(_04594_));
 sky130_fd_sc_hd__a22o_1 _18990_ (.A1(_04585_),
    .A2(net135),
    .B1(_04581_),
    .B2(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__inv_2 _18991_ (.A(_04595_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _18992_ (.A(_04586_),
    .B(net4272),
    .Y(_04596_));
 sky130_fd_sc_hd__a22o_1 _18993_ (.A1(_04585_),
    .A2(_09218_),
    .B1(_04581_),
    .B2(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__inv_2 _18994_ (.A(_04597_),
    .Y(_01505_));
 sky130_fd_sc_hd__nand2_1 _18995_ (.A(_04586_),
    .B(net4261),
    .Y(_04598_));
 sky130_fd_sc_hd__a22o_1 _18996_ (.A1(_04585_),
    .A2(net143),
    .B1(_04579_),
    .B2(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__inv_2 _18997_ (.A(_04599_),
    .Y(_01506_));
 sky130_fd_sc_hd__nand2_1 _18998_ (.A(_04586_),
    .B(net4283),
    .Y(_04600_));
 sky130_fd_sc_hd__a22o_1 _18999_ (.A1(_04585_),
    .A2(_09588_),
    .B1(_04579_),
    .B2(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__inv_2 _19000_ (.A(_04601_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_1 _19001_ (.A(_09232_),
    .B(_04581_),
    .Y(_04602_));
 sky130_fd_sc_hd__a31o_1 _19002_ (.A1(_04542_),
    .A2(net2536),
    .A3(_04580_),
    .B1(_04602_),
    .X(_01508_));
 sky130_fd_sc_hd__nor2_1 _19003_ (.A(_09235_),
    .B(_04581_),
    .Y(_04603_));
 sky130_fd_sc_hd__a31o_1 _19004_ (.A1(_04542_),
    .A2(net2592),
    .A3(_04580_),
    .B1(_04603_),
    .X(_01509_));
 sky130_fd_sc_hd__buf_4 _19005_ (.A(_09226_),
    .X(_04604_));
 sky130_fd_sc_hd__and3_1 _19006_ (.A(_04576_),
    .B(net64),
    .C(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__a31o_1 _19007_ (.A1(_04580_),
    .A2(_04457_),
    .A3(net1729),
    .B1(_04605_),
    .X(_01510_));
 sky130_fd_sc_hd__nand2_1 _19008_ (.A(_04586_),
    .B(net3744),
    .Y(_04606_));
 sky130_fd_sc_hd__a22o_1 _19009_ (.A1(_04585_),
    .A2(_09767_),
    .B1(_04579_),
    .B2(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__inv_2 _19010_ (.A(_04607_),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_1 _19011_ (.A(_03294_),
    .B(_04581_),
    .Y(_04608_));
 sky130_fd_sc_hd__a31o_1 _19012_ (.A1(_04542_),
    .A2(net807),
    .A3(_04581_),
    .B1(_04608_),
    .X(_01416_));
 sky130_fd_sc_hd__and3_1 _19013_ (.A(_04576_),
    .B(net82),
    .C(_04604_),
    .X(_04609_));
 sky130_fd_sc_hd__a31o_1 _19014_ (.A1(_04580_),
    .A2(_04457_),
    .A3(net1121),
    .B1(_04609_),
    .X(_01417_));
 sky130_fd_sc_hd__clkbuf_8 _19015_ (.A(_09164_),
    .X(_04610_));
 sky130_fd_sc_hd__nor2_1 _19016_ (.A(_03482_),
    .B(_04581_),
    .Y(_04611_));
 sky130_fd_sc_hd__a31o_1 _19017_ (.A1(_04610_),
    .A2(net1842),
    .A3(_04581_),
    .B1(_04611_),
    .X(_01418_));
 sky130_fd_sc_hd__nand2_1 _19018_ (.A(_04586_),
    .B(net2853),
    .Y(_04612_));
 sky130_fd_sc_hd__a22o_1 _19019_ (.A1(_04585_),
    .A2(_09255_),
    .B1(_04579_),
    .B2(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__inv_2 _19020_ (.A(_04613_),
    .Y(_01419_));
 sky130_fd_sc_hd__nor2_1 _19021_ (.A(_09259_),
    .B(_04581_),
    .Y(_04614_));
 sky130_fd_sc_hd__a31o_1 _19022_ (.A1(_04610_),
    .A2(net459),
    .A3(_04581_),
    .B1(_04614_),
    .X(_01420_));
 sky130_fd_sc_hd__nand2_1 _19023_ (.A(_04586_),
    .B(net3915),
    .Y(_04615_));
 sky130_fd_sc_hd__a22o_1 _19024_ (.A1(_04585_),
    .A2(net145),
    .B1(_04579_),
    .B2(_04615_),
    .X(_04616_));
 sky130_fd_sc_hd__inv_2 _19025_ (.A(_04616_),
    .Y(_01421_));
 sky130_fd_sc_hd__clkbuf_8 _19026_ (.A(_03834_),
    .X(_04617_));
 sky130_fd_sc_hd__and3_1 _19027_ (.A(_04576_),
    .B(net55),
    .C(_04604_),
    .X(_04618_));
 sky130_fd_sc_hd__a31o_1 _19028_ (.A1(_04580_),
    .A2(_04617_),
    .A3(net783),
    .B1(_04618_),
    .X(_01422_));
 sky130_fd_sc_hd__nand2_1 _19029_ (.A(_04586_),
    .B(net3836),
    .Y(_04619_));
 sky130_fd_sc_hd__a22o_1 _19030_ (.A1(_04585_),
    .A2(net144),
    .B1(_04579_),
    .B2(_04619_),
    .X(_04620_));
 sky130_fd_sc_hd__inv_2 _19031_ (.A(_04620_),
    .Y(_01423_));
 sky130_fd_sc_hd__and3_1 _19032_ (.A(_04576_),
    .B(_03196_),
    .C(_04604_),
    .X(_04621_));
 sky130_fd_sc_hd__a31o_1 _19033_ (.A1(_04580_),
    .A2(_04617_),
    .A3(net1385),
    .B1(_04621_),
    .X(_01328_));
 sky130_fd_sc_hd__nand2_1 _19034_ (.A(_04586_),
    .B(net2919),
    .Y(_04622_));
 sky130_fd_sc_hd__a22o_1 _19035_ (.A1(_04585_),
    .A2(_09365_),
    .B1(_04579_),
    .B2(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__inv_2 _19036_ (.A(_04623_),
    .Y(_01329_));
 sky130_fd_sc_hd__nand2_1 _19037_ (.A(_04586_),
    .B(net3689),
    .Y(_04624_));
 sky130_fd_sc_hd__a22o_1 _19038_ (.A1(_04585_),
    .A2(_10624_),
    .B1(_04579_),
    .B2(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__inv_2 _19039_ (.A(_04625_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _19040_ (.A(_04586_),
    .B(net2916),
    .Y(_04626_));
 sky130_fd_sc_hd__a22o_1 _19041_ (.A1(_04585_),
    .A2(net140),
    .B1(_04579_),
    .B2(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__inv_2 _19042_ (.A(_04627_),
    .Y(_01331_));
 sky130_fd_sc_hd__and3_1 _19043_ (.A(_04576_),
    .B(_03550_),
    .C(_04604_),
    .X(_04628_));
 sky130_fd_sc_hd__a31o_1 _19044_ (.A1(_04580_),
    .A2(_04617_),
    .A3(net1519),
    .B1(_04628_),
    .X(_01332_));
 sky130_fd_sc_hd__clkbuf_8 _19045_ (.A(_08800_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _19046_ (.A(_04629_),
    .B(net3789),
    .Y(_04630_));
 sky130_fd_sc_hd__o2bb2a_1 _19047_ (.A1_N(_04630_),
    .A2_N(_04580_),
    .B1(_09293_),
    .B2(_04577_),
    .X(_01333_));
 sky130_fd_sc_hd__nand2_1 _19048_ (.A(_04629_),
    .B(net3587),
    .Y(_04631_));
 sky130_fd_sc_hd__o2bb2a_1 _19049_ (.A1_N(_04631_),
    .A2_N(_04580_),
    .B1(_09297_),
    .B2(_04577_),
    .X(_01334_));
 sky130_fd_sc_hd__nand2_1 _19050_ (.A(_04629_),
    .B(net3804),
    .Y(_04632_));
 sky130_fd_sc_hd__o2bb2a_1 _19051_ (.A1_N(_04632_),
    .A2_N(_04580_),
    .B1(_09441_),
    .B2(_04577_),
    .X(_01335_));
 sky130_fd_sc_hd__and3_4 _19052_ (.A(_09737_),
    .B(_09444_),
    .C(_09380_),
    .X(_04633_));
 sky130_fd_sc_hd__inv_2 _19053_ (.A(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__nor2_1 _19054_ (.A(_09166_),
    .B(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__clkinv_4 _19055_ (.A(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__buf_4 _19056_ (.A(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__buf_4 _19057_ (.A(_04636_),
    .X(_04638_));
 sky130_fd_sc_hd__nor2_1 _19058_ (.A(_09180_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__a31o_1 _19059_ (.A1(_04610_),
    .A2(net1892),
    .A3(_04637_),
    .B1(_04639_),
    .X(_01240_));
 sky130_fd_sc_hd__nor2_1 _19060_ (.A(_09184_),
    .B(_04638_),
    .Y(_04640_));
 sky130_fd_sc_hd__a31o_1 _19061_ (.A1(_04610_),
    .A2(net1597),
    .A3(_04637_),
    .B1(_04640_),
    .X(_01241_));
 sky130_fd_sc_hd__nor2_1 _19062_ (.A(_03219_),
    .B(_04638_),
    .Y(_04641_));
 sky130_fd_sc_hd__a31o_1 _19063_ (.A1(_04610_),
    .A2(net1325),
    .A3(_04637_),
    .B1(_04641_),
    .X(_01242_));
 sky130_fd_sc_hd__and3_1 _19064_ (.A(_04633_),
    .B(net69),
    .C(_04604_),
    .X(_04642_));
 sky130_fd_sc_hd__a31o_1 _19065_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net1991),
    .B1(_04642_),
    .X(_01243_));
 sky130_fd_sc_hd__nor2_4 _19066_ (.A(_08795_),
    .B(_04634_),
    .Y(_04643_));
 sky130_fd_sc_hd__nand2_1 _19067_ (.A(_04586_),
    .B(net3029),
    .Y(_04644_));
 sky130_fd_sc_hd__a22o_1 _19068_ (.A1(_04643_),
    .A2(_11330_),
    .B1(_04636_),
    .B2(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__inv_2 _19069_ (.A(_04645_),
    .Y(_01244_));
 sky130_fd_sc_hd__and3_1 _19070_ (.A(_04633_),
    .B(net71),
    .C(_04604_),
    .X(_04646_));
 sky130_fd_sc_hd__a31o_1 _19071_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net2572),
    .B1(_04646_),
    .X(_01245_));
 sky130_fd_sc_hd__nand2_1 _19072_ (.A(_04586_),
    .B(net3534),
    .Y(_04647_));
 sky130_fd_sc_hd__a22o_1 _19073_ (.A1(_04643_),
    .A2(_11105_),
    .B1(_04636_),
    .B2(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__inv_2 _19074_ (.A(_04648_),
    .Y(_01246_));
 sky130_fd_sc_hd__and3_1 _19075_ (.A(_04633_),
    .B(net74),
    .C(_04604_),
    .X(_04649_));
 sky130_fd_sc_hd__a31o_1 _19076_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net2640),
    .B1(_04649_),
    .X(_01247_));
 sky130_fd_sc_hd__nor2_1 _19077_ (.A(_03467_),
    .B(_04638_),
    .Y(_04650_));
 sky130_fd_sc_hd__a31o_1 _19078_ (.A1(_04610_),
    .A2(net2278),
    .A3(_04637_),
    .B1(_04650_),
    .X(_01152_));
 sky130_fd_sc_hd__nand2_1 _19079_ (.A(_04586_),
    .B(net3221),
    .Y(_04651_));
 sky130_fd_sc_hd__a22o_1 _19080_ (.A1(_04643_),
    .A2(_09218_),
    .B1(_04636_),
    .B2(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__inv_2 _19081_ (.A(_04652_),
    .Y(_01153_));
 sky130_fd_sc_hd__buf_4 _19082_ (.A(_04184_),
    .X(_04653_));
 sky130_fd_sc_hd__nand2_1 _19083_ (.A(_04653_),
    .B(net3603),
    .Y(_04654_));
 sky130_fd_sc_hd__a22o_1 _19084_ (.A1(_04643_),
    .A2(net143),
    .B1(_04636_),
    .B2(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__inv_2 _19085_ (.A(_04655_),
    .Y(_01154_));
 sky130_fd_sc_hd__nor2_1 _19086_ (.A(_09229_),
    .B(_04638_),
    .Y(_04656_));
 sky130_fd_sc_hd__a31o_1 _19087_ (.A1(_04610_),
    .A2(net2062),
    .A3(_04638_),
    .B1(_04656_),
    .X(_01155_));
 sky130_fd_sc_hd__nor2_1 _19088_ (.A(_09232_),
    .B(_04638_),
    .Y(_04657_));
 sky130_fd_sc_hd__a31o_1 _19089_ (.A1(_04610_),
    .A2(net1205),
    .A3(_04638_),
    .B1(_04657_),
    .X(_01156_));
 sky130_fd_sc_hd__nor2_1 _19090_ (.A(_09235_),
    .B(_04638_),
    .Y(_04658_));
 sky130_fd_sc_hd__a31o_1 _19091_ (.A1(_04610_),
    .A2(net2311),
    .A3(_04638_),
    .B1(_04658_),
    .X(_01157_));
 sky130_fd_sc_hd__and3_1 _19092_ (.A(_04633_),
    .B(net64),
    .C(_04604_),
    .X(_04659_));
 sky130_fd_sc_hd__a31o_1 _19093_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net2446),
    .B1(_04659_),
    .X(_01158_));
 sky130_fd_sc_hd__nand2_1 _19094_ (.A(_04653_),
    .B(net3701),
    .Y(_04660_));
 sky130_fd_sc_hd__a22o_1 _19095_ (.A1(_04643_),
    .A2(_09767_),
    .B1(_04636_),
    .B2(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__inv_2 _19096_ (.A(_04661_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _19097_ (.A(_04653_),
    .B(net3691),
    .Y(_04662_));
 sky130_fd_sc_hd__a22o_1 _19098_ (.A1(_04643_),
    .A2(_09414_),
    .B1(_04636_),
    .B2(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__inv_2 _19099_ (.A(_04663_),
    .Y(_01064_));
 sky130_fd_sc_hd__and3_1 _19100_ (.A(_04633_),
    .B(net82),
    .C(_04604_),
    .X(_04664_));
 sky130_fd_sc_hd__a31o_1 _19101_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net2317),
    .B1(_04664_),
    .X(_01065_));
 sky130_fd_sc_hd__nor2_1 _19102_ (.A(_03482_),
    .B(_04638_),
    .Y(_04665_));
 sky130_fd_sc_hd__a31o_1 _19103_ (.A1(_04610_),
    .A2(net433),
    .A3(_04638_),
    .B1(_04665_),
    .X(_01066_));
 sky130_fd_sc_hd__and3_1 _19104_ (.A(_04633_),
    .B(net52),
    .C(_04604_),
    .X(_04666_));
 sky130_fd_sc_hd__a31o_1 _19105_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net2406),
    .B1(_04666_),
    .X(_01067_));
 sky130_fd_sc_hd__nor2_1 _19106_ (.A(_09259_),
    .B(_04638_),
    .Y(_04667_));
 sky130_fd_sc_hd__a31o_1 _19107_ (.A1(_04610_),
    .A2(net887),
    .A3(_04638_),
    .B1(_04667_),
    .X(_01068_));
 sky130_fd_sc_hd__nand2_1 _19108_ (.A(_04653_),
    .B(net3643),
    .Y(_04668_));
 sky130_fd_sc_hd__a22o_1 _19109_ (.A1(_04643_),
    .A2(_09262_),
    .B1(_04636_),
    .B2(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__inv_2 _19110_ (.A(_04669_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_1 _19111_ (.A(_04653_),
    .B(net2970),
    .Y(_04670_));
 sky130_fd_sc_hd__a22o_1 _19112_ (.A1(_04643_),
    .A2(_09424_),
    .B1(_04636_),
    .B2(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__inv_2 _19113_ (.A(_04671_),
    .Y(_01070_));
 sky130_fd_sc_hd__nand2_1 _19114_ (.A(_04653_),
    .B(net4191),
    .Y(_04672_));
 sky130_fd_sc_hd__a22o_1 _19115_ (.A1(_04643_),
    .A2(_09268_),
    .B1(_04636_),
    .B2(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__inv_2 _19116_ (.A(_04673_),
    .Y(_01071_));
 sky130_fd_sc_hd__and3_1 _19117_ (.A(_04633_),
    .B(net50),
    .C(_04604_),
    .X(_04674_));
 sky130_fd_sc_hd__a31o_1 _19118_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net2481),
    .B1(_04674_),
    .X(_00976_));
 sky130_fd_sc_hd__nor2_1 _19119_ (.A(_03605_),
    .B(_04638_),
    .Y(_04675_));
 sky130_fd_sc_hd__a31o_1 _19120_ (.A1(_04610_),
    .A2(net1922),
    .A3(_04638_),
    .B1(_04675_),
    .X(_00977_));
 sky130_fd_sc_hd__and3_1 _19121_ (.A(_04633_),
    .B(_03199_),
    .C(_04604_),
    .X(_04676_));
 sky130_fd_sc_hd__a31o_1 _19122_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net633),
    .B1(_04676_),
    .X(_00978_));
 sky130_fd_sc_hd__nand2_1 _19123_ (.A(_04653_),
    .B(net3582),
    .Y(_04677_));
 sky130_fd_sc_hd__a22o_1 _19124_ (.A1(_04643_),
    .A2(net140),
    .B1(_04636_),
    .B2(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__inv_2 _19125_ (.A(_04678_),
    .Y(_00979_));
 sky130_fd_sc_hd__and3_1 _19126_ (.A(_04633_),
    .B(_03550_),
    .C(_04604_),
    .X(_04679_));
 sky130_fd_sc_hd__a31o_1 _19127_ (.A1(_04637_),
    .A2(_04617_),
    .A3(net677),
    .B1(_04679_),
    .X(_00980_));
 sky130_fd_sc_hd__nand2_1 _19128_ (.A(_04629_),
    .B(net3007),
    .Y(_04680_));
 sky130_fd_sc_hd__o2bb2a_1 _19129_ (.A1_N(_04680_),
    .A2_N(_04637_),
    .B1(_09293_),
    .B2(_04634_),
    .X(_00981_));
 sky130_fd_sc_hd__nand2_1 _19130_ (.A(_04629_),
    .B(net3239),
    .Y(_04681_));
 sky130_fd_sc_hd__o2bb2a_1 _19131_ (.A1_N(_04681_),
    .A2_N(_04637_),
    .B1(_09297_),
    .B2(_04634_),
    .X(_00982_));
 sky130_fd_sc_hd__nand2_1 _19132_ (.A(_04629_),
    .B(net3391),
    .Y(_04682_));
 sky130_fd_sc_hd__o2bb2a_1 _19133_ (.A1_N(_04682_),
    .A2_N(_04637_),
    .B1(_09441_),
    .B2(_04634_),
    .X(_00983_));
 sky130_fd_sc_hd__nor2_4 _19134_ (.A(_08736_),
    .B(_09925_),
    .Y(_04683_));
 sky130_fd_sc_hd__inv_2 _19135_ (.A(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__nor2_1 _19136_ (.A(_08728_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__inv_2 _19137_ (.A(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__buf_4 _19138_ (.A(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__nor2_1 _19139_ (.A(_09180_),
    .B(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__a31o_1 _19140_ (.A1(_04610_),
    .A2(net757),
    .A3(_04687_),
    .B1(_04688_),
    .X(_00880_));
 sky130_fd_sc_hd__nor2_1 _19141_ (.A(_08797_),
    .B(_04684_),
    .Y(_04689_));
 sky130_fd_sc_hd__buf_4 _19142_ (.A(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__buf_4 _19143_ (.A(_04686_),
    .X(_04691_));
 sky130_fd_sc_hd__nand2_1 _19144_ (.A(_04653_),
    .B(net2980),
    .Y(_04692_));
 sky130_fd_sc_hd__a22o_1 _19145_ (.A1(_04690_),
    .A2(_09314_),
    .B1(_04691_),
    .B2(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__inv_2 _19146_ (.A(_04693_),
    .Y(_00881_));
 sky130_fd_sc_hd__nand2_1 _19147_ (.A(_04653_),
    .B(net3057),
    .Y(_04694_));
 sky130_fd_sc_hd__a22o_1 _19148_ (.A1(_04690_),
    .A2(_09459_),
    .B1(_04691_),
    .B2(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__inv_2 _19149_ (.A(_04695_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _19150_ (.A(_04653_),
    .B(net3334),
    .Y(_04696_));
 sky130_fd_sc_hd__a22o_1 _19151_ (.A1(_04690_),
    .A2(_10983_),
    .B1(_04691_),
    .B2(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__inv_2 _19152_ (.A(_04697_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand2_1 _19153_ (.A(_04653_),
    .B(net3459),
    .Y(_04698_));
 sky130_fd_sc_hd__a22o_1 _19154_ (.A1(_04690_),
    .A2(_11330_),
    .B1(_04691_),
    .B2(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__inv_2 _19155_ (.A(_04699_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _19156_ (.A(_04653_),
    .B(net3299),
    .Y(_04700_));
 sky130_fd_sc_hd__a22o_1 _19157_ (.A1(_04690_),
    .A2(_09204_),
    .B1(_04691_),
    .B2(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__inv_2 _19158_ (.A(_04701_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _19159_ (.A(_04653_),
    .B(net3267),
    .Y(_04702_));
 sky130_fd_sc_hd__a22o_1 _19160_ (.A1(_04690_),
    .A2(_11105_),
    .B1(_04691_),
    .B2(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__inv_2 _19161_ (.A(_04703_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand2_1 _19162_ (.A(_04653_),
    .B(net3314),
    .Y(_04704_));
 sky130_fd_sc_hd__a22o_1 _19163_ (.A1(_04690_),
    .A2(_09211_),
    .B1(_04691_),
    .B2(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__inv_2 _19164_ (.A(_04705_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_1 _19165_ (.A(_03467_),
    .B(_04691_),
    .Y(_04706_));
 sky130_fd_sc_hd__a31o_1 _19166_ (.A1(_04610_),
    .A2(net1631),
    .A3(_04687_),
    .B1(_04706_),
    .X(_00792_));
 sky130_fd_sc_hd__nand2_1 _19167_ (.A(_04653_),
    .B(net3493),
    .Y(_04707_));
 sky130_fd_sc_hd__a22o_1 _19168_ (.A1(_04690_),
    .A2(_09218_),
    .B1(_04691_),
    .B2(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__inv_2 _19169_ (.A(_04708_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_1 _19170_ (.A(_04653_),
    .B(net3511),
    .Y(_04709_));
 sky130_fd_sc_hd__a22o_1 _19171_ (.A1(_04690_),
    .A2(net143),
    .B1(_04691_),
    .B2(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__inv_2 _19172_ (.A(_04710_),
    .Y(_00794_));
 sky130_fd_sc_hd__nor2_1 _19173_ (.A(_09229_),
    .B(_04691_),
    .Y(_04711_));
 sky130_fd_sc_hd__a31o_1 _19174_ (.A1(_04610_),
    .A2(net1257),
    .A3(_04687_),
    .B1(_04711_),
    .X(_00795_));
 sky130_fd_sc_hd__nor2_1 _19175_ (.A(_09232_),
    .B(_04691_),
    .Y(_04712_));
 sky130_fd_sc_hd__a31o_1 _19176_ (.A1(_04610_),
    .A2(net1049),
    .A3(_04687_),
    .B1(_04712_),
    .X(_00796_));
 sky130_fd_sc_hd__buf_6 _19177_ (.A(_09164_),
    .X(_04713_));
 sky130_fd_sc_hd__nor2_1 _19178_ (.A(_09235_),
    .B(_04691_),
    .Y(_04714_));
 sky130_fd_sc_hd__a31o_1 _19179_ (.A1(_04713_),
    .A2(net2152),
    .A3(_04687_),
    .B1(_04714_),
    .X(_00797_));
 sky130_fd_sc_hd__and3_1 _19180_ (.A(_04683_),
    .B(net64),
    .C(_04604_),
    .X(_04715_));
 sky130_fd_sc_hd__a31o_1 _19181_ (.A1(_04687_),
    .A2(_04617_),
    .A3(net1979),
    .B1(_04715_),
    .X(_00798_));
 sky130_fd_sc_hd__nor2_1 _19182_ (.A(_09242_),
    .B(_04691_),
    .Y(_04716_));
 sky130_fd_sc_hd__a31o_1 _19183_ (.A1(_04713_),
    .A2(net1265),
    .A3(_04687_),
    .B1(_04716_),
    .X(_00799_));
 sky130_fd_sc_hd__nor2_1 _19184_ (.A(_03294_),
    .B(_04691_),
    .Y(_04717_));
 sky130_fd_sc_hd__a31o_1 _19185_ (.A1(_04713_),
    .A2(net1747),
    .A3(_04687_),
    .B1(_04717_),
    .X(_00704_));
 sky130_fd_sc_hd__clkbuf_8 _19186_ (.A(_10310_),
    .X(_04718_));
 sky130_fd_sc_hd__nand2_1 _19187_ (.A(_04718_),
    .B(net3248),
    .Y(_04719_));
 sky130_fd_sc_hd__a22o_1 _19188_ (.A1(_04690_),
    .A2(_09248_),
    .B1(_04686_),
    .B2(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__inv_2 _19189_ (.A(_04720_),
    .Y(_00705_));
 sky130_fd_sc_hd__nand2_1 _19190_ (.A(_04718_),
    .B(net3530),
    .Y(_04721_));
 sky130_fd_sc_hd__a22o_1 _19191_ (.A1(_04690_),
    .A2(_09347_),
    .B1(_04686_),
    .B2(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__inv_2 _19192_ (.A(_04722_),
    .Y(_00706_));
 sky130_fd_sc_hd__and3_1 _19193_ (.A(_04683_),
    .B(net52),
    .C(_04604_),
    .X(_04723_));
 sky130_fd_sc_hd__a31o_1 _19194_ (.A1(_04687_),
    .A2(_04617_),
    .A3(net1879),
    .B1(_04723_),
    .X(_00707_));
 sky130_fd_sc_hd__nand2_1 _19195_ (.A(_04718_),
    .B(net3509),
    .Y(_04724_));
 sky130_fd_sc_hd__a22o_1 _19196_ (.A1(_04690_),
    .A2(_11136_),
    .B1(_04686_),
    .B2(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__inv_2 _19197_ (.A(_04725_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _19198_ (.A(_04718_),
    .B(net3446),
    .Y(_04726_));
 sky130_fd_sc_hd__a22o_1 _19199_ (.A1(_04690_),
    .A2(_09262_),
    .B1(_04686_),
    .B2(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__inv_2 _19200_ (.A(_04727_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _19201_ (.A(_04718_),
    .B(net2953),
    .Y(_04728_));
 sky130_fd_sc_hd__a22o_1 _19202_ (.A1(_04690_),
    .A2(_09424_),
    .B1(_04686_),
    .B2(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__inv_2 _19203_ (.A(_04729_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand2_1 _19204_ (.A(_04718_),
    .B(net3636),
    .Y(_04730_));
 sky130_fd_sc_hd__a22o_1 _19205_ (.A1(_04690_),
    .A2(_09268_),
    .B1(_04686_),
    .B2(_04730_),
    .X(_04731_));
 sky130_fd_sc_hd__inv_2 _19206_ (.A(_04731_),
    .Y(_00711_));
 sky130_fd_sc_hd__clkbuf_8 _19207_ (.A(_09226_),
    .X(_04732_));
 sky130_fd_sc_hd__and3_1 _19208_ (.A(_04683_),
    .B(net50),
    .C(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a31o_1 _19209_ (.A1(_04687_),
    .A2(_04617_),
    .A3(net2137),
    .B1(_04733_),
    .X(_00616_));
 sky130_fd_sc_hd__nor2_1 _19210_ (.A(_03605_),
    .B(_04691_),
    .Y(_04734_));
 sky130_fd_sc_hd__a31o_1 _19211_ (.A1(_04713_),
    .A2(net1489),
    .A3(_04687_),
    .B1(_04734_),
    .X(_00617_));
 sky130_fd_sc_hd__nand2_1 _19212_ (.A(_04718_),
    .B(net3064),
    .Y(_04735_));
 sky130_fd_sc_hd__a22o_1 _19213_ (.A1(_04690_),
    .A2(_10624_),
    .B1(_04686_),
    .B2(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__inv_2 _19214_ (.A(_04736_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand2_1 _19215_ (.A(_04718_),
    .B(net3591),
    .Y(_04737_));
 sky130_fd_sc_hd__a22o_1 _19216_ (.A1(_04689_),
    .A2(net140),
    .B1(_04686_),
    .B2(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__inv_2 _19217_ (.A(net3592),
    .Y(_00619_));
 sky130_fd_sc_hd__and3_1 _19218_ (.A(_04683_),
    .B(_03550_),
    .C(_04732_),
    .X(_04739_));
 sky130_fd_sc_hd__a31o_1 _19219_ (.A1(_04687_),
    .A2(_04617_),
    .A3(net2518),
    .B1(_04739_),
    .X(_00620_));
 sky130_fd_sc_hd__clkbuf_8 _19220_ (.A(_03834_),
    .X(_04740_));
 sky130_fd_sc_hd__and3_1 _19221_ (.A(_04683_),
    .B(net78),
    .C(_04732_),
    .X(_04741_));
 sky130_fd_sc_hd__a31o_1 _19222_ (.A1(_04687_),
    .A2(_04740_),
    .A3(net2500),
    .B1(_04741_),
    .X(_00621_));
 sky130_fd_sc_hd__nand2_1 _19223_ (.A(_04629_),
    .B(net3514),
    .Y(_04742_));
 sky130_fd_sc_hd__o2bb2a_1 _19224_ (.A1_N(_04742_),
    .A2_N(_04687_),
    .B1(_09297_),
    .B2(_04684_),
    .X(_00622_));
 sky130_fd_sc_hd__nand2_1 _19225_ (.A(_04629_),
    .B(net3960),
    .Y(_04743_));
 sky130_fd_sc_hd__o2bb2a_1 _19226_ (.A1_N(_04743_),
    .A2_N(_04687_),
    .B1(_09441_),
    .B2(_04684_),
    .X(_00623_));
 sky130_fd_sc_hd__nor2_4 _19227_ (.A(_08736_),
    .B(_09984_),
    .Y(_04744_));
 sky130_fd_sc_hd__inv_2 _19228_ (.A(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__nor2_4 _19229_ (.A(_09190_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__nor2_1 _19230_ (.A(_09304_),
    .B(_04745_),
    .Y(_04747_));
 sky130_fd_sc_hd__clkinv_4 _19231_ (.A(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__clkbuf_8 _19232_ (.A(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__nand2_1 _19233_ (.A(_04718_),
    .B(net4202),
    .Y(_04750_));
 sky130_fd_sc_hd__a22o_1 _19234_ (.A1(_04746_),
    .A2(_10239_),
    .B1(_04749_),
    .B2(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__inv_2 _19235_ (.A(_04751_),
    .Y(_00528_));
 sky130_fd_sc_hd__clkbuf_8 _19236_ (.A(_04748_),
    .X(_04752_));
 sky130_fd_sc_hd__nor2_1 _19237_ (.A(_09184_),
    .B(_04749_),
    .Y(_04753_));
 sky130_fd_sc_hd__a31o_1 _19238_ (.A1(_04713_),
    .A2(net2212),
    .A3(_04752_),
    .B1(_04753_),
    .X(_00529_));
 sky130_fd_sc_hd__nor2_1 _19239_ (.A(_09187_),
    .B(_04749_),
    .Y(_04754_));
 sky130_fd_sc_hd__a31o_1 _19240_ (.A1(_04713_),
    .A2(net2344),
    .A3(_04752_),
    .B1(_04754_),
    .X(_00530_));
 sky130_fd_sc_hd__and3_1 _19241_ (.A(_04744_),
    .B(net69),
    .C(_04732_),
    .X(_04755_));
 sky130_fd_sc_hd__a31o_1 _19242_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net2565),
    .B1(_04755_),
    .X(_00531_));
 sky130_fd_sc_hd__and3_1 _19243_ (.A(_04744_),
    .B(_10586_),
    .C(_04732_),
    .X(_04756_));
 sky130_fd_sc_hd__a31o_1 _19244_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net2583),
    .B1(_04756_),
    .X(_00532_));
 sky130_fd_sc_hd__and3_1 _19245_ (.A(_04744_),
    .B(net71),
    .C(_04732_),
    .X(_04757_));
 sky130_fd_sc_hd__a31o_1 _19246_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net2282),
    .B1(_04757_),
    .X(_00533_));
 sky130_fd_sc_hd__nand2_1 _19247_ (.A(_04718_),
    .B(net4249),
    .Y(_04758_));
 sky130_fd_sc_hd__a22o_1 _19248_ (.A1(_04746_),
    .A2(_09397_),
    .B1(_04749_),
    .B2(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__inv_2 _19249_ (.A(_04759_),
    .Y(_00534_));
 sky130_fd_sc_hd__and3_1 _19250_ (.A(_04744_),
    .B(net74),
    .C(_04732_),
    .X(_04760_));
 sky130_fd_sc_hd__a31o_1 _19251_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net2623),
    .B1(_04760_),
    .X(_00535_));
 sky130_fd_sc_hd__nor2_1 _19252_ (.A(_03467_),
    .B(_04749_),
    .Y(_04761_));
 sky130_fd_sc_hd__a31o_1 _19253_ (.A1(_04713_),
    .A2(net2395),
    .A3(_04752_),
    .B1(_04761_),
    .X(_00440_));
 sky130_fd_sc_hd__nand2_1 _19254_ (.A(_04718_),
    .B(net3354),
    .Y(_04762_));
 sky130_fd_sc_hd__a22o_1 _19255_ (.A1(_04746_),
    .A2(net146),
    .B1(_04749_),
    .B2(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__inv_2 _19256_ (.A(_04763_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _19257_ (.A(_04718_),
    .B(net3298),
    .Y(_04764_));
 sky130_fd_sc_hd__a22o_1 _19258_ (.A1(_04746_),
    .A2(net143),
    .B1(_04748_),
    .B2(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__inv_2 _19259_ (.A(_04765_),
    .Y(_00442_));
 sky130_fd_sc_hd__nor2_1 _19260_ (.A(_09229_),
    .B(_04749_),
    .Y(_04766_));
 sky130_fd_sc_hd__a31o_1 _19261_ (.A1(_04713_),
    .A2(net2193),
    .A3(_04752_),
    .B1(_04766_),
    .X(_00443_));
 sky130_fd_sc_hd__nand2_1 _19262_ (.A(_04718_),
    .B(net3768),
    .Y(_04767_));
 sky130_fd_sc_hd__a22o_1 _19263_ (.A1(_04746_),
    .A2(_09592_),
    .B1(_04748_),
    .B2(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__inv_2 _19264_ (.A(_04768_),
    .Y(_00444_));
 sky130_fd_sc_hd__nor2_1 _19265_ (.A(_09235_),
    .B(_04749_),
    .Y(_04769_));
 sky130_fd_sc_hd__a31o_1 _19266_ (.A1(_04713_),
    .A2(net1864),
    .A3(_04752_),
    .B1(_04769_),
    .X(_00445_));
 sky130_fd_sc_hd__nand2_1 _19267_ (.A(_04718_),
    .B(net3145),
    .Y(_04770_));
 sky130_fd_sc_hd__a22o_1 _19268_ (.A1(_04746_),
    .A2(_09238_),
    .B1(_04748_),
    .B2(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__inv_2 _19269_ (.A(_04771_),
    .Y(_00446_));
 sky130_fd_sc_hd__nor2_1 _19270_ (.A(_09242_),
    .B(_04749_),
    .Y(_04772_));
 sky130_fd_sc_hd__a31o_1 _19271_ (.A1(_04713_),
    .A2(net1537),
    .A3(_04749_),
    .B1(_04772_),
    .X(_00447_));
 sky130_fd_sc_hd__nor2_1 _19272_ (.A(_03294_),
    .B(_04749_),
    .Y(_04773_));
 sky130_fd_sc_hd__a31o_1 _19273_ (.A1(_04713_),
    .A2(net1832),
    .A3(_04749_),
    .B1(_04773_),
    .X(_00352_));
 sky130_fd_sc_hd__and3_1 _19274_ (.A(_04744_),
    .B(net82),
    .C(_04732_),
    .X(_04774_));
 sky130_fd_sc_hd__a31o_1 _19275_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net2281),
    .B1(_04774_),
    .X(_00353_));
 sky130_fd_sc_hd__nand2_1 _19276_ (.A(_04718_),
    .B(net3842),
    .Y(_04775_));
 sky130_fd_sc_hd__a22o_1 _19277_ (.A1(_04746_),
    .A2(_09347_),
    .B1(_04748_),
    .B2(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__inv_2 _19278_ (.A(_04776_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _19279_ (.A(_04718_),
    .B(net3490),
    .Y(_04777_));
 sky130_fd_sc_hd__a22o_1 _19280_ (.A1(_04746_),
    .A2(_09255_),
    .B1(_04748_),
    .B2(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__inv_2 _19281_ (.A(_04778_),
    .Y(_00355_));
 sky130_fd_sc_hd__nor2_1 _19282_ (.A(_09259_),
    .B(_04749_),
    .Y(_04779_));
 sky130_fd_sc_hd__a31o_1 _19283_ (.A1(_04713_),
    .A2(net1487),
    .A3(_04749_),
    .B1(_04779_),
    .X(_00356_));
 sky130_fd_sc_hd__buf_4 _19284_ (.A(_10310_),
    .X(_04780_));
 sky130_fd_sc_hd__nand2_1 _19285_ (.A(_04780_),
    .B(net3801),
    .Y(_04781_));
 sky130_fd_sc_hd__a22o_1 _19286_ (.A1(_04746_),
    .A2(_09262_),
    .B1(_04748_),
    .B2(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__inv_2 _19287_ (.A(_04782_),
    .Y(_00357_));
 sky130_fd_sc_hd__and3_1 _19288_ (.A(_04744_),
    .B(net55),
    .C(_04732_),
    .X(_04783_));
 sky130_fd_sc_hd__a31o_1 _19289_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net1784),
    .B1(_04783_),
    .X(_00358_));
 sky130_fd_sc_hd__nand2_1 _19290_ (.A(_04780_),
    .B(net3563),
    .Y(_04784_));
 sky130_fd_sc_hd__a22o_1 _19291_ (.A1(_04746_),
    .A2(_09268_),
    .B1(_04748_),
    .B2(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__inv_2 _19292_ (.A(_04785_),
    .Y(_00359_));
 sky130_fd_sc_hd__and3_1 _19293_ (.A(_04744_),
    .B(net50),
    .C(_04732_),
    .X(_04786_));
 sky130_fd_sc_hd__a31o_1 _19294_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net1587),
    .B1(_04786_),
    .X(_00264_));
 sky130_fd_sc_hd__nand2_1 _19295_ (.A(_04780_),
    .B(net2773),
    .Y(_04787_));
 sky130_fd_sc_hd__a22o_1 _19296_ (.A1(_04746_),
    .A2(_09365_),
    .B1(_04748_),
    .B2(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__inv_2 _19297_ (.A(_04788_),
    .Y(_00265_));
 sky130_fd_sc_hd__and3_1 _19298_ (.A(_04744_),
    .B(_03199_),
    .C(_04732_),
    .X(_04789_));
 sky130_fd_sc_hd__a31o_1 _19299_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net1219),
    .B1(_04789_),
    .X(_00266_));
 sky130_fd_sc_hd__nand2_1 _19300_ (.A(_04780_),
    .B(net2833),
    .Y(_04790_));
 sky130_fd_sc_hd__a22o_1 _19301_ (.A1(_04746_),
    .A2(net140),
    .B1(_04748_),
    .B2(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__inv_2 _19302_ (.A(_04791_),
    .Y(_00267_));
 sky130_fd_sc_hd__and3_1 _19303_ (.A(_04744_),
    .B(net77),
    .C(_04732_),
    .X(_04792_));
 sky130_fd_sc_hd__a31o_1 _19304_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net617),
    .B1(_04792_),
    .X(_00268_));
 sky130_fd_sc_hd__and3_1 _19305_ (.A(_04744_),
    .B(net78),
    .C(_04732_),
    .X(_04793_));
 sky130_fd_sc_hd__a31o_1 _19306_ (.A1(_04752_),
    .A2(_04740_),
    .A3(net835),
    .B1(_04793_),
    .X(_00269_));
 sky130_fd_sc_hd__nand2_1 _19307_ (.A(_04629_),
    .B(net3233),
    .Y(_04794_));
 sky130_fd_sc_hd__o2bb2a_1 _19308_ (.A1_N(_04794_),
    .A2_N(_04752_),
    .B1(_09297_),
    .B2(_04745_),
    .X(_00270_));
 sky130_fd_sc_hd__nor2_1 _19309_ (.A(_09299_),
    .B(_04749_),
    .Y(_04795_));
 sky130_fd_sc_hd__a31o_1 _19310_ (.A1(_04713_),
    .A2(net517),
    .A3(_04749_),
    .B1(_04795_),
    .X(_00271_));
 sky130_fd_sc_hd__nor2_4 _19311_ (.A(_08736_),
    .B(_10041_),
    .Y(_04796_));
 sky130_fd_sc_hd__inv_2 _19312_ (.A(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__nor2_1 _19313_ (.A(_09625_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__inv_2 _19314_ (.A(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__buf_4 _19315_ (.A(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__buf_4 _19316_ (.A(_04799_),
    .X(_04801_));
 sky130_fd_sc_hd__nor2_1 _19317_ (.A(_09180_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__a31o_1 _19318_ (.A1(_04713_),
    .A2(net863),
    .A3(_04800_),
    .B1(_04802_),
    .X(_00176_));
 sky130_fd_sc_hd__nor2_1 _19319_ (.A(_09184_),
    .B(_04801_),
    .Y(_04803_));
 sky130_fd_sc_hd__a31o_1 _19320_ (.A1(_04713_),
    .A2(net1609),
    .A3(_04800_),
    .B1(_04803_),
    .X(_00177_));
 sky130_fd_sc_hd__nor2_1 _19321_ (.A(_09187_),
    .B(_04801_),
    .Y(_04804_));
 sky130_fd_sc_hd__a31o_1 _19322_ (.A1(_04713_),
    .A2(net1544),
    .A3(_04800_),
    .B1(_04804_),
    .X(_00178_));
 sky130_fd_sc_hd__and3_1 _19323_ (.A(_04796_),
    .B(net69),
    .C(_04732_),
    .X(_04805_));
 sky130_fd_sc_hd__a31o_1 _19324_ (.A1(_04800_),
    .A2(_04740_),
    .A3(net2293),
    .B1(_04805_),
    .X(_00179_));
 sky130_fd_sc_hd__and3_1 _19325_ (.A(_04796_),
    .B(_10586_),
    .C(_04732_),
    .X(_04806_));
 sky130_fd_sc_hd__a31o_1 _19326_ (.A1(_04800_),
    .A2(_04740_),
    .A3(net1731),
    .B1(_04806_),
    .X(_00180_));
 sky130_fd_sc_hd__nor2_4 _19327_ (.A(_08797_),
    .B(_04797_),
    .Y(_04807_));
 sky130_fd_sc_hd__nand2_1 _19328_ (.A(_04780_),
    .B(net3351),
    .Y(_04808_));
 sky130_fd_sc_hd__a22o_1 _19329_ (.A1(_04807_),
    .A2(_09204_),
    .B1(_04801_),
    .B2(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__inv_2 _19330_ (.A(_04809_),
    .Y(_00181_));
 sky130_fd_sc_hd__nor2_1 _19331_ (.A(_09208_),
    .B(_04801_),
    .Y(_04810_));
 sky130_fd_sc_hd__a31o_1 _19332_ (.A1(_09224_),
    .A2(net1187),
    .A3(_04800_),
    .B1(_04810_),
    .X(_00182_));
 sky130_fd_sc_hd__nand2_1 _19333_ (.A(_04780_),
    .B(net3160),
    .Y(_04811_));
 sky130_fd_sc_hd__a22o_1 _19334_ (.A1(_04807_),
    .A2(_09211_),
    .B1(_04801_),
    .B2(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__inv_2 _19335_ (.A(_04812_),
    .Y(_00183_));
 sky130_fd_sc_hd__nor2_1 _19336_ (.A(_03467_),
    .B(_04801_),
    .Y(_04813_));
 sky130_fd_sc_hd__a31o_1 _19337_ (.A1(_09224_),
    .A2(net1107),
    .A3(_04800_),
    .B1(_04813_),
    .X(_00088_));
 sky130_fd_sc_hd__nand2_1 _19338_ (.A(_04780_),
    .B(net2989),
    .Y(_04814_));
 sky130_fd_sc_hd__a22o_1 _19339_ (.A1(_04807_),
    .A2(net146),
    .B1(_04801_),
    .B2(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__inv_2 _19340_ (.A(_04815_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_1 _19341_ (.A(_04780_),
    .B(net2938),
    .Y(_04816_));
 sky130_fd_sc_hd__a22o_1 _19342_ (.A1(_04807_),
    .A2(net143),
    .B1(_04801_),
    .B2(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__inv_2 _19343_ (.A(_04817_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_1 _19344_ (.A(_04780_),
    .B(net3330),
    .Y(_04818_));
 sky130_fd_sc_hd__a22o_1 _19345_ (.A1(_04807_),
    .A2(_09588_),
    .B1(_04801_),
    .B2(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__inv_2 _19346_ (.A(_04819_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor2_1 _19347_ (.A(_09232_),
    .B(_04801_),
    .Y(_04820_));
 sky130_fd_sc_hd__a31o_1 _19348_ (.A1(_09224_),
    .A2(net639),
    .A3(_04800_),
    .B1(_04820_),
    .X(_00092_));
 sky130_fd_sc_hd__nand2_1 _19349_ (.A(_04780_),
    .B(net3017),
    .Y(_04821_));
 sky130_fd_sc_hd__a22o_1 _19350_ (.A1(_04807_),
    .A2(_09337_),
    .B1(_04801_),
    .B2(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__inv_2 _19351_ (.A(_04822_),
    .Y(_00093_));
 sky130_fd_sc_hd__and3_1 _19352_ (.A(_04796_),
    .B(net64),
    .C(_04732_),
    .X(_04823_));
 sky130_fd_sc_hd__a31o_1 _19353_ (.A1(_04800_),
    .A2(_04740_),
    .A3(net1871),
    .B1(_04823_),
    .X(_00094_));
 sky130_fd_sc_hd__nand2_1 _19354_ (.A(_04780_),
    .B(net3844),
    .Y(_04824_));
 sky130_fd_sc_hd__a22o_1 _19355_ (.A1(_04807_),
    .A2(_09767_),
    .B1(_04799_),
    .B2(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__inv_2 _19356_ (.A(_04825_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_1 _19357_ (.A(_04780_),
    .B(net3460),
    .Y(_04826_));
 sky130_fd_sc_hd__a22o_1 _19358_ (.A1(_04807_),
    .A2(_09414_),
    .B1(_04799_),
    .B2(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__inv_2 _19359_ (.A(_04827_),
    .Y(_02552_));
 sky130_fd_sc_hd__buf_4 _19360_ (.A(_09226_),
    .X(_04828_));
 sky130_fd_sc_hd__and3_1 _19361_ (.A(_04796_),
    .B(net82),
    .C(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__a31o_1 _19362_ (.A1(_04800_),
    .A2(_04740_),
    .A3(net1872),
    .B1(_04829_),
    .X(_02553_));
 sky130_fd_sc_hd__nor2_1 _19363_ (.A(_09252_),
    .B(_04801_),
    .Y(_04830_));
 sky130_fd_sc_hd__a31o_1 _19364_ (.A1(_09224_),
    .A2(net957),
    .A3(_04800_),
    .B1(_04830_),
    .X(_02554_));
 sky130_fd_sc_hd__nand2_1 _19365_ (.A(_04780_),
    .B(net3265),
    .Y(_04831_));
 sky130_fd_sc_hd__a22o_1 _19366_ (.A1(_04807_),
    .A2(_09255_),
    .B1(_04799_),
    .B2(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__inv_2 _19367_ (.A(_04832_),
    .Y(_02555_));
 sky130_fd_sc_hd__nand2_1 _19368_ (.A(_04780_),
    .B(net2926),
    .Y(_04833_));
 sky130_fd_sc_hd__a22o_1 _19369_ (.A1(_04807_),
    .A2(_11136_),
    .B1(_04799_),
    .B2(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__inv_2 _19370_ (.A(_04834_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _19371_ (.A(_04780_),
    .B(net3146),
    .Y(_04835_));
 sky130_fd_sc_hd__a22o_1 _19372_ (.A1(_04807_),
    .A2(_09262_),
    .B1(_04799_),
    .B2(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__inv_2 _19373_ (.A(_04836_),
    .Y(_02557_));
 sky130_fd_sc_hd__and3_1 _19374_ (.A(_04796_),
    .B(net55),
    .C(_04828_),
    .X(_04837_));
 sky130_fd_sc_hd__a31o_1 _19375_ (.A1(_04800_),
    .A2(_04740_),
    .A3(net1067),
    .B1(_04837_),
    .X(_02558_));
 sky130_fd_sc_hd__nand2_1 _19376_ (.A(_04780_),
    .B(net3491),
    .Y(_04838_));
 sky130_fd_sc_hd__a22o_1 _19377_ (.A1(_04807_),
    .A2(_09268_),
    .B1(_04799_),
    .B2(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__inv_2 _19378_ (.A(_04839_),
    .Y(_02559_));
 sky130_fd_sc_hd__buf_4 _19379_ (.A(_10310_),
    .X(_04840_));
 sky130_fd_sc_hd__nand2_1 _19380_ (.A(_04840_),
    .B(net2996),
    .Y(_04841_));
 sky130_fd_sc_hd__a22o_1 _19381_ (.A1(_04807_),
    .A2(_09494_),
    .B1(_04799_),
    .B2(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__inv_2 _19382_ (.A(_04842_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor2_1 _19383_ (.A(_09276_),
    .B(_04801_),
    .Y(_04843_));
 sky130_fd_sc_hd__a31o_1 _19384_ (.A1(_09224_),
    .A2(net1957),
    .A3(_04800_),
    .B1(_04843_),
    .X(_02465_));
 sky130_fd_sc_hd__and3_1 _19385_ (.A(_04796_),
    .B(_03199_),
    .C(_04828_),
    .X(_04844_));
 sky130_fd_sc_hd__a31o_1 _19386_ (.A1(_04800_),
    .A2(_08801_),
    .A3(net2628),
    .B1(_04844_),
    .X(_02466_));
 sky130_fd_sc_hd__nand2_1 _19387_ (.A(_04840_),
    .B(net3895),
    .Y(_04845_));
 sky130_fd_sc_hd__a22o_1 _19388_ (.A1(_04807_),
    .A2(net140),
    .B1(_04799_),
    .B2(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__inv_2 _19389_ (.A(_04846_),
    .Y(_02467_));
 sky130_fd_sc_hd__nand2_1 _19390_ (.A(_04840_),
    .B(net3929),
    .Y(_04847_));
 sky130_fd_sc_hd__a22o_1 _19391_ (.A1(_04807_),
    .A2(_09287_),
    .B1(_04799_),
    .B2(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__inv_2 _19392_ (.A(_04848_),
    .Y(_02468_));
 sky130_fd_sc_hd__nand2_1 _19393_ (.A(_04629_),
    .B(net4105),
    .Y(_04849_));
 sky130_fd_sc_hd__o2bb2a_1 _19394_ (.A1_N(_04849_),
    .A2_N(_04800_),
    .B1(_09293_),
    .B2(_04797_),
    .X(_02469_));
 sky130_fd_sc_hd__nand2_1 _19395_ (.A(_04629_),
    .B(net4017),
    .Y(_04850_));
 sky130_fd_sc_hd__o2bb2a_1 _19396_ (.A1_N(_04850_),
    .A2_N(_04800_),
    .B1(_09297_),
    .B2(_04797_),
    .X(_02470_));
 sky130_fd_sc_hd__nor2_1 _19397_ (.A(_09299_),
    .B(_04801_),
    .Y(_04851_));
 sky130_fd_sc_hd__a31o_1 _19398_ (.A1(_09224_),
    .A2(net1676),
    .A3(_04801_),
    .B1(_04851_),
    .X(_02471_));
 sky130_fd_sc_hd__nor2_1 _19399_ (.A(_08736_),
    .B(_10096_),
    .Y(_04852_));
 sky130_fd_sc_hd__inv_2 _19400_ (.A(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__nor2_4 _19401_ (.A(_08794_),
    .B(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__clkbuf_8 _19402_ (.A(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__nor2_1 _19403_ (.A(_09166_),
    .B(_04853_),
    .Y(_04856_));
 sky130_fd_sc_hd__inv_2 _19404_ (.A(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__buf_4 _19405_ (.A(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__nand2_1 _19406_ (.A(_04840_),
    .B(net2932),
    .Y(_04859_));
 sky130_fd_sc_hd__a22o_1 _19407_ (.A1(_04855_),
    .A2(_10239_),
    .B1(_04858_),
    .B2(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__inv_2 _19408_ (.A(_04860_),
    .Y(_02376_));
 sky130_fd_sc_hd__nand2_1 _19409_ (.A(_04840_),
    .B(net2910),
    .Y(_04861_));
 sky130_fd_sc_hd__a22o_1 _19410_ (.A1(_04855_),
    .A2(_09314_),
    .B1(_04858_),
    .B2(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__inv_2 _19411_ (.A(_04862_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_1 _19412_ (.A(_04840_),
    .B(net3909),
    .Y(_04863_));
 sky130_fd_sc_hd__a22o_1 _19413_ (.A1(_04855_),
    .A2(_09459_),
    .B1(_04858_),
    .B2(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__inv_2 _19414_ (.A(_04864_),
    .Y(_02378_));
 sky130_fd_sc_hd__nand2_1 _19415_ (.A(_04840_),
    .B(net3863),
    .Y(_04865_));
 sky130_fd_sc_hd__a22o_1 _19416_ (.A1(_04855_),
    .A2(_10983_),
    .B1(_04858_),
    .B2(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__inv_2 _19417_ (.A(_04866_),
    .Y(_02379_));
 sky130_fd_sc_hd__nand2_1 _19418_ (.A(_04840_),
    .B(net3865),
    .Y(_04867_));
 sky130_fd_sc_hd__a22o_1 _19419_ (.A1(_04855_),
    .A2(_09200_),
    .B1(_04858_),
    .B2(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__inv_2 _19420_ (.A(_04868_),
    .Y(_02380_));
 sky130_fd_sc_hd__nand2_1 _19421_ (.A(_04840_),
    .B(net3002),
    .Y(_04869_));
 sky130_fd_sc_hd__a22o_1 _19422_ (.A1(_04855_),
    .A2(_09204_),
    .B1(_04858_),
    .B2(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__inv_2 _19423_ (.A(_04870_),
    .Y(_02381_));
 sky130_fd_sc_hd__nand2_1 _19424_ (.A(_04840_),
    .B(net3826),
    .Y(_04871_));
 sky130_fd_sc_hd__a22o_1 _19425_ (.A1(_04855_),
    .A2(_09397_),
    .B1(_04858_),
    .B2(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__inv_2 _19426_ (.A(_04872_),
    .Y(_02382_));
 sky130_fd_sc_hd__nand2_1 _19427_ (.A(_04840_),
    .B(net3204),
    .Y(_04873_));
 sky130_fd_sc_hd__a22o_1 _19428_ (.A1(_04855_),
    .A2(_09211_),
    .B1(_04858_),
    .B2(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__inv_2 _19429_ (.A(_04874_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _19430_ (.A(_04840_),
    .B(net3986),
    .Y(_04875_));
 sky130_fd_sc_hd__a22o_1 _19431_ (.A1(_04855_),
    .A2(_09530_),
    .B1(_04858_),
    .B2(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__inv_2 _19432_ (.A(_04876_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2_1 _19433_ (.A(_04840_),
    .B(net3638),
    .Y(_04877_));
 sky130_fd_sc_hd__a22o_1 _19434_ (.A1(_04855_),
    .A2(net146),
    .B1(_04858_),
    .B2(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__inv_2 _19435_ (.A(_04878_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _19436_ (.A(_04840_),
    .B(net3846),
    .Y(_04879_));
 sky130_fd_sc_hd__a22o_1 _19437_ (.A1(_04855_),
    .A2(net143),
    .B1(_04858_),
    .B2(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__inv_2 _19438_ (.A(_04880_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _19439_ (.A(_04840_),
    .B(net3607),
    .Y(_04881_));
 sky130_fd_sc_hd__a22o_1 _19440_ (.A1(_04855_),
    .A2(_09588_),
    .B1(_04858_),
    .B2(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__inv_2 _19441_ (.A(_04882_),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_1 _19442_ (.A(_04840_),
    .B(net3340),
    .Y(_04883_));
 sky130_fd_sc_hd__a22o_1 _19443_ (.A1(_04855_),
    .A2(_09592_),
    .B1(_04858_),
    .B2(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__inv_2 _19444_ (.A(_04884_),
    .Y(_02292_));
 sky130_fd_sc_hd__buf_4 _19445_ (.A(_04857_),
    .X(_04885_));
 sky130_fd_sc_hd__buf_4 _19446_ (.A(_10310_),
    .X(_04886_));
 sky130_fd_sc_hd__nand2_1 _19447_ (.A(_04886_),
    .B(net3119),
    .Y(_04887_));
 sky130_fd_sc_hd__a22o_1 _19448_ (.A1(_04855_),
    .A2(_09337_),
    .B1(_04885_),
    .B2(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__inv_2 _19449_ (.A(_04888_),
    .Y(_02293_));
 sky130_fd_sc_hd__nand2_1 _19450_ (.A(_04886_),
    .B(net2995),
    .Y(_04889_));
 sky130_fd_sc_hd__a22o_1 _19451_ (.A1(_04855_),
    .A2(_09238_),
    .B1(_04885_),
    .B2(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__inv_2 _19452_ (.A(_04890_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_1 _19453_ (.A(_04886_),
    .B(net2873),
    .Y(_04891_));
 sky130_fd_sc_hd__a22o_1 _19454_ (.A1(_04855_),
    .A2(_09767_),
    .B1(_04885_),
    .B2(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__inv_2 _19455_ (.A(_04892_),
    .Y(_02295_));
 sky130_fd_sc_hd__nand2_1 _19456_ (.A(_04886_),
    .B(net3268),
    .Y(_04893_));
 sky130_fd_sc_hd__a22o_1 _19457_ (.A1(_04854_),
    .A2(_09414_),
    .B1(_04885_),
    .B2(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__inv_2 _19458_ (.A(_04894_),
    .Y(_02200_));
 sky130_fd_sc_hd__nand2_1 _19459_ (.A(_04886_),
    .B(net3035),
    .Y(_04895_));
 sky130_fd_sc_hd__a22o_1 _19460_ (.A1(_04854_),
    .A2(_09248_),
    .B1(_04885_),
    .B2(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__inv_2 _19461_ (.A(_04896_),
    .Y(_02201_));
 sky130_fd_sc_hd__nand2_1 _19462_ (.A(_04886_),
    .B(net3237),
    .Y(_04897_));
 sky130_fd_sc_hd__a22o_1 _19463_ (.A1(_04854_),
    .A2(_09347_),
    .B1(_04885_),
    .B2(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__inv_2 _19464_ (.A(_04898_),
    .Y(_02202_));
 sky130_fd_sc_hd__nand2_1 _19465_ (.A(_04886_),
    .B(net3308),
    .Y(_04899_));
 sky130_fd_sc_hd__a22o_1 _19466_ (.A1(_04854_),
    .A2(_09255_),
    .B1(_04885_),
    .B2(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__inv_2 _19467_ (.A(_04900_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2_1 _19468_ (.A(_04886_),
    .B(net3255),
    .Y(_04901_));
 sky130_fd_sc_hd__a22o_1 _19469_ (.A1(_04854_),
    .A2(_11136_),
    .B1(_04885_),
    .B2(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__inv_2 _19470_ (.A(_04902_),
    .Y(_02204_));
 sky130_fd_sc_hd__nand2_1 _19471_ (.A(_04886_),
    .B(net3544),
    .Y(_04903_));
 sky130_fd_sc_hd__a22o_1 _19472_ (.A1(_04854_),
    .A2(net145),
    .B1(_04885_),
    .B2(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__inv_2 _19473_ (.A(_04904_),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _19474_ (.A(_04886_),
    .B(net3167),
    .Y(_04905_));
 sky130_fd_sc_hd__a22o_1 _19475_ (.A1(_04854_),
    .A2(_09424_),
    .B1(_04885_),
    .B2(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__inv_2 _19476_ (.A(_04906_),
    .Y(_02206_));
 sky130_fd_sc_hd__nand2_1 _19477_ (.A(_04886_),
    .B(net2867),
    .Y(_04907_));
 sky130_fd_sc_hd__a22o_1 _19478_ (.A1(_04854_),
    .A2(net144),
    .B1(_04885_),
    .B2(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__inv_2 _19479_ (.A(_04908_),
    .Y(_02207_));
 sky130_fd_sc_hd__nand2_1 _19480_ (.A(_04886_),
    .B(net3163),
    .Y(_04909_));
 sky130_fd_sc_hd__a22o_1 _19481_ (.A1(_04854_),
    .A2(_09494_),
    .B1(_04885_),
    .B2(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__inv_2 _19482_ (.A(_04910_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _19483_ (.A(_04886_),
    .B(net3075),
    .Y(_04911_));
 sky130_fd_sc_hd__a22o_1 _19484_ (.A1(_04854_),
    .A2(_09365_),
    .B1(_04885_),
    .B2(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__inv_2 _19485_ (.A(_04912_),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_1 _19486_ (.A(_04886_),
    .B(net3155),
    .Y(_04913_));
 sky130_fd_sc_hd__a22o_1 _19487_ (.A1(_04854_),
    .A2(_10624_),
    .B1(_04885_),
    .B2(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__inv_2 _19488_ (.A(_04914_),
    .Y(_02114_));
 sky130_fd_sc_hd__nand2_1 _19489_ (.A(_04886_),
    .B(net3317),
    .Y(_04915_));
 sky130_fd_sc_hd__a22o_1 _19490_ (.A1(_04854_),
    .A2(net140),
    .B1(_04885_),
    .B2(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__inv_2 _19491_ (.A(_04916_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _19492_ (.A(_04886_),
    .B(net3348),
    .Y(_04917_));
 sky130_fd_sc_hd__a22o_1 _19493_ (.A1(_04854_),
    .A2(_09287_),
    .B1(_04885_),
    .B2(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__inv_2 _19494_ (.A(_04918_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2_1 _19495_ (.A(_04629_),
    .B(net3489),
    .Y(_04919_));
 sky130_fd_sc_hd__o2bb2a_1 _19496_ (.A1_N(_04919_),
    .A2_N(_04858_),
    .B1(_09293_),
    .B2(_04853_),
    .X(_02117_));
 sky130_fd_sc_hd__nand2_1 _19497_ (.A(_04629_),
    .B(net3684),
    .Y(_04920_));
 sky130_fd_sc_hd__o2bb2a_1 _19498_ (.A1_N(_04920_),
    .A2_N(_04858_),
    .B1(_09297_),
    .B2(_04853_),
    .X(_02118_));
 sky130_fd_sc_hd__nand2_1 _19499_ (.A(_04629_),
    .B(net3629),
    .Y(_04921_));
 sky130_fd_sc_hd__o2bb2a_1 _19500_ (.A1_N(_04921_),
    .A2_N(_04858_),
    .B1(_09441_),
    .B2(_04853_),
    .X(_02119_));
 sky130_fd_sc_hd__nor2_4 _19501_ (.A(_08736_),
    .B(_10173_),
    .Y(_04922_));
 sky130_fd_sc_hd__inv_2 _19502_ (.A(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__nor2_4 _19503_ (.A(_08795_),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__nor2_1 _19504_ (.A(_09625_),
    .B(_04923_),
    .Y(_04925_));
 sky130_fd_sc_hd__inv_2 _19505_ (.A(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__buf_4 _19506_ (.A(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__nand2_1 _19507_ (.A(_08777_),
    .B(net2798),
    .Y(_04928_));
 sky130_fd_sc_hd__a22o_1 _19508_ (.A1(_04924_),
    .A2(_10239_),
    .B1(_04927_),
    .B2(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__inv_2 _19509_ (.A(_04929_),
    .Y(_02024_));
 sky130_fd_sc_hd__buf_4 _19510_ (.A(_04926_),
    .X(_04930_));
 sky130_fd_sc_hd__nor2_1 _19511_ (.A(_09184_),
    .B(_04927_),
    .Y(_04931_));
 sky130_fd_sc_hd__a31o_1 _19512_ (.A1(_09224_),
    .A2(net765),
    .A3(_04930_),
    .B1(_04931_),
    .X(_02025_));
 sky130_fd_sc_hd__nor2_1 _19513_ (.A(_09187_),
    .B(_04927_),
    .Y(_04932_));
 sky130_fd_sc_hd__a31o_1 _19514_ (.A1(_09224_),
    .A2(net491),
    .A3(_04930_),
    .B1(_04932_),
    .X(_02026_));
 sky130_fd_sc_hd__and3_1 _19515_ (.A(_04922_),
    .B(net69),
    .C(_04828_),
    .X(_04933_));
 sky130_fd_sc_hd__a31o_1 _19516_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net929),
    .B1(_04933_),
    .X(_02027_));
 sky130_fd_sc_hd__and3_1 _19517_ (.A(_04922_),
    .B(_10586_),
    .C(_04828_),
    .X(_04934_));
 sky130_fd_sc_hd__a31o_1 _19518_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net1665),
    .B1(_04934_),
    .X(_02028_));
 sky130_fd_sc_hd__and3_1 _19519_ (.A(_04922_),
    .B(net71),
    .C(_04828_),
    .X(_04935_));
 sky130_fd_sc_hd__a31o_1 _19520_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net849),
    .B1(_04935_),
    .X(_02029_));
 sky130_fd_sc_hd__nor2_1 _19521_ (.A(_09208_),
    .B(_04927_),
    .Y(_04936_));
 sky130_fd_sc_hd__a31o_1 _19522_ (.A1(_09224_),
    .A2(net531),
    .A3(_04927_),
    .B1(_04936_),
    .X(_02030_));
 sky130_fd_sc_hd__and3_1 _19523_ (.A(_04922_),
    .B(net74),
    .C(_04828_),
    .X(_04937_));
 sky130_fd_sc_hd__a31o_1 _19524_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net623),
    .B1(_04937_),
    .X(_02031_));
 sky130_fd_sc_hd__nor2_1 _19525_ (.A(_03467_),
    .B(_04927_),
    .Y(_04938_));
 sky130_fd_sc_hd__a31o_1 _19526_ (.A1(_09224_),
    .A2(net443),
    .A3(_04927_),
    .B1(_04938_),
    .X(_01776_));
 sky130_fd_sc_hd__nand2_1 _19527_ (.A(_08777_),
    .B(net2820),
    .Y(_04939_));
 sky130_fd_sc_hd__a22o_1 _19528_ (.A1(_04924_),
    .A2(net146),
    .B1(_04927_),
    .B2(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__inv_2 _19529_ (.A(_04940_),
    .Y(_01777_));
 sky130_fd_sc_hd__nand2_1 _19530_ (.A(_08777_),
    .B(net2829),
    .Y(_04941_));
 sky130_fd_sc_hd__a22o_1 _19531_ (.A1(_04924_),
    .A2(net143),
    .B1(_04926_),
    .B2(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__inv_2 _19532_ (.A(_04942_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _19533_ (.A(_09229_),
    .B(_04927_),
    .Y(_04943_));
 sky130_fd_sc_hd__a31o_1 _19534_ (.A1(_09224_),
    .A2(net505),
    .A3(_04927_),
    .B1(_04943_),
    .X(_01779_));
 sky130_fd_sc_hd__nand2_1 _19535_ (.A(_08777_),
    .B(net2789),
    .Y(_04944_));
 sky130_fd_sc_hd__a22o_1 _19536_ (.A1(_04924_),
    .A2(_09592_),
    .B1(_04926_),
    .B2(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__inv_2 _19537_ (.A(_04945_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _19538_ (.A(_08777_),
    .B(net2929),
    .Y(_04946_));
 sky130_fd_sc_hd__a22o_1 _19539_ (.A1(_04924_),
    .A2(_09337_),
    .B1(_04926_),
    .B2(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__inv_2 _19540_ (.A(_04947_),
    .Y(_01781_));
 sky130_fd_sc_hd__and3_1 _19541_ (.A(_04922_),
    .B(net64),
    .C(_04828_),
    .X(_04948_));
 sky130_fd_sc_hd__a31o_1 _19542_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net2595),
    .B1(_04948_),
    .X(_01782_));
 sky130_fd_sc_hd__nor2_1 _19543_ (.A(_09242_),
    .B(_04927_),
    .Y(_04949_));
 sky130_fd_sc_hd__a31o_1 _19544_ (.A1(_09224_),
    .A2(net809),
    .A3(_04927_),
    .B1(_04949_),
    .X(_01783_));
 sky130_fd_sc_hd__nand2_1 _19545_ (.A(_08777_),
    .B(net2917),
    .Y(_04950_));
 sky130_fd_sc_hd__a22o_1 _19546_ (.A1(_04924_),
    .A2(_09414_),
    .B1(_04926_),
    .B2(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__inv_2 _19547_ (.A(_04951_),
    .Y(_00888_));
 sky130_fd_sc_hd__and3_1 _19548_ (.A(_04922_),
    .B(net82),
    .C(_04828_),
    .X(_04952_));
 sky130_fd_sc_hd__a31o_1 _19549_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net647),
    .B1(_04952_),
    .X(_00889_));
 sky130_fd_sc_hd__nor2_1 _19550_ (.A(_09252_),
    .B(_04927_),
    .Y(_04953_));
 sky130_fd_sc_hd__a31o_1 _19551_ (.A1(_09224_),
    .A2(net471),
    .A3(_04927_),
    .B1(_04953_),
    .X(_00890_));
 sky130_fd_sc_hd__and3_1 _19552_ (.A(_04922_),
    .B(net52),
    .C(_04828_),
    .X(_04954_));
 sky130_fd_sc_hd__a31o_1 _19553_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net1359),
    .B1(_04954_),
    .X(_00891_));
 sky130_fd_sc_hd__nand2_1 _19554_ (.A(_08777_),
    .B(net3143),
    .Y(_04955_));
 sky130_fd_sc_hd__a22o_1 _19555_ (.A1(_04924_),
    .A2(_09353_),
    .B1(_04926_),
    .B2(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__inv_2 _19556_ (.A(_04956_),
    .Y(_00892_));
 sky130_fd_sc_hd__nand2_1 _19557_ (.A(_08777_),
    .B(net3140),
    .Y(_04957_));
 sky130_fd_sc_hd__a22o_1 _19558_ (.A1(_04924_),
    .A2(net145),
    .B1(_04926_),
    .B2(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__inv_2 _19559_ (.A(_04958_),
    .Y(_00893_));
 sky130_fd_sc_hd__nand2_1 _19560_ (.A(_08777_),
    .B(net2900),
    .Y(_04959_));
 sky130_fd_sc_hd__a22o_1 _19561_ (.A1(_04924_),
    .A2(_09424_),
    .B1(_04926_),
    .B2(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__inv_2 _19562_ (.A(_04960_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_1 _19563_ (.A(_08777_),
    .B(net2828),
    .Y(_04961_));
 sky130_fd_sc_hd__a22o_1 _19564_ (.A1(_04924_),
    .A2(net144),
    .B1(_04926_),
    .B2(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__inv_2 _19565_ (.A(_04962_),
    .Y(_00895_));
 sky130_fd_sc_hd__and3_1 _19566_ (.A(_04922_),
    .B(net50),
    .C(_04828_),
    .X(_04963_));
 sky130_fd_sc_hd__a31o_1 _19567_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net607),
    .B1(_04963_),
    .X(_00000_));
 sky130_fd_sc_hd__nor2_1 _19568_ (.A(_09276_),
    .B(_04927_),
    .Y(_04964_));
 sky130_fd_sc_hd__a31o_1 _19569_ (.A1(_09224_),
    .A2(net2705),
    .A3(_04927_),
    .B1(_04964_),
    .X(_00001_));
 sky130_fd_sc_hd__and3_1 _19570_ (.A(_04922_),
    .B(_03199_),
    .C(_04828_),
    .X(_04965_));
 sky130_fd_sc_hd__a31o_1 _19571_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net1745),
    .B1(_04965_),
    .X(_00002_));
 sky130_fd_sc_hd__and3_1 _19572_ (.A(_04922_),
    .B(net76),
    .C(_04828_),
    .X(_04966_));
 sky130_fd_sc_hd__a31o_1 _19573_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net2547),
    .B1(_04966_),
    .X(_00003_));
 sky130_fd_sc_hd__and3_1 _19574_ (.A(_04922_),
    .B(net77),
    .C(_04828_),
    .X(_04967_));
 sky130_fd_sc_hd__a31o_1 _19575_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net695),
    .B1(_04967_),
    .X(_00004_));
 sky130_fd_sc_hd__and3_1 _19576_ (.A(_04922_),
    .B(net78),
    .C(_04828_),
    .X(_04968_));
 sky130_fd_sc_hd__a31o_1 _19577_ (.A1(_04930_),
    .A2(_08801_),
    .A3(net2378),
    .B1(_04968_),
    .X(_00005_));
 sky130_fd_sc_hd__nand2_1 _19578_ (.A(_04629_),
    .B(net4302),
    .Y(_04969_));
 sky130_fd_sc_hd__o2bb2a_1 _19579_ (.A1_N(_04969_),
    .A2_N(_04930_),
    .B1(_09297_),
    .B2(_04923_),
    .X(_00006_));
 sky130_fd_sc_hd__nand2_1 _19580_ (.A(_04629_),
    .B(net4295),
    .Y(_04970_));
 sky130_fd_sc_hd__o2bb2a_1 _19581_ (.A1_N(_04970_),
    .A2_N(_04930_),
    .B1(_09441_),
    .B2(_04923_),
    .X(_00007_));
 sky130_fd_sc_hd__buf_6 _19582_ (.A(_08792_),
    .X(_04971_));
 sky130_fd_sc_hd__or2_1 _19583_ (.A(net3436),
    .B(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__inv_2 _19584_ (.A(_04972_),
    .Y(_02560_));
 sky130_fd_sc_hd__nand2_1 _19585_ (.A(net3436),
    .B(net4294),
    .Y(_04973_));
 sky130_fd_sc_hd__inv_2 _19586_ (.A(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__nor2_1 _19587_ (.A(net3436),
    .B(net4294),
    .Y(_04975_));
 sky130_fd_sc_hd__or3_1 _19588_ (.A(_04974_),
    .B(_04975_),
    .C(_04971_),
    .X(_04976_));
 sky130_fd_sc_hd__inv_2 _19589_ (.A(_04976_),
    .Y(_02561_));
 sky130_fd_sc_hd__and3_1 _19590_ (.A(net3436),
    .B(net4294),
    .C(net4322),
    .X(_04977_));
 sky130_fd_sc_hd__nor2_1 _19591_ (.A(net4322),
    .B(_04974_),
    .Y(_04978_));
 sky130_fd_sc_hd__or3_1 _19592_ (.A(_04977_),
    .B(_04978_),
    .C(_04971_),
    .X(_04979_));
 sky130_fd_sc_hd__inv_2 _19593_ (.A(_04979_),
    .Y(_02562_));
 sky130_fd_sc_hd__and3_1 _19594_ (.A(_04974_),
    .B(net4322),
    .C(net4314),
    .X(_04980_));
 sky130_fd_sc_hd__or2_1 _19595_ (.A(net4314),
    .B(_04977_),
    .X(_04981_));
 sky130_fd_sc_hd__or3b_1 _19596_ (.A(_04980_),
    .B(_04971_),
    .C_N(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__inv_2 _19597_ (.A(_04982_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_1 _19598_ (.A(net4276),
    .B(_04980_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_1 _19599_ (.A(_04980_),
    .B(net4276),
    .Y(_04984_));
 sky130_fd_sc_hd__or3b_1 _19600_ (.A(_08723_),
    .B(net4277),
    .C_N(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__inv_2 _19601_ (.A(net4278),
    .Y(_02564_));
 sky130_fd_sc_hd__inv_2 _19602_ (.A(net2905),
    .Y(_04986_));
 sky130_fd_sc_hd__or2_1 _19603_ (.A(_04986_),
    .B(_04984_),
    .X(_04987_));
 sky130_fd_sc_hd__nand2_1 _19604_ (.A(_04984_),
    .B(_04986_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand3_1 _19605_ (.A(_04987_),
    .B(_09165_),
    .C(net2906),
    .Y(_04989_));
 sky130_fd_sc_hd__inv_2 _19606_ (.A(net2907),
    .Y(_02565_));
 sky130_fd_sc_hd__inv_2 _19607_ (.A(net4324),
    .Y(_04990_));
 sky130_fd_sc_hd__and2_1 _19608_ (.A(_04987_),
    .B(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__or2_1 _19609_ (.A(_04990_),
    .B(_04987_),
    .X(_04992_));
 sky130_fd_sc_hd__inv_2 _19610_ (.A(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__or3_1 _19611_ (.A(_08723_),
    .B(_04991_),
    .C(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__inv_2 _19612_ (.A(_04994_),
    .Y(_02566_));
 sky130_fd_sc_hd__or2_1 _19613_ (.A(net2762),
    .B(_04993_),
    .X(_04995_));
 sky130_fd_sc_hd__nand2_1 _19614_ (.A(_04993_),
    .B(net2762),
    .Y(_04996_));
 sky130_fd_sc_hd__nand3_1 _19615_ (.A(net2763),
    .B(_09165_),
    .C(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__inv_2 _19616_ (.A(net2764),
    .Y(_02567_));
 sky130_fd_sc_hd__or2_1 _19617_ (.A(net2695),
    .B(_04996_),
    .X(_04998_));
 sky130_fd_sc_hd__nand2_1 _19618_ (.A(_04996_),
    .B(net2695),
    .Y(_04999_));
 sky130_fd_sc_hd__a21oi_1 _19619_ (.A1(net2696),
    .A2(_04999_),
    .B1(_08723_),
    .Y(_02568_));
 sky130_fd_sc_hd__nor2_2 _19620_ (.A(\res_h_counter[0] ),
    .B(\res_h_counter[1] ),
    .Y(_05000_));
 sky130_fd_sc_hd__nor2_2 _19621_ (.A(\res_h_counter[2] ),
    .B(\res_h_counter[3] ),
    .Y(_05001_));
 sky130_fd_sc_hd__and2_2 _19622_ (.A(_05000_),
    .B(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__inv_2 _19623_ (.A(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__nor2_8 _19624_ (.A(\res_h_counter[4] ),
    .B(_08713_),
    .Y(_05004_));
 sky130_fd_sc_hd__and3_4 _19625_ (.A(_05004_),
    .B(_08709_),
    .C(_08662_),
    .X(_05005_));
 sky130_fd_sc_hd__buf_4 _19626_ (.A(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__inv_2 _19627_ (.A(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__nor2_1 _19628_ (.A(_05003_),
    .B(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__clkbuf_8 _19629_ (.A(_08676_),
    .X(_05009_));
 sky130_fd_sc_hd__buf_6 _19630_ (.A(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__nand2_2 _19631_ (.A(_05008_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__nor2_2 _19632_ (.A(net3038),
    .B(_08696_),
    .Y(_05012_));
 sky130_fd_sc_hd__nand2_2 _19633_ (.A(_05012_),
    .B(_05001_),
    .Y(_05013_));
 sky130_fd_sc_hd__nor2_1 _19634_ (.A(_05013_),
    .B(_05007_),
    .Y(_05014_));
 sky130_fd_sc_hd__nand2_2 _19635_ (.A(_05014_),
    .B(_05010_),
    .Y(_05015_));
 sky130_fd_sc_hd__nand2_1 _19636_ (.A(_05011_),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__nor2b_4 _19637_ (.A(net2770),
    .B_N(net3038),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_4 _19638_ (.A(_05017_),
    .B(_05001_),
    .Y(_05018_));
 sky130_fd_sc_hd__nor2_1 _19639_ (.A(_05018_),
    .B(_05007_),
    .Y(_05019_));
 sky130_fd_sc_hd__buf_6 _19640_ (.A(_05009_),
    .X(_05020_));
 sky130_fd_sc_hd__clkbuf_8 _19641_ (.A(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__nand2_2 _19642_ (.A(_05019_),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand2_4 _19643_ (.A(net2770),
    .B(net3038),
    .Y(_05023_));
 sky130_fd_sc_hd__clkinv_4 _19644_ (.A(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_4 _19645_ (.A(_05024_),
    .B(_05001_),
    .Y(_05025_));
 sky130_fd_sc_hd__nor2_1 _19646_ (.A(_05025_),
    .B(_05007_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_2 _19647_ (.A(_05026_),
    .B(_05010_),
    .Y(_05027_));
 sky130_fd_sc_hd__nand2_1 _19648_ (.A(_05022_),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__inv_2 _19649_ (.A(net3919),
    .Y(_05029_));
 sky130_fd_sc_hd__nor2_2 _19650_ (.A(\res_h_counter[3] ),
    .B(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__and2_4 _19651_ (.A(_05012_),
    .B(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__inv_2 _19652_ (.A(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__nor2_1 _19653_ (.A(_05032_),
    .B(_05007_),
    .Y(_05033_));
 sky130_fd_sc_hd__buf_4 _19654_ (.A(_05010_),
    .X(_05034_));
 sky130_fd_sc_hd__nand2_1 _19655_ (.A(_05033_),
    .B(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__and2_4 _19656_ (.A(_05030_),
    .B(_05000_),
    .X(_05036_));
 sky130_fd_sc_hd__inv_2 _19657_ (.A(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nor2_1 _19658_ (.A(_05037_),
    .B(_05007_),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _19659_ (.A(_05038_),
    .B(_05034_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_1 _19660_ (.A(_05035_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__and2_1 _19661_ (.A(_05017_),
    .B(_05030_),
    .X(_05041_));
 sky130_fd_sc_hd__buf_8 _19662_ (.A(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__and3_4 _19663_ (.A(_05006_),
    .B(_05020_),
    .C(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__nand2_4 _19664_ (.A(_05030_),
    .B(_05024_),
    .Y(_05044_));
 sky130_fd_sc_hd__inv_2 _19665_ (.A(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__and3_4 _19666_ (.A(_05006_),
    .B(_05045_),
    .C(_05020_),
    .X(_05046_));
 sky130_fd_sc_hd__or2_1 _19667_ (.A(_05043_),
    .B(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__or4_1 _19668_ (.A(_05016_),
    .B(_05028_),
    .C(_05040_),
    .D(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_2 _19669_ (.A(\res_h_counter[2] ),
    .B(net2785),
    .Y(_05049_));
 sky130_fd_sc_hd__inv_2 _19670_ (.A(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__nand2_4 _19671_ (.A(_05050_),
    .B(_05000_),
    .Y(_05051_));
 sky130_fd_sc_hd__clkinv_4 _19672_ (.A(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__and3_2 _19673_ (.A(_05006_),
    .B(_05052_),
    .C(_05009_),
    .X(_05053_));
 sky130_fd_sc_hd__and2_4 _19674_ (.A(_05012_),
    .B(_05050_),
    .X(_05054_));
 sky130_fd_sc_hd__and3_1 _19675_ (.A(_05006_),
    .B(_05009_),
    .C(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_4 _19676_ (.A(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__nand2_4 _19677_ (.A(_05017_),
    .B(_05050_),
    .Y(_05057_));
 sky130_fd_sc_hd__nor2_2 _19678_ (.A(_05057_),
    .B(_05007_),
    .Y(_05058_));
 sky130_fd_sc_hd__buf_6 _19679_ (.A(_05010_),
    .X(_05059_));
 sky130_fd_sc_hd__nand2_1 _19680_ (.A(_05058_),
    .B(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__nor2_8 _19681_ (.A(_05023_),
    .B(_05049_),
    .Y(_05061_));
 sky130_fd_sc_hd__inv_4 _19682_ (.A(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__nor2_2 _19683_ (.A(_05062_),
    .B(_05007_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _19684_ (.A(_05063_),
    .B(_05059_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand2_1 _19685_ (.A(_05060_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__nor2_4 _19686_ (.A(\res_h_counter[2] ),
    .B(_08705_),
    .Y(_05066_));
 sky130_fd_sc_hd__nand2_2 _19687_ (.A(_05066_),
    .B(_05000_),
    .Y(_05067_));
 sky130_fd_sc_hd__inv_6 _19688_ (.A(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__and3_4 _19689_ (.A(_05006_),
    .B(_05009_),
    .C(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__nand2_8 _19690_ (.A(_05066_),
    .B(_05024_),
    .Y(_05070_));
 sky130_fd_sc_hd__inv_2 _19691_ (.A(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__and3_1 _19692_ (.A(_05006_),
    .B(_05071_),
    .C(_08676_),
    .X(_05072_));
 sky130_fd_sc_hd__clkbuf_4 _19693_ (.A(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__nand2_4 _19694_ (.A(_05012_),
    .B(_05066_),
    .Y(_05074_));
 sky130_fd_sc_hd__inv_2 _19695_ (.A(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__and3_4 _19696_ (.A(_05006_),
    .B(_05009_),
    .C(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__nand2_4 _19697_ (.A(_05017_),
    .B(_05066_),
    .Y(_05077_));
 sky130_fd_sc_hd__inv_2 _19698_ (.A(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__and3_4 _19699_ (.A(_05006_),
    .B(_05009_),
    .C(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__or4_1 _19700_ (.A(_05069_),
    .B(_05073_),
    .C(_05076_),
    .D(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__or4_1 _19701_ (.A(_05053_),
    .B(_05056_),
    .C(_05065_),
    .D(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__nor2_1 _19702_ (.A(_05048_),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__nor2_8 _19703_ (.A(\res_h_counter[4] ),
    .B(\res_h_counter[5] ),
    .Y(_05083_));
 sky130_fd_sc_hd__and3_1 _19704_ (.A(_05083_),
    .B(_08709_),
    .C(_08662_),
    .X(_05084_));
 sky130_fd_sc_hd__clkbuf_8 _19705_ (.A(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__nand2_1 _19706_ (.A(_05085_),
    .B(_05021_),
    .Y(_05086_));
 sky130_fd_sc_hd__nand2_4 _19707_ (.A(\res_h_counter[4] ),
    .B(\res_h_counter[5] ),
    .Y(_05087_));
 sky130_fd_sc_hd__clkinv_4 _19708_ (.A(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__and3_1 _19709_ (.A(_05088_),
    .B(_08709_),
    .C(_08662_),
    .X(_05089_));
 sky130_fd_sc_hd__clkbuf_4 _19710_ (.A(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__buf_4 _19711_ (.A(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__and3_1 _19712_ (.A(_05091_),
    .B(_05009_),
    .C(_05031_),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_4 _19713_ (.A(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__inv_2 _19714_ (.A(_05090_),
    .Y(_05094_));
 sky130_fd_sc_hd__nor2_2 _19715_ (.A(_05044_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _19716_ (.A(_05095_),
    .B(_05010_),
    .Y(_05096_));
 sky130_fd_sc_hd__inv_2 _19717_ (.A(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__and3_4 _19718_ (.A(_05091_),
    .B(_05036_),
    .C(_05020_),
    .X(_05098_));
 sky130_fd_sc_hd__buf_12 _19719_ (.A(_08677_),
    .X(_05099_));
 sky130_fd_sc_hd__buf_8 _19720_ (.A(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__inv_2 _19721_ (.A(_05042_),
    .Y(_05101_));
 sky130_fd_sc_hd__or3_1 _19722_ (.A(_05100_),
    .B(_05101_),
    .C(_05094_),
    .X(_05102_));
 sky130_fd_sc_hd__inv_2 _19723_ (.A(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__or4_1 _19724_ (.A(_05093_),
    .B(_05097_),
    .C(_05098_),
    .D(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__and3_1 _19725_ (.A(_05091_),
    .B(_05009_),
    .C(_05054_),
    .X(_05105_));
 sky130_fd_sc_hd__buf_2 _19726_ (.A(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__and3_1 _19727_ (.A(_05091_),
    .B(_05009_),
    .C(_05052_),
    .X(_05107_));
 sky130_fd_sc_hd__clkbuf_4 _19728_ (.A(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__nor2_2 _19729_ (.A(_05057_),
    .B(_05094_),
    .Y(_05109_));
 sky130_fd_sc_hd__nand2_1 _19730_ (.A(_05109_),
    .B(_05059_),
    .Y(_05110_));
 sky130_fd_sc_hd__nor2_2 _19731_ (.A(_05062_),
    .B(_05094_),
    .Y(_05111_));
 sky130_fd_sc_hd__clkbuf_4 _19732_ (.A(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__buf_8 _19733_ (.A(_05059_),
    .X(_05113_));
 sky130_fd_sc_hd__nand2_1 _19734_ (.A(_05112_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__nand2_1 _19735_ (.A(_05110_),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__nor3_1 _19736_ (.A(_05106_),
    .B(_05108_),
    .C(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__nor2_2 _19737_ (.A(_05070_),
    .B(_05094_),
    .Y(_05117_));
 sky130_fd_sc_hd__and3_1 _19738_ (.A(_05091_),
    .B(_05068_),
    .C(_05009_),
    .X(_05118_));
 sky130_fd_sc_hd__clkbuf_4 _19739_ (.A(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__and3_1 _19740_ (.A(_05091_),
    .B(_05009_),
    .C(_05075_),
    .X(_05120_));
 sky130_fd_sc_hd__clkbuf_4 _19741_ (.A(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__and3_1 _19742_ (.A(_05091_),
    .B(_05020_),
    .C(_05078_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_4 _19743_ (.A(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__a2111oi_1 _19744_ (.A1(_05113_),
    .A2(_05117_),
    .B1(_05119_),
    .C1(_05121_),
    .D1(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__inv_6 _19745_ (.A(_05013_),
    .Y(_05125_));
 sky130_fd_sc_hd__and3_1 _19746_ (.A(_05091_),
    .B(_05009_),
    .C(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__buf_2 _19747_ (.A(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__and3_1 _19748_ (.A(_05091_),
    .B(_05002_),
    .C(_05009_),
    .X(_05128_));
 sky130_fd_sc_hd__buf_2 _19749_ (.A(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__inv_4 _19750_ (.A(_05018_),
    .Y(_05130_));
 sky130_fd_sc_hd__and3_1 _19751_ (.A(_05091_),
    .B(_05020_),
    .C(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__clkbuf_4 _19752_ (.A(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__inv_2 _19753_ (.A(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__clkinv_4 _19754_ (.A(_05025_),
    .Y(_05134_));
 sky130_fd_sc_hd__and3_1 _19755_ (.A(_05091_),
    .B(_05020_),
    .C(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__clkbuf_4 _19756_ (.A(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__inv_2 _19757_ (.A(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand2_1 _19758_ (.A(_05133_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__nor3_1 _19759_ (.A(_05127_),
    .B(_05129_),
    .C(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__and4b_1 _19760_ (.A_N(_05104_),
    .B(_05116_),
    .C(_05124_),
    .D(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__nor2_8 _19761_ (.A(\res_h_counter[5] ),
    .B(_08684_),
    .Y(_05141_));
 sky130_fd_sc_hd__and3_4 _19762_ (.A(_05141_),
    .B(_08709_),
    .C(_08662_),
    .X(_05142_));
 sky130_fd_sc_hd__and3_1 _19763_ (.A(_05142_),
    .B(_05020_),
    .C(_05068_),
    .X(_05143_));
 sky130_fd_sc_hd__buf_4 _19764_ (.A(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__clkinv_16 _19765_ (.A(_05142_),
    .Y(_05145_));
 sky130_fd_sc_hd__nor2_8 _19766_ (.A(_05074_),
    .B(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_2 _19767_ (.A(_05146_),
    .B(_05010_),
    .Y(_05147_));
 sky130_fd_sc_hd__nor2_4 _19768_ (.A(_05077_),
    .B(_05145_),
    .Y(_05148_));
 sky130_fd_sc_hd__nand2_2 _19769_ (.A(_05148_),
    .B(_05034_),
    .Y(_05149_));
 sky130_fd_sc_hd__nor2_4 _19770_ (.A(_05070_),
    .B(_05145_),
    .Y(_05150_));
 sky130_fd_sc_hd__buf_6 _19771_ (.A(_05021_),
    .X(_05151_));
 sky130_fd_sc_hd__nand2_1 _19772_ (.A(_05150_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__and4b_1 _19773_ (.A_N(_05144_),
    .B(_05147_),
    .C(_05149_),
    .D(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__nor2_1 _19774_ (.A(_05003_),
    .B(_05145_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand2_2 _19775_ (.A(_05154_),
    .B(_05010_),
    .Y(_05155_));
 sky130_fd_sc_hd__nor2_2 _19776_ (.A(_05025_),
    .B(_05145_),
    .Y(_05156_));
 sky130_fd_sc_hd__nand2_4 _19777_ (.A(_05156_),
    .B(_05020_),
    .Y(_05157_));
 sky130_fd_sc_hd__nor2_1 _19778_ (.A(_05013_),
    .B(_05145_),
    .Y(_05158_));
 sky130_fd_sc_hd__nand2_2 _19779_ (.A(_05158_),
    .B(_05010_),
    .Y(_05159_));
 sky130_fd_sc_hd__nor2_1 _19780_ (.A(_05018_),
    .B(_05145_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_2 _19781_ (.A(_05160_),
    .B(_05020_),
    .Y(_05161_));
 sky130_fd_sc_hd__and4_1 _19782_ (.A(_05155_),
    .B(_05157_),
    .C(_05159_),
    .D(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__nor2_8 _19783_ (.A(_05032_),
    .B(_05145_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2_2 _19784_ (.A(_05163_),
    .B(_05009_),
    .Y(_05164_));
 sky130_fd_sc_hd__nor2_8 _19785_ (.A(_05101_),
    .B(_05145_),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_1 _19786_ (.A(_05165_),
    .B(_05151_),
    .Y(_05166_));
 sky130_fd_sc_hd__nor2_8 _19787_ (.A(_05037_),
    .B(_05145_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand2_2 _19788_ (.A(_05167_),
    .B(_05010_),
    .Y(_05168_));
 sky130_fd_sc_hd__nor2_2 _19789_ (.A(_05044_),
    .B(_05145_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_2 _19790_ (.A(_05169_),
    .B(_05010_),
    .Y(_05170_));
 sky130_fd_sc_hd__and4_1 _19791_ (.A(_05164_),
    .B(_05166_),
    .C(_05168_),
    .D(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__inv_2 _19792_ (.A(_05054_),
    .Y(_05172_));
 sky130_fd_sc_hd__nor2_4 _19793_ (.A(_05172_),
    .B(_05145_),
    .Y(_05173_));
 sky130_fd_sc_hd__nand2_2 _19794_ (.A(_05173_),
    .B(_05034_),
    .Y(_05174_));
 sky130_fd_sc_hd__nor2_4 _19795_ (.A(_05057_),
    .B(_05145_),
    .Y(_05175_));
 sky130_fd_sc_hd__clkbuf_8 _19796_ (.A(_05010_),
    .X(_05176_));
 sky130_fd_sc_hd__nand2_2 _19797_ (.A(_05175_),
    .B(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__nor2_2 _19798_ (.A(_05051_),
    .B(_05145_),
    .Y(_05178_));
 sky130_fd_sc_hd__nand2_1 _19799_ (.A(_05178_),
    .B(_05151_),
    .Y(_05179_));
 sky130_fd_sc_hd__nor2_4 _19800_ (.A(_05062_),
    .B(_05145_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand2_2 _19801_ (.A(_05180_),
    .B(_05059_),
    .Y(_05181_));
 sky130_fd_sc_hd__and4_1 _19802_ (.A(_05174_),
    .B(_05177_),
    .C(_05179_),
    .D(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__and4_1 _19803_ (.A(_05153_),
    .B(_05162_),
    .C(_05171_),
    .D(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__and4_2 _19804_ (.A(_05082_),
    .B(_05086_),
    .C(_05140_),
    .D(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__buf_8 _19805_ (.A(_08678_),
    .X(_05185_));
 sky130_fd_sc_hd__clkbuf_16 _19806_ (.A(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__buf_6 _19807_ (.A(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__buf_6 _19808_ (.A(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__nand2_4 _19809_ (.A(\res_h_counter[6] ),
    .B(\res_h_counter[7] ),
    .Y(_05189_));
 sky130_fd_sc_hd__inv_4 _19810_ (.A(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand2_8 _19811_ (.A(_05004_),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__inv_2 _19812_ (.A(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__clkbuf_4 _19813_ (.A(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__buf_4 _19814_ (.A(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__nand2_8 _19815_ (.A(_05141_),
    .B(_05190_),
    .Y(_05195_));
 sky130_fd_sc_hd__nand2_8 _19816_ (.A(_05190_),
    .B(_05083_),
    .Y(_05196_));
 sky130_fd_sc_hd__a21oi_1 _19817_ (.A1(_05195_),
    .A2(_05196_),
    .B1(_05113_),
    .Y(_05197_));
 sky130_fd_sc_hd__nor2_4 _19818_ (.A(_05189_),
    .B(_05087_),
    .Y(_05198_));
 sky130_fd_sc_hd__inv_8 _19819_ (.A(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__nor2_8 _19820_ (.A(_08676_),
    .B(_05077_),
    .Y(_05200_));
 sky130_fd_sc_hd__clkinv_16 _19821_ (.A(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__nor2_4 _19822_ (.A(_05199_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__nor2_8 _19823_ (.A(_08676_),
    .B(_05070_),
    .Y(_05203_));
 sky130_fd_sc_hd__inv_16 _19824_ (.A(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__nor2_4 _19825_ (.A(_05199_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__buf_4 _19826_ (.A(_05198_),
    .X(_05206_));
 sky130_fd_sc_hd__nor2_8 _19827_ (.A(_08676_),
    .B(_05074_),
    .Y(_05207_));
 sky130_fd_sc_hd__inv_16 _19828_ (.A(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__nor2_4 _19829_ (.A(_05199_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__a31o_1 _19830_ (.A1(_05187_),
    .A2(_05068_),
    .A3(_05206_),
    .B1(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__nand2_8 _19831_ (.A(_05052_),
    .B(_08678_),
    .Y(_05211_));
 sky130_fd_sc_hd__nor2_2 _19832_ (.A(_05199_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_8 _19833_ (.A(_05054_),
    .B(_05099_),
    .Y(_05213_));
 sky130_fd_sc_hd__nor2_4 _19834_ (.A(_05199_),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__nor2_4 _19835_ (.A(_08676_),
    .B(_05057_),
    .Y(_05215_));
 sky130_fd_sc_hd__inv_12 _19836_ (.A(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nor2_2 _19837_ (.A(_05199_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__nor2_1 _19838_ (.A(_05062_),
    .B(_05199_),
    .Y(_05218_));
 sky130_fd_sc_hd__inv_2 _19839_ (.A(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__nor2_8 _19840_ (.A(_05020_),
    .B(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__or4_1 _19841_ (.A(_05212_),
    .B(_05214_),
    .C(_05217_),
    .D(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__or4_1 _19842_ (.A(_05202_),
    .B(_05205_),
    .C(_05210_),
    .D(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__nand2_8 _19843_ (.A(_05036_),
    .B(_08677_),
    .Y(_05223_));
 sky130_fd_sc_hd__nor2_4 _19844_ (.A(_05199_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__nand2_8 _19845_ (.A(_05031_),
    .B(_05099_),
    .Y(_05225_));
 sky130_fd_sc_hd__nor2_4 _19846_ (.A(_05199_),
    .B(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__nor2_8 _19847_ (.A(_08676_),
    .B(_05044_),
    .Y(_05227_));
 sky130_fd_sc_hd__inv_16 _19848_ (.A(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__nor2_4 _19849_ (.A(_05199_),
    .B(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__a31o_1 _19850_ (.A1(_05187_),
    .A2(_05042_),
    .A3(_05206_),
    .B1(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__nor2_8 _19851_ (.A(_08676_),
    .B(_05003_),
    .Y(_05231_));
 sky130_fd_sc_hd__clkinv_16 _19852_ (.A(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_4 _19853_ (.A(_05199_),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__nand2_8 _19854_ (.A(_05134_),
    .B(_05099_),
    .Y(_05234_));
 sky130_fd_sc_hd__nor2_2 _19855_ (.A(_05199_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__a31o_1 _19856_ (.A1(_05186_),
    .A2(_05130_),
    .A3(_05206_),
    .B1(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__a311o_1 _19857_ (.A1(_05187_),
    .A2(_05125_),
    .A3(_05206_),
    .B1(_05233_),
    .C1(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__or4_1 _19858_ (.A(_05224_),
    .B(_05226_),
    .C(_05230_),
    .D(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__a2111oi_2 _19859_ (.A1(_05188_),
    .A2(_05194_),
    .B1(_05197_),
    .C1(_05222_),
    .D1(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__nor2_8 _19860_ (.A(\res_h_counter[7] ),
    .B(_08709_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2_4 _19861_ (.A(_05240_),
    .B(_05004_),
    .Y(_05241_));
 sky130_fd_sc_hd__buf_12 _19862_ (.A(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__nand2_2 _19863_ (.A(_05240_),
    .B(_05141_),
    .Y(_05243_));
 sky130_fd_sc_hd__clkbuf_16 _19864_ (.A(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__nand2_8 _19865_ (.A(_05240_),
    .B(_05083_),
    .Y(_05245_));
 sky130_fd_sc_hd__nand2_8 _19866_ (.A(_05240_),
    .B(_05088_),
    .Y(_05246_));
 sky130_fd_sc_hd__a41o_1 _19867_ (.A1(_05242_),
    .A2(_05244_),
    .A3(_05245_),
    .A4(_05246_),
    .B1(_05113_),
    .X(_05247_));
 sky130_fd_sc_hd__nor2_8 _19868_ (.A(\res_h_counter[6] ),
    .B(_08662_),
    .Y(_05248_));
 sky130_fd_sc_hd__nand2_4 _19869_ (.A(_05004_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__buf_12 _19870_ (.A(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__nand2_2 _19871_ (.A(_05141_),
    .B(_05248_),
    .Y(_05251_));
 sky130_fd_sc_hd__buf_12 _19872_ (.A(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__nand2_8 _19873_ (.A(_05248_),
    .B(_05083_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2_2 _19874_ (.A(_05248_),
    .B(_05088_),
    .Y(_05254_));
 sky130_fd_sc_hd__buf_12 _19875_ (.A(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__a41o_1 _19876_ (.A1(_05250_),
    .A2(_05252_),
    .A3(_05253_),
    .A4(_05255_),
    .B1(_05113_),
    .X(_05256_));
 sky130_fd_sc_hd__and2_1 _19877_ (.A(_05247_),
    .B(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__nand3_4 _19878_ (.A(_05184_),
    .B(_05239_),
    .C(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__and3_1 _19879_ (.A(_05005_),
    .B(_05099_),
    .C(_05002_),
    .X(_05259_));
 sky130_fd_sc_hd__buf_2 _19880_ (.A(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__and3_4 _19881_ (.A(_05006_),
    .B(_05134_),
    .C(_08678_),
    .X(_05261_));
 sky130_fd_sc_hd__and3_4 _19882_ (.A(_05006_),
    .B(_08678_),
    .C(_05125_),
    .X(_05262_));
 sky130_fd_sc_hd__and3_4 _19883_ (.A(_05006_),
    .B(_05100_),
    .C(_05130_),
    .X(_05263_));
 sky130_fd_sc_hd__or4_1 _19884_ (.A(_05260_),
    .B(_05261_),
    .C(_05262_),
    .D(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__and3_1 _19885_ (.A(_05005_),
    .B(_05099_),
    .C(_05036_),
    .X(_05265_));
 sky130_fd_sc_hd__clkbuf_4 _19886_ (.A(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__and3_1 _19887_ (.A(_05005_),
    .B(_05045_),
    .C(_05099_),
    .X(_05267_));
 sky130_fd_sc_hd__clkbuf_4 _19888_ (.A(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__and3_1 _19889_ (.A(_05005_),
    .B(_05099_),
    .C(_05042_),
    .X(_05269_));
 sky130_fd_sc_hd__clkbuf_4 _19890_ (.A(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__and3_1 _19891_ (.A(_05005_),
    .B(_08678_),
    .C(_05031_),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_4 _19892_ (.A(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__or4_1 _19893_ (.A(_05266_),
    .B(_05268_),
    .C(_05270_),
    .D(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__and3_1 _19894_ (.A(_05005_),
    .B(_05099_),
    .C(_05068_),
    .X(_05274_));
 sky130_fd_sc_hd__clkbuf_4 _19895_ (.A(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__and3_1 _19896_ (.A(_05005_),
    .B(_05071_),
    .C(_05099_),
    .X(_05276_));
 sky130_fd_sc_hd__clkbuf_4 _19897_ (.A(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__and3_1 _19898_ (.A(_05005_),
    .B(_05099_),
    .C(_05075_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_4 _19899_ (.A(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__and3_1 _19900_ (.A(_05006_),
    .B(_08678_),
    .C(_05078_),
    .X(_05280_));
 sky130_fd_sc_hd__clkbuf_4 _19901_ (.A(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__or4_1 _19902_ (.A(_05275_),
    .B(_05277_),
    .C(_05279_),
    .D(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__and3_4 _19903_ (.A(_05006_),
    .B(_05100_),
    .C(_05054_),
    .X(_05283_));
 sky130_fd_sc_hd__inv_2 _19904_ (.A(_05057_),
    .Y(_05284_));
 sky130_fd_sc_hd__and3_4 _19905_ (.A(_05006_),
    .B(_05100_),
    .C(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__and3_1 _19906_ (.A(_05006_),
    .B(_05052_),
    .C(_08678_),
    .X(_05286_));
 sky130_fd_sc_hd__clkbuf_4 _19907_ (.A(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__nand2_1 _19908_ (.A(_05063_),
    .B(_05185_),
    .Y(_05288_));
 sky130_fd_sc_hd__or4b_1 _19909_ (.A(_05283_),
    .B(_05285_),
    .C(_05287_),
    .D_N(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__or4_1 _19910_ (.A(_05264_),
    .B(_05273_),
    .C(_05282_),
    .D(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__and3_1 _19911_ (.A(_05090_),
    .B(_08678_),
    .C(_05054_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_4 _19912_ (.A(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__and3_1 _19913_ (.A(_05090_),
    .B(_05100_),
    .C(_05052_),
    .X(_05293_));
 sky130_fd_sc_hd__clkbuf_4 _19914_ (.A(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__and3_1 _19915_ (.A(_05091_),
    .B(_05100_),
    .C(_05284_),
    .X(_05295_));
 sky130_fd_sc_hd__clkbuf_4 _19916_ (.A(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__a2111o_1 _19917_ (.A1(_05111_),
    .A2(_05186_),
    .B1(_05292_),
    .C1(_05294_),
    .D1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__and3_4 _19918_ (.A(_05090_),
    .B(_05002_),
    .C(_08678_),
    .X(_05298_));
 sky130_fd_sc_hd__and3_1 _19919_ (.A(_05090_),
    .B(_05099_),
    .C(_05125_),
    .X(_05299_));
 sky130_fd_sc_hd__clkbuf_4 _19920_ (.A(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__and3_4 _19921_ (.A(_05091_),
    .B(_05100_),
    .C(_05130_),
    .X(_05301_));
 sky130_fd_sc_hd__and3_4 _19922_ (.A(_05091_),
    .B(_05100_),
    .C(_05134_),
    .X(_05302_));
 sky130_fd_sc_hd__or4_1 _19923_ (.A(_05298_),
    .B(_05300_),
    .C(_05301_),
    .D(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__and3_4 _19924_ (.A(_05090_),
    .B(_05036_),
    .C(_08678_),
    .X(_05304_));
 sky130_fd_sc_hd__and3_1 _19925_ (.A(_05090_),
    .B(_08678_),
    .C(_05031_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_4 _19926_ (.A(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__and3_4 _19927_ (.A(_05091_),
    .B(_05100_),
    .C(_05042_),
    .X(_05307_));
 sky130_fd_sc_hd__nand2_1 _19928_ (.A(_05095_),
    .B(_05185_),
    .Y(_05308_));
 sky130_fd_sc_hd__clkinv_4 _19929_ (.A(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__or4_1 _19930_ (.A(_05304_),
    .B(_05306_),
    .C(_05307_),
    .D(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__and3_1 _19931_ (.A(_05090_),
    .B(_08678_),
    .C(_05078_),
    .X(_05311_));
 sky130_fd_sc_hd__clkbuf_4 _19932_ (.A(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__and3_1 _19933_ (.A(_05090_),
    .B(_05068_),
    .C(_08678_),
    .X(_05313_));
 sky130_fd_sc_hd__clkbuf_4 _19934_ (.A(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__and3_4 _19935_ (.A(_05091_),
    .B(_05185_),
    .C(_05075_),
    .X(_05315_));
 sky130_fd_sc_hd__nand2_1 _19936_ (.A(_05117_),
    .B(_05185_),
    .Y(_05316_));
 sky130_fd_sc_hd__inv_2 _19937_ (.A(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__or4_1 _19938_ (.A(_05312_),
    .B(_05314_),
    .C(_05315_),
    .D(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__or4_1 _19939_ (.A(_05297_),
    .B(_05303_),
    .C(_05310_),
    .D(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__nor2_4 _19940_ (.A(_05067_),
    .B(_05145_),
    .Y(_05320_));
 sky130_fd_sc_hd__o41a_1 _19941_ (.A1(_05146_),
    .A2(_05148_),
    .A3(_05150_),
    .A4(_05320_),
    .B1(_05186_),
    .X(_05321_));
 sky130_fd_sc_hd__nand2_2 _19942_ (.A(_05165_),
    .B(_05100_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand2_4 _19943_ (.A(_05169_),
    .B(_05100_),
    .Y(_05323_));
 sky130_fd_sc_hd__nand2_1 _19944_ (.A(_05322_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__nand2_2 _19945_ (.A(_05160_),
    .B(_05100_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_4 _19946_ (.A(_05156_),
    .B(_05100_),
    .Y(_05326_));
 sky130_fd_sc_hd__nand2_1 _19947_ (.A(_05325_),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__o21a_1 _19948_ (.A1(_05167_),
    .A2(_05163_),
    .B1(_05100_),
    .X(_05328_));
 sky130_fd_sc_hd__and3_4 _19949_ (.A(_05142_),
    .B(_08677_),
    .C(_05002_),
    .X(_05329_));
 sky130_fd_sc_hd__and3_4 _19950_ (.A(_05142_),
    .B(_08677_),
    .C(_05125_),
    .X(_05330_));
 sky130_fd_sc_hd__or2_1 _19951_ (.A(_05329_),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__or4_1 _19952_ (.A(_05324_),
    .B(_05327_),
    .C(_05328_),
    .D(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__nand2_1 _19953_ (.A(_05175_),
    .B(_05185_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand2_1 _19954_ (.A(_05173_),
    .B(_05185_),
    .Y(_05334_));
 sky130_fd_sc_hd__nand2_1 _19955_ (.A(_05178_),
    .B(_05185_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand2_1 _19956_ (.A(_05180_),
    .B(_05185_),
    .Y(_05336_));
 sky130_fd_sc_hd__and4_1 _19957_ (.A(_05333_),
    .B(_05334_),
    .C(_05335_),
    .D(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__or3b_1 _19958_ (.A(_05321_),
    .B(_05332_),
    .C_N(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__o311a_1 _19959_ (.A1(_05134_),
    .A2(_05125_),
    .A3(_05130_),
    .B1(_05186_),
    .C1(_05085_),
    .X(_05339_));
 sky130_fd_sc_hd__inv_6 _19960_ (.A(_05085_),
    .Y(_05340_));
 sky130_fd_sc_hd__nor2_1 _19961_ (.A(_05037_),
    .B(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__and3_1 _19962_ (.A(_05085_),
    .B(_05099_),
    .C(_05031_),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_4 _19963_ (.A(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__nor2_1 _19964_ (.A(_05044_),
    .B(_05340_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand2_1 _19965_ (.A(_05344_),
    .B(_05100_),
    .Y(_05345_));
 sky130_fd_sc_hd__clkinv_4 _19966_ (.A(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__and3_1 _19967_ (.A(_05085_),
    .B(_05099_),
    .C(_05042_),
    .X(_05347_));
 sky130_fd_sc_hd__clkbuf_4 _19968_ (.A(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__a2111o_1 _19969_ (.A1(_05185_),
    .A2(_05341_),
    .B1(_05343_),
    .C1(_05346_),
    .D1(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__and3_1 _19970_ (.A(_05085_),
    .B(_08677_),
    .C(_05075_),
    .X(_05350_));
 sky130_fd_sc_hd__clkbuf_4 _19971_ (.A(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__and3_1 _19972_ (.A(_05085_),
    .B(_08677_),
    .C(_05078_),
    .X(_05352_));
 sky130_fd_sc_hd__clkbuf_4 _19973_ (.A(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__and3_1 _19974_ (.A(_05085_),
    .B(_08677_),
    .C(_05068_),
    .X(_05354_));
 sky130_fd_sc_hd__clkbuf_4 _19975_ (.A(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__nor2_4 _19976_ (.A(_05070_),
    .B(_05340_),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_1 _19977_ (.A(_05356_),
    .B(_08678_),
    .Y(_05357_));
 sky130_fd_sc_hd__inv_2 _19978_ (.A(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__or4_1 _19979_ (.A(_05351_),
    .B(_05353_),
    .C(_05355_),
    .D(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__nor2_1 _19980_ (.A(_05172_),
    .B(_05340_),
    .Y(_05360_));
 sky130_fd_sc_hd__nand2_1 _19981_ (.A(_05360_),
    .B(_05185_),
    .Y(_05361_));
 sky130_fd_sc_hd__nor2_1 _19982_ (.A(_05057_),
    .B(_05340_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_1 _19983_ (.A(_05362_),
    .B(_05185_),
    .Y(_05363_));
 sky130_fd_sc_hd__nor2_8 _19984_ (.A(_05051_),
    .B(_05340_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_4 _19985_ (.A(_05364_),
    .B(_05185_),
    .Y(_05365_));
 sky130_fd_sc_hd__nor2_1 _19986_ (.A(_05062_),
    .B(_05340_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _19987_ (.A(_05366_),
    .B(_05185_),
    .Y(_05367_));
 sky130_fd_sc_hd__and4_1 _19988_ (.A(_05361_),
    .B(_05363_),
    .C(_05365_),
    .D(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__or4b_1 _19989_ (.A(_05339_),
    .B(_05349_),
    .C(_05359_),
    .D_N(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__or2_1 _19990_ (.A(_05338_),
    .B(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__or3_2 _19991_ (.A(_05290_),
    .B(_05319_),
    .C(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__buf_2 _19992_ (.A(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__nor3b_1 _19993_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][0] ),
    .Y(_05373_));
 sky130_fd_sc_hd__nor2_4 _19994_ (.A(_05253_),
    .B(_05216_),
    .Y(_05374_));
 sky130_fd_sc_hd__nor2_4 _19995_ (.A(_05253_),
    .B(_05213_),
    .Y(_05375_));
 sky130_fd_sc_hd__nor2_4 _19996_ (.A(_05253_),
    .B(_05211_),
    .Y(_05376_));
 sky130_fd_sc_hd__nor2_4 _19997_ (.A(_05253_),
    .B(_05204_),
    .Y(_05377_));
 sky130_fd_sc_hd__a22o_1 _19998_ (.A1(_05376_),
    .A2(\line_cache[140][0] ),
    .B1(_05377_),
    .B2(\line_cache[139][0] ),
    .X(_05378_));
 sky130_fd_sc_hd__a221o_1 _19999_ (.A1(\line_cache[142][0] ),
    .A2(_05374_),
    .B1(\line_cache[141][0] ),
    .B2(_05375_),
    .C1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__nor2_4 _20000_ (.A(_05252_),
    .B(_05232_),
    .Y(_05380_));
 sky130_fd_sc_hd__clkinv_4 _20001_ (.A(_05253_),
    .Y(_05381_));
 sky130_fd_sc_hd__and3_4 _20002_ (.A(_05381_),
    .B(_05185_),
    .C(_05061_),
    .X(_05382_));
 sky130_fd_sc_hd__nand2_8 _20003_ (.A(_05125_),
    .B(_05099_),
    .Y(_05383_));
 sky130_fd_sc_hd__nor2_4 _20004_ (.A(_05252_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__nand2_8 _20005_ (.A(_05130_),
    .B(_08677_),
    .Y(_05385_));
 sky130_fd_sc_hd__nor2_2 _20006_ (.A(_05252_),
    .B(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__a22o_1 _20007_ (.A1(_05384_),
    .A2(\line_cache[145][0] ),
    .B1(\line_cache[146][0] ),
    .B2(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__a221o_1 _20008_ (.A1(\line_cache[144][0] ),
    .A2(_05380_),
    .B1(\line_cache[143][0] ),
    .B2(_05382_),
    .C1(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__nand2_8 _20009_ (.A(_05042_),
    .B(_05099_),
    .Y(_05389_));
 sky130_fd_sc_hd__nor2_4 _20010_ (.A(_05252_),
    .B(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__nor2_2 _20011_ (.A(_05252_),
    .B(_05225_),
    .Y(_05391_));
 sky130_fd_sc_hd__nor2_4 _20012_ (.A(_05252_),
    .B(_05234_),
    .Y(_05392_));
 sky130_fd_sc_hd__nor2_4 _20013_ (.A(_05252_),
    .B(_05223_),
    .Y(_05393_));
 sky130_fd_sc_hd__a22o_1 _20014_ (.A1(_05392_),
    .A2(\line_cache[147][0] ),
    .B1(_05393_),
    .B2(\line_cache[148][0] ),
    .X(_05394_));
 sky130_fd_sc_hd__a221o_1 _20015_ (.A1(\line_cache[150][0] ),
    .A2(_05390_),
    .B1(\line_cache[149][0] ),
    .B2(_05391_),
    .C1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__nand2_8 _20016_ (.A(_05068_),
    .B(_08678_),
    .Y(_05396_));
 sky130_fd_sc_hd__nor2_4 _20017_ (.A(_05252_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__nor2_4 _20018_ (.A(_05252_),
    .B(_05228_),
    .Y(_05398_));
 sky130_fd_sc_hd__nor2_4 _20019_ (.A(_05252_),
    .B(_05208_),
    .Y(_05399_));
 sky130_fd_sc_hd__inv_2 _20020_ (.A(_05251_),
    .Y(_05400_));
 sky130_fd_sc_hd__and3_1 _20021_ (.A(_05200_),
    .B(\line_cache[154][0] ),
    .C(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__a21o_1 _20022_ (.A1(\line_cache[153][0] ),
    .A2(_05399_),
    .B1(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__a221oi_1 _20023_ (.A1(\line_cache[152][0] ),
    .A2(_05397_),
    .B1(\line_cache[151][0] ),
    .B2(_05398_),
    .C1(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__or2b_1 _20024_ (.A(_05395_),
    .B_N(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__or3_1 _20025_ (.A(_05379_),
    .B(_05388_),
    .C(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__nor2_4 _20026_ (.A(_05250_),
    .B(_05383_),
    .Y(_05406_));
 sky130_fd_sc_hd__inv_2 _20027_ (.A(_05385_),
    .Y(_05407_));
 sky130_fd_sc_hd__clkbuf_8 _20028_ (.A(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__buf_6 _20029_ (.A(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__inv_2 _20030_ (.A(_05250_),
    .Y(_05410_));
 sky130_fd_sc_hd__and3_1 _20031_ (.A(_05409_),
    .B(\line_cache[162][0] ),
    .C(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__and3_1 _20032_ (.A(_05400_),
    .B(_05186_),
    .C(_05061_),
    .X(_05412_));
 sky130_fd_sc_hd__buf_2 _20033_ (.A(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__nor2_4 _20034_ (.A(_05250_),
    .B(_05232_),
    .Y(_05414_));
 sky130_fd_sc_hd__a22o_1 _20035_ (.A1(_05413_),
    .A2(\line_cache[159][0] ),
    .B1(_05414_),
    .B2(\line_cache[160][0] ),
    .X(_05415_));
 sky130_fd_sc_hd__nor2_4 _20036_ (.A(_05252_),
    .B(_05216_),
    .Y(_05416_));
 sky130_fd_sc_hd__nor2_4 _20037_ (.A(_05252_),
    .B(_05213_),
    .Y(_05417_));
 sky130_fd_sc_hd__nor2_4 _20038_ (.A(_05252_),
    .B(_05211_),
    .Y(_05418_));
 sky130_fd_sc_hd__nor2_4 _20039_ (.A(_05252_),
    .B(_05204_),
    .Y(_05419_));
 sky130_fd_sc_hd__a22o_1 _20040_ (.A1(_05418_),
    .A2(\line_cache[156][0] ),
    .B1(_05419_),
    .B2(\line_cache[155][0] ),
    .X(_05420_));
 sky130_fd_sc_hd__a221o_1 _20041_ (.A1(\line_cache[158][0] ),
    .A2(_05416_),
    .B1(\line_cache[157][0] ),
    .B2(_05417_),
    .C1(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__a2111oi_1 _20042_ (.A1(\line_cache[161][0] ),
    .A2(_05406_),
    .B1(_05411_),
    .C1(_05415_),
    .D1(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__nor2_2 _20043_ (.A(_05250_),
    .B(_05208_),
    .Y(_05423_));
 sky130_fd_sc_hd__nor2_4 _20044_ (.A(_05250_),
    .B(_05201_),
    .Y(_05424_));
 sky130_fd_sc_hd__nor2_4 _20045_ (.A(_05250_),
    .B(_05228_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _20046_ (.A(_05425_),
    .B(\line_cache[167][0] ),
    .Y(_05426_));
 sky130_fd_sc_hd__nor2_2 _20047_ (.A(_05250_),
    .B(_05396_),
    .Y(_05427_));
 sky130_fd_sc_hd__nand2_1 _20048_ (.A(_05427_),
    .B(\line_cache[168][0] ),
    .Y(_05428_));
 sky130_fd_sc_hd__nand2_1 _20049_ (.A(_05426_),
    .B(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__a221oi_2 _20050_ (.A1(_05423_),
    .A2(\line_cache[169][0] ),
    .B1(\line_cache[170][0] ),
    .B2(_05424_),
    .C1(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__nor2_4 _20051_ (.A(_05250_),
    .B(_05389_),
    .Y(_05431_));
 sky130_fd_sc_hd__nor2_2 _20052_ (.A(_05250_),
    .B(_05225_),
    .Y(_05432_));
 sky130_fd_sc_hd__nor2_4 _20053_ (.A(_05250_),
    .B(_05234_),
    .Y(_05433_));
 sky130_fd_sc_hd__nor2_4 _20054_ (.A(_05250_),
    .B(_05223_),
    .Y(_05434_));
 sky130_fd_sc_hd__a22o_1 _20055_ (.A1(_05433_),
    .A2(\line_cache[163][0] ),
    .B1(_05434_),
    .B2(\line_cache[164][0] ),
    .X(_05435_));
 sky130_fd_sc_hd__a221oi_1 _20056_ (.A1(\line_cache[166][0] ),
    .A2(_05431_),
    .B1(\line_cache[165][0] ),
    .B2(_05432_),
    .C1(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__and4b_2 _20057_ (.A_N(_05405_),
    .B(_05422_),
    .C(_05430_),
    .D(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__nor2_4 _20058_ (.A(_05255_),
    .B(_05396_),
    .Y(_05438_));
 sky130_fd_sc_hd__nor2_4 _20059_ (.A(_05255_),
    .B(_05228_),
    .Y(_05439_));
 sky130_fd_sc_hd__nor2_4 _20060_ (.A(_05255_),
    .B(_05208_),
    .Y(_05440_));
 sky130_fd_sc_hd__inv_2 _20061_ (.A(_05254_),
    .Y(_05441_));
 sky130_fd_sc_hd__and3_1 _20062_ (.A(_05200_),
    .B(\line_cache[186][0] ),
    .C(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__a21o_1 _20063_ (.A1(\line_cache[185][0] ),
    .A2(_05440_),
    .B1(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__a221o_1 _20064_ (.A1(\line_cache[184][0] ),
    .A2(_05438_),
    .B1(\line_cache[183][0] ),
    .B2(_05439_),
    .C1(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__nor2_4 _20065_ (.A(_05255_),
    .B(_05389_),
    .Y(_05445_));
 sky130_fd_sc_hd__nor2_2 _20066_ (.A(_05255_),
    .B(_05225_),
    .Y(_05446_));
 sky130_fd_sc_hd__nor2_4 _20067_ (.A(_05255_),
    .B(_05234_),
    .Y(_05447_));
 sky130_fd_sc_hd__and2_1 _20068_ (.A(_05447_),
    .B(\line_cache[179][0] ),
    .X(_05448_));
 sky130_fd_sc_hd__nor2_2 _20069_ (.A(_05255_),
    .B(_05223_),
    .Y(_05449_));
 sky130_fd_sc_hd__and2_1 _20070_ (.A(_05449_),
    .B(\line_cache[180][0] ),
    .X(_05450_));
 sky130_fd_sc_hd__or2_1 _20071_ (.A(_05448_),
    .B(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__a221o_1 _20072_ (.A1(\line_cache[182][0] ),
    .A2(_05445_),
    .B1(\line_cache[181][0] ),
    .B2(_05446_),
    .C1(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__nor2_4 _20073_ (.A(_05255_),
    .B(_05232_),
    .Y(_05453_));
 sky130_fd_sc_hd__nor2_8 _20074_ (.A(_08676_),
    .B(_05062_),
    .Y(_05454_));
 sky130_fd_sc_hd__inv_4 _20075_ (.A(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__nor2_4 _20076_ (.A(_05250_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__nor2_4 _20077_ (.A(_05255_),
    .B(_05383_),
    .Y(_05457_));
 sky130_fd_sc_hd__nor2_4 _20078_ (.A(_05255_),
    .B(_05385_),
    .Y(_05458_));
 sky130_fd_sc_hd__a22o_1 _20079_ (.A1(_05457_),
    .A2(\line_cache[177][0] ),
    .B1(\line_cache[178][0] ),
    .B2(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__a221o_1 _20080_ (.A1(\line_cache[176][0] ),
    .A2(_05453_),
    .B1(\line_cache[175][0] ),
    .B2(_05456_),
    .C1(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__nor2_4 _20081_ (.A(_05250_),
    .B(_05216_),
    .Y(_05461_));
 sky130_fd_sc_hd__nor2_2 _20082_ (.A(_05250_),
    .B(_05213_),
    .Y(_05462_));
 sky130_fd_sc_hd__nor2_4 _20083_ (.A(_05249_),
    .B(_05211_),
    .Y(_05463_));
 sky130_fd_sc_hd__nor2_4 _20084_ (.A(_05250_),
    .B(_05204_),
    .Y(_05464_));
 sky130_fd_sc_hd__a22o_1 _20085_ (.A1(_05463_),
    .A2(\line_cache[172][0] ),
    .B1(_05464_),
    .B2(\line_cache[171][0] ),
    .X(_05465_));
 sky130_fd_sc_hd__a221o_1 _20086_ (.A1(\line_cache[174][0] ),
    .A2(_05461_),
    .B1(\line_cache[173][0] ),
    .B2(_05462_),
    .C1(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__or4_1 _20087_ (.A(_05444_),
    .B(_05452_),
    .C(_05460_),
    .D(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__nor2_4 _20088_ (.A(_05255_),
    .B(_05455_),
    .Y(_05468_));
 sky130_fd_sc_hd__inv_2 _20089_ (.A(_05383_),
    .Y(_05469_));
 sky130_fd_sc_hd__buf_4 _20090_ (.A(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__inv_2 _20091_ (.A(_05196_),
    .Y(_05471_));
 sky130_fd_sc_hd__clkbuf_4 _20092_ (.A(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__and3_1 _20093_ (.A(_05470_),
    .B(\line_cache[193][0] ),
    .C(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__and3_1 _20094_ (.A(_05409_),
    .B(\line_cache[194][0] ),
    .C(_05472_),
    .X(_05474_));
 sky130_fd_sc_hd__buf_4 _20095_ (.A(_05231_),
    .X(_05475_));
 sky130_fd_sc_hd__and3_1 _20096_ (.A(_05475_),
    .B(\line_cache[192][0] ),
    .C(_05472_),
    .X(_05476_));
 sky130_fd_sc_hd__a2111o_1 _20097_ (.A1(\line_cache[191][0] ),
    .A2(_05468_),
    .B1(_05473_),
    .C1(_05474_),
    .D1(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__nor2_4 _20098_ (.A(_05255_),
    .B(_05216_),
    .Y(_05478_));
 sky130_fd_sc_hd__nor2_4 _20099_ (.A(_05255_),
    .B(_05213_),
    .Y(_05479_));
 sky130_fd_sc_hd__nor2_4 _20100_ (.A(_05255_),
    .B(_05211_),
    .Y(_05480_));
 sky130_fd_sc_hd__nor2_4 _20101_ (.A(_05255_),
    .B(_05204_),
    .Y(_05481_));
 sky130_fd_sc_hd__a22o_1 _20102_ (.A1(_05480_),
    .A2(\line_cache[188][0] ),
    .B1(_05481_),
    .B2(\line_cache[187][0] ),
    .X(_05482_));
 sky130_fd_sc_hd__a221o_2 _20103_ (.A1(\line_cache[190][0] ),
    .A2(_05478_),
    .B1(\line_cache[189][0] ),
    .B2(_05479_),
    .C1(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__nor2_2 _20104_ (.A(_05196_),
    .B(_05234_),
    .Y(_05484_));
 sky130_fd_sc_hd__nor2_4 _20105_ (.A(_05196_),
    .B(_05223_),
    .Y(_05485_));
 sky130_fd_sc_hd__a22o_1 _20106_ (.A1(_05484_),
    .A2(\line_cache[195][0] ),
    .B1(_05485_),
    .B2(\line_cache[196][0] ),
    .X(_05486_));
 sky130_fd_sc_hd__nor2_2 _20107_ (.A(_05196_),
    .B(_05389_),
    .Y(_05487_));
 sky130_fd_sc_hd__and2_1 _20108_ (.A(_05487_),
    .B(\line_cache[198][0] ),
    .X(_05488_));
 sky130_fd_sc_hd__nor2_4 _20109_ (.A(_05196_),
    .B(_05225_),
    .Y(_05489_));
 sky130_fd_sc_hd__and2_1 _20110_ (.A(_05489_),
    .B(\line_cache[197][0] ),
    .X(_05490_));
 sky130_fd_sc_hd__nor2_2 _20111_ (.A(_05196_),
    .B(_05208_),
    .Y(_05491_));
 sky130_fd_sc_hd__nor2_2 _20112_ (.A(_05196_),
    .B(_05201_),
    .Y(_05492_));
 sky130_fd_sc_hd__nor2_2 _20113_ (.A(_05196_),
    .B(_05228_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(_05493_),
    .B(\line_cache[199][0] ),
    .Y(_05494_));
 sky130_fd_sc_hd__nor2_2 _20115_ (.A(_05196_),
    .B(_05396_),
    .Y(_05495_));
 sky130_fd_sc_hd__nand2_1 _20116_ (.A(_05495_),
    .B(\line_cache[200][0] ),
    .Y(_05496_));
 sky130_fd_sc_hd__nand2_1 _20117_ (.A(_05494_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__a221oi_1 _20118_ (.A1(_05491_),
    .A2(\line_cache[201][0] ),
    .B1(\line_cache[202][0] ),
    .B2(_05492_),
    .C1(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__or4b_1 _20119_ (.A(_05486_),
    .B(_05488_),
    .C(_05490_),
    .D_N(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__or3_4 _20120_ (.A(_05477_),
    .B(_05483_),
    .C(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__nor2_1 _20121_ (.A(_05467_),
    .B(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hd__nor2_2 _20122_ (.A(_05241_),
    .B(_05389_),
    .Y(_05502_));
 sky130_fd_sc_hd__nor2_4 _20123_ (.A(_05242_),
    .B(_05396_),
    .Y(_05503_));
 sky130_fd_sc_hd__nor2_4 _20124_ (.A(_05242_),
    .B(_05228_),
    .Y(_05504_));
 sky130_fd_sc_hd__a22o_1 _20125_ (.A1(_05503_),
    .A2(\line_cache[104][0] ),
    .B1(_05504_),
    .B2(\line_cache[103][0] ),
    .X(_05505_));
 sky130_fd_sc_hd__nor2_4 _20126_ (.A(_05242_),
    .B(_05201_),
    .Y(_05506_));
 sky130_fd_sc_hd__and2_1 _20127_ (.A(_05506_),
    .B(\line_cache[106][0] ),
    .X(_05507_));
 sky130_fd_sc_hd__nor2_4 _20128_ (.A(_05242_),
    .B(_05208_),
    .Y(_05508_));
 sky130_fd_sc_hd__nor2_2 _20129_ (.A(_05242_),
    .B(_05225_),
    .Y(_05509_));
 sky130_fd_sc_hd__nor2_4 _20130_ (.A(_05242_),
    .B(_05234_),
    .Y(_05510_));
 sky130_fd_sc_hd__nor2_2 _20131_ (.A(_05242_),
    .B(_05223_),
    .Y(_05511_));
 sky130_fd_sc_hd__a22o_1 _20132_ (.A1(_05510_),
    .A2(\line_cache[99][0] ),
    .B1(_05511_),
    .B2(\line_cache[100][0] ),
    .X(_05512_));
 sky130_fd_sc_hd__a221o_1 _20133_ (.A1(\line_cache[105][0] ),
    .A2(_05508_),
    .B1(\line_cache[101][0] ),
    .B2(_05509_),
    .C1(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__a2111o_1 _20134_ (.A1(\line_cache[102][0] ),
    .A2(_05502_),
    .B1(_05505_),
    .C1(_05507_),
    .D1(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__nor2_4 _20135_ (.A(_05242_),
    .B(_05383_),
    .Y(_05515_));
 sky130_fd_sc_hd__nor2_4 _20136_ (.A(_05242_),
    .B(_05385_),
    .Y(_05516_));
 sky130_fd_sc_hd__and2_1 _20137_ (.A(_05516_),
    .B(\line_cache[98][0] ),
    .X(_05517_));
 sky130_fd_sc_hd__inv_2 _20138_ (.A(_05243_),
    .Y(_05518_));
 sky130_fd_sc_hd__and3_4 _20139_ (.A(_05518_),
    .B(_05185_),
    .C(_05061_),
    .X(_05519_));
 sky130_fd_sc_hd__nor2_4 _20140_ (.A(_05242_),
    .B(_05232_),
    .Y(_05520_));
 sky130_fd_sc_hd__a22o_1 _20141_ (.A1(_05519_),
    .A2(\line_cache[95][0] ),
    .B1(_05520_),
    .B2(\line_cache[96][0] ),
    .X(_05521_));
 sky130_fd_sc_hd__nor2_4 _20142_ (.A(_05244_),
    .B(_05216_),
    .Y(_05522_));
 sky130_fd_sc_hd__nor2_4 _20143_ (.A(_05244_),
    .B(_05213_),
    .Y(_05523_));
 sky130_fd_sc_hd__nor2_2 _20144_ (.A(_05244_),
    .B(_05211_),
    .Y(_05524_));
 sky130_fd_sc_hd__nor2_4 _20145_ (.A(_05244_),
    .B(_05204_),
    .Y(_05525_));
 sky130_fd_sc_hd__a22o_1 _20146_ (.A1(_05524_),
    .A2(\line_cache[92][0] ),
    .B1(_05525_),
    .B2(\line_cache[91][0] ),
    .X(_05526_));
 sky130_fd_sc_hd__a221o_1 _20147_ (.A1(\line_cache[94][0] ),
    .A2(_05522_),
    .B1(\line_cache[93][0] ),
    .B2(_05523_),
    .C1(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__a2111oi_1 _20148_ (.A1(\line_cache[97][0] ),
    .A2(_05515_),
    .B1(_05517_),
    .C1(_05521_),
    .D1(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__nor2_2 _20149_ (.A(_05244_),
    .B(_05389_),
    .Y(_05529_));
 sky130_fd_sc_hd__nor2_2 _20150_ (.A(_05244_),
    .B(_05225_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_4 _20151_ (.A(_05244_),
    .B(_05234_),
    .Y(_05531_));
 sky130_fd_sc_hd__nor2_2 _20152_ (.A(_05244_),
    .B(_05223_),
    .Y(_05532_));
 sky130_fd_sc_hd__a22o_1 _20153_ (.A1(_05531_),
    .A2(\line_cache[83][0] ),
    .B1(_05532_),
    .B2(\line_cache[84][0] ),
    .X(_05533_));
 sky130_fd_sc_hd__a221o_1 _20154_ (.A1(\line_cache[86][0] ),
    .A2(_05529_),
    .B1(\line_cache[85][0] ),
    .B2(_05530_),
    .C1(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__nor2_4 _20155_ (.A(_05244_),
    .B(_05232_),
    .Y(_05535_));
 sky130_fd_sc_hd__clkinv_4 _20156_ (.A(_05245_),
    .Y(_05536_));
 sky130_fd_sc_hd__and3_4 _20157_ (.A(_05536_),
    .B(_05100_),
    .C(_05061_),
    .X(_05537_));
 sky130_fd_sc_hd__nor2_4 _20158_ (.A(_05244_),
    .B(_05383_),
    .Y(_05538_));
 sky130_fd_sc_hd__nor2_4 _20159_ (.A(_05244_),
    .B(_05385_),
    .Y(_05539_));
 sky130_fd_sc_hd__a22o_1 _20160_ (.A1(_05538_),
    .A2(\line_cache[81][0] ),
    .B1(\line_cache[82][0] ),
    .B2(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__a221o_1 _20161_ (.A1(\line_cache[80][0] ),
    .A2(_05535_),
    .B1(\line_cache[79][0] ),
    .B2(_05537_),
    .C1(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__nor2_4 _20162_ (.A(_05245_),
    .B(_05211_),
    .Y(_05542_));
 sky130_fd_sc_hd__nor2_4 _20163_ (.A(_05245_),
    .B(_05204_),
    .Y(_05543_));
 sky130_fd_sc_hd__inv_2 _20164_ (.A(_05213_),
    .Y(_05544_));
 sky130_fd_sc_hd__nor2_4 _20165_ (.A(_05245_),
    .B(_05216_),
    .Y(_05545_));
 sky130_fd_sc_hd__a32o_1 _20166_ (.A1(_05544_),
    .A2(\line_cache[77][0] ),
    .A3(_05536_),
    .B1(_05545_),
    .B2(\line_cache[78][0] ),
    .X(_05546_));
 sky130_fd_sc_hd__a221o_1 _20167_ (.A1(\line_cache[76][0] ),
    .A2(_05542_),
    .B1(\line_cache[75][0] ),
    .B2(_05543_),
    .C1(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__nor2_1 _20168_ (.A(_05541_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__nor2_2 _20169_ (.A(_05244_),
    .B(_05208_),
    .Y(_05549_));
 sky130_fd_sc_hd__nor2_4 _20170_ (.A(_05244_),
    .B(_05201_),
    .Y(_05550_));
 sky130_fd_sc_hd__nor2_2 _20171_ (.A(_05244_),
    .B(_05228_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_1 _20172_ (.A(_05551_),
    .B(\line_cache[87][0] ),
    .Y(_05552_));
 sky130_fd_sc_hd__nor2_2 _20173_ (.A(_05244_),
    .B(_05396_),
    .Y(_05553_));
 sky130_fd_sc_hd__nand2_1 _20174_ (.A(_05553_),
    .B(\line_cache[88][0] ),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_1 _20175_ (.A(_05552_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__a221oi_2 _20176_ (.A1(_05549_),
    .A2(\line_cache[89][0] ),
    .B1(\line_cache[90][0] ),
    .B2(_05550_),
    .C1(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__and3b_1 _20177_ (.A_N(_05534_),
    .B(_05548_),
    .C(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__and3b_1 _20178_ (.A_N(_05514_),
    .B(_05528_),
    .C(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__nor2_4 _20179_ (.A(_05246_),
    .B(_05201_),
    .Y(_05559_));
 sky130_fd_sc_hd__nor2_1 _20180_ (.A(_05246_),
    .B(_05208_),
    .Y(_05560_));
 sky130_fd_sc_hd__nor2_4 _20181_ (.A(_05246_),
    .B(_05396_),
    .Y(_05561_));
 sky130_fd_sc_hd__clkinv_4 _20182_ (.A(_05246_),
    .Y(_05562_));
 sky130_fd_sc_hd__and3_1 _20183_ (.A(_05227_),
    .B(\line_cache[119][0] ),
    .C(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__a21o_1 _20184_ (.A1(\line_cache[120][0] ),
    .A2(_05561_),
    .B1(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__a221o_1 _20185_ (.A1(\line_cache[122][0] ),
    .A2(_05559_),
    .B1(\line_cache[121][0] ),
    .B2(_05560_),
    .C1(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__nor2_4 _20186_ (.A(_05246_),
    .B(_05389_),
    .Y(_05566_));
 sky130_fd_sc_hd__nor2_2 _20187_ (.A(_05246_),
    .B(_05225_),
    .Y(_05567_));
 sky130_fd_sc_hd__nor2_2 _20188_ (.A(_05246_),
    .B(_05223_),
    .Y(_05568_));
 sky130_fd_sc_hd__nor2_2 _20189_ (.A(_05246_),
    .B(_05234_),
    .Y(_05569_));
 sky130_fd_sc_hd__and2_1 _20190_ (.A(_05569_),
    .B(\line_cache[115][0] ),
    .X(_05570_));
 sky130_fd_sc_hd__a21o_1 _20191_ (.A1(\line_cache[116][0] ),
    .A2(_05568_),
    .B1(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__a221o_1 _20192_ (.A1(\line_cache[118][0] ),
    .A2(_05566_),
    .B1(\line_cache[117][0] ),
    .B2(_05567_),
    .C1(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__nor2_4 _20193_ (.A(_05242_),
    .B(_05216_),
    .Y(_05573_));
 sky130_fd_sc_hd__nor2_4 _20194_ (.A(_05242_),
    .B(_05213_),
    .Y(_05574_));
 sky130_fd_sc_hd__nor2_4 _20195_ (.A(_05242_),
    .B(_05211_),
    .Y(_05575_));
 sky130_fd_sc_hd__nor2_4 _20196_ (.A(_05242_),
    .B(_05204_),
    .Y(_05576_));
 sky130_fd_sc_hd__a22o_1 _20197_ (.A1(_05575_),
    .A2(\line_cache[108][0] ),
    .B1(_05576_),
    .B2(\line_cache[107][0] ),
    .X(_05577_));
 sky130_fd_sc_hd__a221o_1 _20198_ (.A1(\line_cache[110][0] ),
    .A2(_05573_),
    .B1(\line_cache[109][0] ),
    .B2(_05574_),
    .C1(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__nor2_2 _20199_ (.A(_05246_),
    .B(_05232_),
    .Y(_05579_));
 sky130_fd_sc_hd__nor2_4 _20200_ (.A(_05242_),
    .B(_05455_),
    .Y(_05580_));
 sky130_fd_sc_hd__nor2_2 _20201_ (.A(_05246_),
    .B(_05383_),
    .Y(_05581_));
 sky130_fd_sc_hd__nor2_2 _20202_ (.A(_05246_),
    .B(_05385_),
    .Y(_05582_));
 sky130_fd_sc_hd__a22o_1 _20203_ (.A1(_05581_),
    .A2(\line_cache[113][0] ),
    .B1(\line_cache[114][0] ),
    .B2(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__a221o_1 _20204_ (.A1(\line_cache[112][0] ),
    .A2(_05579_),
    .B1(\line_cache[111][0] ),
    .B2(_05580_),
    .C1(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__or4_1 _20205_ (.A(_05565_),
    .B(_05572_),
    .C(_05578_),
    .D(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_8 _20206_ (.A(_05215_),
    .X(_05586_));
 sky130_fd_sc_hd__nand2_1 _20207_ (.A(_05586_),
    .B(_05562_),
    .Y(_05587_));
 sky130_fd_sc_hd__inv_2 _20208_ (.A(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__nor2_2 _20209_ (.A(_05246_),
    .B(_05213_),
    .Y(_05589_));
 sky130_fd_sc_hd__nor2_4 _20210_ (.A(_05246_),
    .B(_05211_),
    .Y(_05590_));
 sky130_fd_sc_hd__nor2_4 _20211_ (.A(_05246_),
    .B(_05204_),
    .Y(_05591_));
 sky130_fd_sc_hd__a22o_1 _20212_ (.A1(_05590_),
    .A2(\line_cache[124][0] ),
    .B1(_05591_),
    .B2(\line_cache[123][0] ),
    .X(_05592_));
 sky130_fd_sc_hd__a221o_1 _20213_ (.A1(\line_cache[126][0] ),
    .A2(_05588_),
    .B1(\line_cache[125][0] ),
    .B2(_05589_),
    .C1(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__nor2_4 _20214_ (.A(_05253_),
    .B(_05232_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_1 _20215_ (.A(_05454_),
    .B(_05562_),
    .Y(_05595_));
 sky130_fd_sc_hd__inv_2 _20216_ (.A(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__nor2_2 _20217_ (.A(_05253_),
    .B(_05383_),
    .Y(_05597_));
 sky130_fd_sc_hd__nor2_4 _20218_ (.A(_05253_),
    .B(_05385_),
    .Y(_05598_));
 sky130_fd_sc_hd__and2_1 _20219_ (.A(_05598_),
    .B(\line_cache[130][0] ),
    .X(_05599_));
 sky130_fd_sc_hd__a21o_1 _20220_ (.A1(\line_cache[129][0] ),
    .A2(_05597_),
    .B1(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__a221o_1 _20221_ (.A1(\line_cache[128][0] ),
    .A2(_05594_),
    .B1(\line_cache[127][0] ),
    .B2(_05596_),
    .C1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__nor2_2 _20222_ (.A(_05253_),
    .B(_05201_),
    .Y(_05602_));
 sky130_fd_sc_hd__nor2_2 _20223_ (.A(_05253_),
    .B(_05208_),
    .Y(_05603_));
 sky130_fd_sc_hd__nor2_4 _20224_ (.A(_05253_),
    .B(_05396_),
    .Y(_05604_));
 sky130_fd_sc_hd__nor2_4 _20225_ (.A(_05253_),
    .B(_05228_),
    .Y(_05605_));
 sky130_fd_sc_hd__a22o_1 _20226_ (.A1(_05604_),
    .A2(\line_cache[136][0] ),
    .B1(_05605_),
    .B2(\line_cache[135][0] ),
    .X(_05606_));
 sky130_fd_sc_hd__a221o_1 _20227_ (.A1(\line_cache[138][0] ),
    .A2(_05602_),
    .B1(\line_cache[137][0] ),
    .B2(_05603_),
    .C1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__nor2_4 _20228_ (.A(_05253_),
    .B(_05389_),
    .Y(_05608_));
 sky130_fd_sc_hd__nor2_2 _20229_ (.A(_05253_),
    .B(_05225_),
    .Y(_05609_));
 sky130_fd_sc_hd__inv_6 _20230_ (.A(_05223_),
    .Y(_05610_));
 sky130_fd_sc_hd__buf_8 _20231_ (.A(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__nor2_2 _20232_ (.A(_05253_),
    .B(_05234_),
    .Y(_05612_));
 sky130_fd_sc_hd__a32o_1 _20233_ (.A1(_05611_),
    .A2(\line_cache[132][0] ),
    .A3(_05381_),
    .B1(\line_cache[131][0] ),
    .B2(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__a221o_1 _20234_ (.A1(\line_cache[134][0] ),
    .A2(_05608_),
    .B1(\line_cache[133][0] ),
    .B2(_05609_),
    .C1(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__or4_1 _20235_ (.A(_05593_),
    .B(_05601_),
    .C(_05607_),
    .D(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__nor2_1 _20236_ (.A(_05585_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__and4_2 _20237_ (.A(_05437_),
    .B(_05501_),
    .C(_05558_),
    .D(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__a22o_1 _20238_ (.A1(_05056_),
    .A2(\line_cache[301][0] ),
    .B1(\line_cache[300][0] ),
    .B2(_05053_),
    .X(_05618_));
 sky130_fd_sc_hd__a22o_1 _20239_ (.A1(_05073_),
    .A2(\line_cache[299][0] ),
    .B1(\line_cache[298][0] ),
    .B2(_05079_),
    .X(_05619_));
 sky130_fd_sc_hd__a22o_1 _20240_ (.A1(_05046_),
    .A2(\line_cache[295][0] ),
    .B1(\line_cache[294][0] ),
    .B2(_05043_),
    .X(_05620_));
 sky130_fd_sc_hd__a22o_1 _20241_ (.A1(_05069_),
    .A2(\line_cache[296][0] ),
    .B1(\line_cache[297][0] ),
    .B2(_05076_),
    .X(_05621_));
 sky130_fd_sc_hd__or4_1 _20242_ (.A(_05618_),
    .B(_05619_),
    .C(_05620_),
    .D(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__inv_2 _20243_ (.A(_05027_),
    .Y(_05623_));
 sky130_fd_sc_hd__inv_2 _20244_ (.A(_05022_),
    .Y(_05624_));
 sky130_fd_sc_hd__a22o_1 _20245_ (.A1(_05623_),
    .A2(\line_cache[291][0] ),
    .B1(\line_cache[290][0] ),
    .B2(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__inv_2 _20246_ (.A(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__inv_2 _20247_ (.A(_05039_),
    .Y(_05627_));
 sky130_fd_sc_hd__inv_2 _20248_ (.A(_05035_),
    .Y(_05628_));
 sky130_fd_sc_hd__a22oi_1 _20249_ (.A1(_05627_),
    .A2(\line_cache[292][0] ),
    .B1(\line_cache[293][0] ),
    .B2(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__clkinv_4 _20250_ (.A(_05177_),
    .Y(_05630_));
 sky130_fd_sc_hd__inv_2 _20251_ (.A(_05174_),
    .Y(_05631_));
 sky130_fd_sc_hd__inv_2 _20252_ (.A(_05011_),
    .Y(_05632_));
 sky130_fd_sc_hd__inv_2 _20253_ (.A(_05015_),
    .Y(_05633_));
 sky130_fd_sc_hd__a22o_1 _20254_ (.A1(_05632_),
    .A2(\line_cache[288][0] ),
    .B1(\line_cache[289][0] ),
    .B2(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__a221oi_4 _20255_ (.A1(\line_cache[286][0] ),
    .A2(_05630_),
    .B1(\line_cache[285][0] ),
    .B2(_05631_),
    .C1(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__and4b_1 _20256_ (.A_N(_05622_),
    .B(_05626_),
    .C(_05629_),
    .D(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__a22o_1 _20257_ (.A1(_05098_),
    .A2(\line_cache[308][0] ),
    .B1(\line_cache[307][0] ),
    .B2(_05136_),
    .X(_05637_));
 sky130_fd_sc_hd__a221oi_1 _20258_ (.A1(\line_cache[309][0] ),
    .A2(_05093_),
    .B1(\line_cache[310][0] ),
    .B2(_05103_),
    .C1(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__or2b_1 _20259_ (.A(_05060_),
    .B_N(\line_cache[302][0] ),
    .X(_05639_));
 sky130_fd_sc_hd__nand2_1 _20260_ (.A(_05129_),
    .B(\line_cache[304][0] ),
    .Y(_05640_));
 sky130_fd_sc_hd__nand2_1 _20261_ (.A(_05639_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__a221oi_1 _20262_ (.A1(\line_cache[306][0] ),
    .A2(_05132_),
    .B1(\line_cache[305][0] ),
    .B2(_05127_),
    .C1(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__nand2_1 _20263_ (.A(_05117_),
    .B(_05021_),
    .Y(_05643_));
 sky130_fd_sc_hd__inv_2 _20264_ (.A(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__or2b_1 _20265_ (.A(_05110_),
    .B_N(\line_cache[318][0] ),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_1 _20266_ (.A(_05106_),
    .B(\line_cache[317][0] ),
    .Y(_05646_));
 sky130_fd_sc_hd__nand2_1 _20267_ (.A(_05645_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__a221oi_4 _20268_ (.A1(\line_cache[316][0] ),
    .A2(_05108_),
    .B1(\line_cache[315][0] ),
    .B2(_05644_),
    .C1(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__nand2_1 _20269_ (.A(_05123_),
    .B(\line_cache[314][0] ),
    .Y(_05649_));
 sky130_fd_sc_hd__nand2_1 _20270_ (.A(_05121_),
    .B(\line_cache[313][0] ),
    .Y(_05650_));
 sky130_fd_sc_hd__nand2_1 _20271_ (.A(_05649_),
    .B(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__a221oi_1 _20272_ (.A1(_05119_),
    .A2(\line_cache[312][0] ),
    .B1(_05097_),
    .B2(\line_cache[311][0] ),
    .C1(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__and4_1 _20273_ (.A(_05638_),
    .B(_05642_),
    .C(_05648_),
    .D(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__inv_2 _20274_ (.A(_05170_),
    .Y(_05654_));
 sky130_fd_sc_hd__inv_2 _20275_ (.A(_05164_),
    .Y(_05655_));
 sky130_fd_sc_hd__a32o_1 _20276_ (.A1(_05059_),
    .A2(_05165_),
    .A3(\line_cache[278][0] ),
    .B1(_05655_),
    .B2(\line_cache[277][0] ),
    .X(_05656_));
 sky130_fd_sc_hd__a221o_1 _20277_ (.A1(\line_cache[280][0] ),
    .A2(_05144_),
    .B1(\line_cache[279][0] ),
    .B2(_05654_),
    .C1(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__inv_2 _20278_ (.A(_05168_),
    .Y(_05658_));
 sky130_fd_sc_hd__inv_2 _20279_ (.A(_05157_),
    .Y(_05659_));
 sky130_fd_sc_hd__inv_2 _20280_ (.A(_05159_),
    .Y(_05660_));
 sky130_fd_sc_hd__nand2_1 _20281_ (.A(_05660_),
    .B(\line_cache[273][0] ),
    .Y(_05661_));
 sky130_fd_sc_hd__inv_2 _20282_ (.A(_05161_),
    .Y(_05662_));
 sky130_fd_sc_hd__nand2_1 _20283_ (.A(_05662_),
    .B(\line_cache[274][0] ),
    .Y(_05663_));
 sky130_fd_sc_hd__nand2_1 _20284_ (.A(_05661_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__a221oi_1 _20285_ (.A1(_05658_),
    .A2(\line_cache[276][0] ),
    .B1(\line_cache[275][0] ),
    .B2(_05659_),
    .C1(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__inv_2 _20286_ (.A(_05155_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_2 _20287_ (.A(_05362_),
    .B(_05020_),
    .Y(_05667_));
 sky130_fd_sc_hd__inv_2 _20288_ (.A(_05667_),
    .Y(_05668_));
 sky130_fd_sc_hd__nand2_2 _20289_ (.A(_05360_),
    .B(_05009_),
    .Y(_05669_));
 sky130_fd_sc_hd__inv_2 _20290_ (.A(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__a32o_1 _20291_ (.A1(_05113_),
    .A2(_05364_),
    .A3(\line_cache[268][0] ),
    .B1(_05670_),
    .B2(\line_cache[269][0] ),
    .X(_05671_));
 sky130_fd_sc_hd__a221oi_2 _20292_ (.A1(\line_cache[272][0] ),
    .A2(_05666_),
    .B1(\line_cache[270][0] ),
    .B2(_05668_),
    .C1(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__and3_1 _20293_ (.A(_05142_),
    .B(_05052_),
    .C(_05020_),
    .X(_05673_));
 sky130_fd_sc_hd__clkbuf_4 _20294_ (.A(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__and3_2 _20295_ (.A(_05142_),
    .B(_05071_),
    .C(_05020_),
    .X(_05675_));
 sky130_fd_sc_hd__buf_2 _20296_ (.A(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__inv_2 _20297_ (.A(_05147_),
    .Y(_05677_));
 sky130_fd_sc_hd__inv_2 _20298_ (.A(_05149_),
    .Y(_05678_));
 sky130_fd_sc_hd__a22o_1 _20299_ (.A1(_05677_),
    .A2(\line_cache[281][0] ),
    .B1(\line_cache[282][0] ),
    .B2(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__a221oi_2 _20300_ (.A1(\line_cache[284][0] ),
    .A2(_05674_),
    .B1(\line_cache[283][0] ),
    .B2(_05676_),
    .C1(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__and4b_1 _20301_ (.A_N(_05657_),
    .B(_05665_),
    .C(_05672_),
    .D(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__and3_1 _20302_ (.A(_05636_),
    .B(_05653_),
    .C(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__nor2_4 _20303_ (.A(_05196_),
    .B(_05213_),
    .Y(_05683_));
 sky130_fd_sc_hd__and3_1 _20304_ (.A(_05203_),
    .B(\line_cache[203][0] ),
    .C(_05471_),
    .X(_05684_));
 sky130_fd_sc_hd__buf_4 _20305_ (.A(_05471_),
    .X(_05685_));
 sky130_fd_sc_hd__and3_1 _20306_ (.A(_05586_),
    .B(\line_cache[206][0] ),
    .C(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__or2_2 _20307_ (.A(_05196_),
    .B(_05211_),
    .X(_05687_));
 sky130_fd_sc_hd__and2b_1 _20308_ (.A_N(_05687_),
    .B(\line_cache[204][0] ),
    .X(_05688_));
 sky130_fd_sc_hd__a2111o_1 _20309_ (.A1(\line_cache[205][0] ),
    .A2(_05683_),
    .B1(_05684_),
    .C1(_05686_),
    .D1(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__nor2_2 _20310_ (.A(_05195_),
    .B(_05201_),
    .Y(_05690_));
 sky130_fd_sc_hd__nor2_4 _20311_ (.A(_05195_),
    .B(_05208_),
    .Y(_05691_));
 sky130_fd_sc_hd__nor2_2 _20312_ (.A(_05195_),
    .B(_05396_),
    .Y(_05692_));
 sky130_fd_sc_hd__inv_2 _20313_ (.A(_05195_),
    .Y(_05693_));
 sky130_fd_sc_hd__buf_4 _20314_ (.A(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__and3_1 _20315_ (.A(_05227_),
    .B(\line_cache[215][0] ),
    .C(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__a21o_1 _20316_ (.A1(\line_cache[216][0] ),
    .A2(_05692_),
    .B1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__a221o_1 _20317_ (.A1(\line_cache[218][0] ),
    .A2(_05690_),
    .B1(\line_cache[217][0] ),
    .B2(_05691_),
    .C1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__nor2_2 _20318_ (.A(_05195_),
    .B(_05232_),
    .Y(_05698_));
 sky130_fd_sc_hd__and3_2 _20319_ (.A(_05471_),
    .B(_05186_),
    .C(_05061_),
    .X(_05699_));
 sky130_fd_sc_hd__nor2_2 _20320_ (.A(_05195_),
    .B(_05383_),
    .Y(_05700_));
 sky130_fd_sc_hd__nor2_2 _20321_ (.A(_05195_),
    .B(_05385_),
    .Y(_05701_));
 sky130_fd_sc_hd__a22o_1 _20322_ (.A1(_05700_),
    .A2(\line_cache[209][0] ),
    .B1(\line_cache[210][0] ),
    .B2(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__a221o_1 _20323_ (.A1(\line_cache[208][0] ),
    .A2(_05698_),
    .B1(\line_cache[207][0] ),
    .B2(_05699_),
    .C1(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__clkinv_4 _20324_ (.A(_05234_),
    .Y(_05704_));
 sky130_fd_sc_hd__and3_1 _20325_ (.A(_05704_),
    .B(\line_cache[211][0] ),
    .C(_05694_),
    .X(_05705_));
 sky130_fd_sc_hd__clkbuf_4 _20326_ (.A(_05693_),
    .X(_05706_));
 sky130_fd_sc_hd__and3_1 _20327_ (.A(_05611_),
    .B(\line_cache[212][0] ),
    .C(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__clkinv_4 _20328_ (.A(_05389_),
    .Y(_05708_));
 sky130_fd_sc_hd__and3_1 _20329_ (.A(_05708_),
    .B(\line_cache[214][0] ),
    .C(_05706_),
    .X(_05709_));
 sky130_fd_sc_hd__clkinv_4 _20330_ (.A(_05225_),
    .Y(_05710_));
 sky130_fd_sc_hd__and3_1 _20331_ (.A(_05710_),
    .B(\line_cache[213][0] ),
    .C(_05706_),
    .X(_05711_));
 sky130_fd_sc_hd__or4_1 _20332_ (.A(_05705_),
    .B(_05707_),
    .C(_05709_),
    .D(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__or4_2 _20333_ (.A(_05689_),
    .B(_05697_),
    .C(_05703_),
    .D(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__nor2_2 _20334_ (.A(_05195_),
    .B(_05216_),
    .Y(_05714_));
 sky130_fd_sc_hd__nor2_4 _20335_ (.A(_05195_),
    .B(_05213_),
    .Y(_05715_));
 sky130_fd_sc_hd__nor2_2 _20336_ (.A(_05195_),
    .B(_05211_),
    .Y(_05716_));
 sky130_fd_sc_hd__nor2_2 _20337_ (.A(_05195_),
    .B(_05204_),
    .Y(_05717_));
 sky130_fd_sc_hd__a22o_1 _20338_ (.A1(_05716_),
    .A2(\line_cache[220][0] ),
    .B1(_05717_),
    .B2(\line_cache[219][0] ),
    .X(_05718_));
 sky130_fd_sc_hd__a221o_1 _20339_ (.A1(\line_cache[222][0] ),
    .A2(_05714_),
    .B1(\line_cache[221][0] ),
    .B2(_05715_),
    .C1(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__and3_2 _20340_ (.A(_05694_),
    .B(_05186_),
    .C(_05061_),
    .X(_05720_));
 sky130_fd_sc_hd__buf_4 _20341_ (.A(_05192_),
    .X(_05721_));
 sky130_fd_sc_hd__and3_1 _20342_ (.A(_05470_),
    .B(\line_cache[225][0] ),
    .C(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__and3_1 _20343_ (.A(_05408_),
    .B(\line_cache[226][0] ),
    .C(_05194_),
    .X(_05723_));
 sky130_fd_sc_hd__and3_1 _20344_ (.A(_05475_),
    .B(\line_cache[224][0] ),
    .C(_05194_),
    .X(_05724_));
 sky130_fd_sc_hd__a2111o_1 _20345_ (.A1(\line_cache[223][0] ),
    .A2(_05720_),
    .B1(_05722_),
    .C1(_05723_),
    .D1(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__nor2_2 _20346_ (.A(_05191_),
    .B(_05201_),
    .Y(_05726_));
 sky130_fd_sc_hd__nor2_4 _20347_ (.A(_05191_),
    .B(_05208_),
    .Y(_05727_));
 sky130_fd_sc_hd__nor2_2 _20348_ (.A(_05191_),
    .B(_05396_),
    .Y(_05728_));
 sky130_fd_sc_hd__nor2_2 _20349_ (.A(_05191_),
    .B(_05228_),
    .Y(_05729_));
 sky130_fd_sc_hd__a22o_1 _20350_ (.A1(_05728_),
    .A2(\line_cache[232][0] ),
    .B1(_05729_),
    .B2(\line_cache[231][0] ),
    .X(_05730_));
 sky130_fd_sc_hd__a221o_1 _20351_ (.A1(\line_cache[234][0] ),
    .A2(_05726_),
    .B1(\line_cache[233][0] ),
    .B2(_05727_),
    .C1(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__buf_4 _20352_ (.A(_05192_),
    .X(_05732_));
 sky130_fd_sc_hd__and3_1 _20353_ (.A(_05704_),
    .B(\line_cache[227][0] ),
    .C(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__and3_1 _20354_ (.A(_05611_),
    .B(\line_cache[228][0] ),
    .C(_05732_),
    .X(_05734_));
 sky130_fd_sc_hd__and3_1 _20355_ (.A(_05708_),
    .B(\line_cache[230][0] ),
    .C(_05721_),
    .X(_05735_));
 sky130_fd_sc_hd__and3_1 _20356_ (.A(_05710_),
    .B(\line_cache[229][0] ),
    .C(_05194_),
    .X(_05736_));
 sky130_fd_sc_hd__or4_1 _20357_ (.A(_05733_),
    .B(_05734_),
    .C(_05735_),
    .D(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__or4_1 _20358_ (.A(_05719_),
    .B(_05725_),
    .C(_05731_),
    .D(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__nor2_1 _20359_ (.A(_05713_),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__and3_1 _20360_ (.A(_05454_),
    .B(\line_cache[239][0] ),
    .C(_05721_),
    .X(_05740_));
 sky130_fd_sc_hd__and3_1 _20361_ (.A(_05470_),
    .B(\line_cache[241][0] ),
    .C(_05206_),
    .X(_05741_));
 sky130_fd_sc_hd__and3_1 _20362_ (.A(_05408_),
    .B(\line_cache[242][0] ),
    .C(_05206_),
    .X(_05742_));
 sky130_fd_sc_hd__a2111o_1 _20363_ (.A1(_05233_),
    .A2(\line_cache[240][0] ),
    .B1(_05740_),
    .C1(_05741_),
    .D1(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__nor2_2 _20364_ (.A(_05191_),
    .B(_05216_),
    .Y(_05744_));
 sky130_fd_sc_hd__nor2_2 _20365_ (.A(_05191_),
    .B(_05213_),
    .Y(_05745_));
 sky130_fd_sc_hd__nor2_2 _20366_ (.A(_05191_),
    .B(_05211_),
    .Y(_05746_));
 sky130_fd_sc_hd__nor2_2 _20367_ (.A(_05191_),
    .B(_05204_),
    .Y(_05747_));
 sky130_fd_sc_hd__a22o_1 _20368_ (.A1(_05746_),
    .A2(\line_cache[236][0] ),
    .B1(_05747_),
    .B2(\line_cache[235][0] ),
    .X(_05748_));
 sky130_fd_sc_hd__a221o_1 _20369_ (.A1(\line_cache[238][0] ),
    .A2(_05744_),
    .B1(\line_cache[237][0] ),
    .B2(_05745_),
    .C1(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__nor2_2 _20370_ (.A(_05199_),
    .B(_05396_),
    .Y(_05750_));
 sky130_fd_sc_hd__a22o_1 _20371_ (.A1(_05750_),
    .A2(\line_cache[248][0] ),
    .B1(_05229_),
    .B2(\line_cache[247][0] ),
    .X(_05751_));
 sky130_fd_sc_hd__a221o_1 _20372_ (.A1(\line_cache[250][0] ),
    .A2(_05202_),
    .B1(\line_cache[249][0] ),
    .B2(_05209_),
    .C1(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__nor2_4 _20373_ (.A(_05199_),
    .B(_05389_),
    .Y(_05753_));
 sky130_fd_sc_hd__a22o_1 _20374_ (.A1(_05235_),
    .A2(\line_cache[243][0] ),
    .B1(_05224_),
    .B2(\line_cache[244][0] ),
    .X(_05754_));
 sky130_fd_sc_hd__a221o_1 _20375_ (.A1(\line_cache[246][0] ),
    .A2(_05753_),
    .B1(\line_cache[245][0] ),
    .B2(_05226_),
    .C1(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__or4_1 _20376_ (.A(_05743_),
    .B(_05749_),
    .C(_05752_),
    .D(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__and3_1 _20377_ (.A(_05586_),
    .B(\line_cache[254][0] ),
    .C(_05198_),
    .X(_05757_));
 sky130_fd_sc_hd__a21o_1 _20378_ (.A1(\line_cache[253][0] ),
    .A2(_05214_),
    .B1(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__a221o_1 _20379_ (.A1(\line_cache[252][0] ),
    .A2(_05212_),
    .B1(\line_cache[251][0] ),
    .B2(_05205_),
    .C1(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__and3_4 _20380_ (.A(_05085_),
    .B(_05010_),
    .C(_05078_),
    .X(_05760_));
 sky130_fd_sc_hd__and3_1 _20381_ (.A(_05356_),
    .B(_05176_),
    .C(\line_cache[267][0] ),
    .X(_05761_));
 sky130_fd_sc_hd__and3_1 _20382_ (.A(_05085_),
    .B(_05020_),
    .C(_05068_),
    .X(_05762_));
 sky130_fd_sc_hd__clkbuf_4 _20383_ (.A(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__and3_4 _20384_ (.A(_05085_),
    .B(_05010_),
    .C(_05075_),
    .X(_05764_));
 sky130_fd_sc_hd__a22o_1 _20385_ (.A1(_05763_),
    .A2(\line_cache[264][0] ),
    .B1(\line_cache[265][0] ),
    .B2(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__a211o_1 _20386_ (.A1(\line_cache[266][0] ),
    .A2(_05760_),
    .B1(_05761_),
    .C1(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__and3_1 _20387_ (.A(_05085_),
    .B(_05010_),
    .C(_05042_),
    .X(_05767_));
 sky130_fd_sc_hd__buf_2 _20388_ (.A(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__nand2_2 _20389_ (.A(_05344_),
    .B(_05176_),
    .Y(_05769_));
 sky130_fd_sc_hd__inv_2 _20390_ (.A(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__clkbuf_8 _20391_ (.A(_05341_),
    .X(_05771_));
 sky130_fd_sc_hd__and3_1 _20392_ (.A(_05085_),
    .B(_05020_),
    .C(_05031_),
    .X(_05772_));
 sky130_fd_sc_hd__buf_2 _20393_ (.A(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__a32o_1 _20394_ (.A1(_05771_),
    .A2(_05176_),
    .A3(\line_cache[260][0] ),
    .B1(_05773_),
    .B2(\line_cache[261][0] ),
    .X(_05774_));
 sky130_fd_sc_hd__a221o_1 _20395_ (.A1(\line_cache[262][0] ),
    .A2(_05768_),
    .B1(_05770_),
    .B2(\line_cache[263][0] ),
    .C1(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__and3_4 _20396_ (.A(_05085_),
    .B(_05010_),
    .C(_05125_),
    .X(_05776_));
 sky130_fd_sc_hd__nor2_2 _20397_ (.A(_05003_),
    .B(_05086_),
    .Y(_05777_));
 sky130_fd_sc_hd__nor2_8 _20398_ (.A(_05025_),
    .B(_05340_),
    .Y(_05778_));
 sky130_fd_sc_hd__nor2_8 _20399_ (.A(_05018_),
    .B(_05340_),
    .Y(_05779_));
 sky130_fd_sc_hd__and3_1 _20400_ (.A(_05779_),
    .B(_05021_),
    .C(\line_cache[258][0] ),
    .X(_05780_));
 sky130_fd_sc_hd__a31o_1 _20401_ (.A1(_05151_),
    .A2(\line_cache[259][0] ),
    .A3(_05778_),
    .B1(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__a221o_1 _20402_ (.A1(\line_cache[257][0] ),
    .A2(_05776_),
    .B1(\line_cache[256][0] ),
    .B2(_05777_),
    .C1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__or4_1 _20403_ (.A(_05759_),
    .B(_05766_),
    .C(_05775_),
    .D(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__nor2_1 _20404_ (.A(_05756_),
    .B(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__and3_2 _20405_ (.A(_05682_),
    .B(_05739_),
    .C(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__and3_1 _20406_ (.A(_05112_),
    .B(_05113_),
    .C(\line_cache[319][0] ),
    .X(_05786_));
 sky130_fd_sc_hd__inv_2 _20407_ (.A(_05064_),
    .Y(_05787_));
 sky130_fd_sc_hd__inv_6 _20408_ (.A(_05181_),
    .Y(_05788_));
 sky130_fd_sc_hd__a22o_1 _20409_ (.A1(_05787_),
    .A2(\line_cache[303][0] ),
    .B1(\line_cache[287][0] ),
    .B2(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _20410_ (.A(_05366_),
    .B(_05176_),
    .Y(_05790_));
 sky130_fd_sc_hd__inv_2 _20411_ (.A(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__buf_4 _20412_ (.A(_05186_),
    .X(_05792_));
 sky130_fd_sc_hd__and3_1 _20413_ (.A(_05111_),
    .B(_05792_),
    .C(\line_cache[63][0] ),
    .X(_05793_));
 sky130_fd_sc_hd__and3_1 _20414_ (.A(_05063_),
    .B(_05187_),
    .C(\line_cache[47][0] ),
    .X(_05794_));
 sky130_fd_sc_hd__and3_1 _20415_ (.A(_05180_),
    .B(_05187_),
    .C(\line_cache[31][0] ),
    .X(_05795_));
 sky130_fd_sc_hd__a2111o_1 _20416_ (.A1(_05791_),
    .A2(\line_cache[271][0] ),
    .B1(_05793_),
    .C1(_05794_),
    .D1(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__and3_2 _20417_ (.A(_05085_),
    .B(_05186_),
    .C(_05125_),
    .X(_05797_));
 sky130_fd_sc_hd__inv_2 _20418_ (.A(_05367_),
    .Y(_05798_));
 sky130_fd_sc_hd__and3_1 _20419_ (.A(_05779_),
    .B(_05187_),
    .C(\line_cache[2][0] ),
    .X(_05799_));
 sky130_fd_sc_hd__a221o_1 _20420_ (.A1(_05797_),
    .A2(\line_cache[1][0] ),
    .B1(_05798_),
    .B2(\line_cache[15][0] ),
    .C1(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__and3_1 _20421_ (.A(_05778_),
    .B(_05186_),
    .C(\line_cache[3][0] ),
    .X(_05801_));
 sky130_fd_sc_hd__a31o_1 _20422_ (.A1(_05187_),
    .A2(\line_cache[4][0] ),
    .A3(_05771_),
    .B1(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__a221o_1 _20423_ (.A1(_05343_),
    .A2(\line_cache[5][0] ),
    .B1(\line_cache[6][0] ),
    .B2(_05348_),
    .C1(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__or3_1 _20424_ (.A(_05796_),
    .B(_05800_),
    .C(_05803_),
    .X(_05804_));
 sky130_fd_sc_hd__a2111oi_2 _20425_ (.A1(\line_cache[255][0] ),
    .A2(_05220_),
    .B1(_05786_),
    .C1(_05789_),
    .D1(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__and2_1 _20426_ (.A(_05261_),
    .B(\line_cache[35][0] ),
    .X(_05806_));
 sky130_fd_sc_hd__a22o_1 _20427_ (.A1(_05262_),
    .A2(\line_cache[33][0] ),
    .B1(\line_cache[34][0] ),
    .B2(_05263_),
    .X(_05807_));
 sky130_fd_sc_hd__and2_1 _20428_ (.A(_05275_),
    .B(\line_cache[40][0] ),
    .X(_05808_));
 sky130_fd_sc_hd__a21o_1 _20429_ (.A1(\line_cache[39][0] ),
    .A2(_05268_),
    .B1(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__a221o_1 _20430_ (.A1(\line_cache[38][0] ),
    .A2(_05270_),
    .B1(\line_cache[37][0] ),
    .B2(_05272_),
    .C1(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__a2111oi_1 _20431_ (.A1(\line_cache[36][0] ),
    .A2(_05266_),
    .B1(_05806_),
    .C1(_05807_),
    .D1(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__buf_4 _20432_ (.A(_05186_),
    .X(_05812_));
 sky130_fd_sc_hd__and3_1 _20433_ (.A(_05178_),
    .B(_05812_),
    .C(\line_cache[28][0] ),
    .X(_05813_));
 sky130_fd_sc_hd__a31o_1 _20434_ (.A1(_05188_),
    .A2(\line_cache[29][0] ),
    .A3(_05173_),
    .B1(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__and3_1 _20435_ (.A(_05175_),
    .B(_05188_),
    .C(\line_cache[30][0] ),
    .X(_05815_));
 sky130_fd_sc_hd__nand2_1 _20436_ (.A(_05150_),
    .B(_05187_),
    .Y(_05816_));
 sky130_fd_sc_hd__inv_4 _20437_ (.A(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _20438_ (.A(_05148_),
    .B(_05187_),
    .Y(_05818_));
 sky130_fd_sc_hd__inv_4 _20439_ (.A(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__and3_1 _20440_ (.A(_05320_),
    .B(_05186_),
    .C(\line_cache[24][0] ),
    .X(_05820_));
 sky130_fd_sc_hd__and3_1 _20441_ (.A(_05146_),
    .B(_05186_),
    .C(\line_cache[25][0] ),
    .X(_05821_));
 sky130_fd_sc_hd__or2_1 _20442_ (.A(_05820_),
    .B(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__a221o_1 _20443_ (.A1(\line_cache[27][0] ),
    .A2(_05817_),
    .B1(\line_cache[26][0] ),
    .B2(_05819_),
    .C1(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__a2111oi_1 _20444_ (.A1(\line_cache[32][0] ),
    .A2(_05260_),
    .B1(_05814_),
    .C1(_05815_),
    .D1(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__inv_2 _20445_ (.A(_05323_),
    .Y(_05825_));
 sky130_fd_sc_hd__inv_2 _20446_ (.A(_05322_),
    .Y(_05826_));
 sky130_fd_sc_hd__and3_1 _20447_ (.A(_05163_),
    .B(_05186_),
    .C(\line_cache[21][0] ),
    .X(_05827_));
 sky130_fd_sc_hd__and3_1 _20448_ (.A(_05167_),
    .B(_05792_),
    .C(\line_cache[20][0] ),
    .X(_05828_));
 sky130_fd_sc_hd__or2_1 _20449_ (.A(_05827_),
    .B(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__a221o_1 _20450_ (.A1(\line_cache[23][0] ),
    .A2(_05825_),
    .B1(\line_cache[22][0] ),
    .B2(_05826_),
    .C1(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__inv_2 _20451_ (.A(_05326_),
    .Y(_05831_));
 sky130_fd_sc_hd__inv_2 _20452_ (.A(_05325_),
    .Y(_05832_));
 sky130_fd_sc_hd__a22o_1 _20453_ (.A1(_05329_),
    .A2(\line_cache[16][0] ),
    .B1(\line_cache[17][0] ),
    .B2(_05330_),
    .X(_05833_));
 sky130_fd_sc_hd__a221o_1 _20454_ (.A1(\line_cache[19][0] ),
    .A2(_05831_),
    .B1(\line_cache[18][0] ),
    .B2(_05832_),
    .C1(_05833_),
    .X(_05834_));
 sky130_fd_sc_hd__nor2_1 _20455_ (.A(_05830_),
    .B(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__a22o_1 _20456_ (.A1(_05351_),
    .A2(\line_cache[9][0] ),
    .B1(\line_cache[10][0] ),
    .B2(_05353_),
    .X(_05836_));
 sky130_fd_sc_hd__a221o_1 _20457_ (.A1(\line_cache[8][0] ),
    .A2(_05355_),
    .B1(\line_cache[7][0] ),
    .B2(_05346_),
    .C1(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__inv_2 _20458_ (.A(_05363_),
    .Y(_05838_));
 sky130_fd_sc_hd__inv_2 _20459_ (.A(_05361_),
    .Y(_05839_));
 sky130_fd_sc_hd__clkbuf_8 _20460_ (.A(_05187_),
    .X(_05840_));
 sky130_fd_sc_hd__a32o_1 _20461_ (.A1(_05840_),
    .A2(_05364_),
    .A3(\line_cache[12][0] ),
    .B1(_05358_),
    .B2(\line_cache[11][0] ),
    .X(_05841_));
 sky130_fd_sc_hd__a221o_1 _20462_ (.A1(\line_cache[14][0] ),
    .A2(_05838_),
    .B1(\line_cache[13][0] ),
    .B2(_05839_),
    .C1(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__nor2_1 _20463_ (.A(_05837_),
    .B(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__and4_2 _20464_ (.A(_05811_),
    .B(_05824_),
    .C(_05835_),
    .D(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__a22o_1 _20465_ (.A1(_05301_),
    .A2(\line_cache[50][0] ),
    .B1(\line_cache[51][0] ),
    .B2(_05302_),
    .X(_05845_));
 sky130_fd_sc_hd__a22o_1 _20466_ (.A1(_05304_),
    .A2(\line_cache[52][0] ),
    .B1(\line_cache[53][0] ),
    .B2(_05306_),
    .X(_05846_));
 sky130_fd_sc_hd__a22o_1 _20467_ (.A1(_05314_),
    .A2(\line_cache[56][0] ),
    .B1(\line_cache[57][0] ),
    .B2(_05315_),
    .X(_05847_));
 sky130_fd_sc_hd__a221o_1 _20468_ (.A1(\line_cache[55][0] ),
    .A2(_05309_),
    .B1(\line_cache[54][0] ),
    .B2(_05307_),
    .C1(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__or3_1 _20469_ (.A(_05845_),
    .B(_05846_),
    .C(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__a22o_1 _20470_ (.A1(_05283_),
    .A2(\line_cache[45][0] ),
    .B1(\line_cache[46][0] ),
    .B2(_05285_),
    .X(_05850_));
 sky130_fd_sc_hd__a22o_1 _20471_ (.A1(_05298_),
    .A2(\line_cache[48][0] ),
    .B1(\line_cache[49][0] ),
    .B2(_05300_),
    .X(_05851_));
 sky130_fd_sc_hd__and2_1 _20472_ (.A(_05287_),
    .B(\line_cache[44][0] ),
    .X(_05852_));
 sky130_fd_sc_hd__a21o_1 _20473_ (.A1(\line_cache[43][0] ),
    .A2(_05277_),
    .B1(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__a221o_1 _20474_ (.A1(\line_cache[42][0] ),
    .A2(_05281_),
    .B1(\line_cache[41][0] ),
    .B2(_05279_),
    .C1(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__or3_1 _20475_ (.A(_05850_),
    .B(_05851_),
    .C(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__nor2_1 _20476_ (.A(_05849_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__a22o_1 _20477_ (.A1(_05292_),
    .A2(\line_cache[61][0] ),
    .B1(\line_cache[60][0] ),
    .B2(_05294_),
    .X(_05857_));
 sky130_fd_sc_hd__nor2_4 _20478_ (.A(_05245_),
    .B(_05232_),
    .Y(_05858_));
 sky130_fd_sc_hd__a22oi_1 _20479_ (.A1(_05858_),
    .A2(\line_cache[64][0] ),
    .B1(_05296_),
    .B2(\line_cache[62][0] ),
    .Y(_05859_));
 sky130_fd_sc_hd__nor2_2 _20480_ (.A(_05245_),
    .B(_05383_),
    .Y(_05860_));
 sky130_fd_sc_hd__nor2_2 _20481_ (.A(_05245_),
    .B(_05385_),
    .Y(_05861_));
 sky130_fd_sc_hd__a22oi_1 _20482_ (.A1(_05860_),
    .A2(\line_cache[65][0] ),
    .B1(\line_cache[66][0] ),
    .B2(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__a22oi_1 _20483_ (.A1(_05312_),
    .A2(\line_cache[58][0] ),
    .B1(_05317_),
    .B2(\line_cache[59][0] ),
    .Y(_05863_));
 sky130_fd_sc_hd__and4b_1 _20484_ (.A_N(_05857_),
    .B(_05859_),
    .C(_05862_),
    .D(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__nor2_2 _20485_ (.A(_05245_),
    .B(_05201_),
    .Y(_05865_));
 sky130_fd_sc_hd__nor2_4 _20486_ (.A(_05245_),
    .B(_05208_),
    .Y(_05866_));
 sky130_fd_sc_hd__nor2_2 _20487_ (.A(_05245_),
    .B(_05396_),
    .Y(_05867_));
 sky130_fd_sc_hd__nor2_4 _20488_ (.A(_05245_),
    .B(_05228_),
    .Y(_05868_));
 sky130_fd_sc_hd__a22o_1 _20489_ (.A1(_05867_),
    .A2(\line_cache[72][0] ),
    .B1(_05868_),
    .B2(\line_cache[71][0] ),
    .X(_05869_));
 sky130_fd_sc_hd__a221oi_2 _20490_ (.A1(\line_cache[74][0] ),
    .A2(_05865_),
    .B1(\line_cache[73][0] ),
    .B2(_05866_),
    .C1(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__nor2_2 _20491_ (.A(_05245_),
    .B(_05389_),
    .Y(_05871_));
 sky130_fd_sc_hd__nor2_4 _20492_ (.A(_05245_),
    .B(_05225_),
    .Y(_05872_));
 sky130_fd_sc_hd__nor2_2 _20493_ (.A(_05245_),
    .B(_05223_),
    .Y(_05873_));
 sky130_fd_sc_hd__nand2_1 _20494_ (.A(_05873_),
    .B(\line_cache[68][0] ),
    .Y(_05874_));
 sky130_fd_sc_hd__nor2_4 _20495_ (.A(_05245_),
    .B(_05234_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand2_1 _20496_ (.A(_05875_),
    .B(\line_cache[67][0] ),
    .Y(_05876_));
 sky130_fd_sc_hd__nand2_1 _20497_ (.A(_05874_),
    .B(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__a221oi_1 _20498_ (.A1(_05871_),
    .A2(\line_cache[70][0] ),
    .B1(\line_cache[69][0] ),
    .B2(_05872_),
    .C1(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__and4_1 _20499_ (.A(_05856_),
    .B(_05864_),
    .C(_05870_),
    .D(_05878_),
    .X(_05879_));
 sky130_fd_sc_hd__and3_1 _20500_ (.A(_05805_),
    .B(_05844_),
    .C(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__nand3_1 _20501_ (.A(_05617_),
    .B(_05785_),
    .C(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__nor2_1 _20502_ (.A(_08723_),
    .B(_08614_),
    .Y(_05882_));
 sky130_fd_sc_hd__nand2_4 _20503_ (.A(_05882_),
    .B(net168),
    .Y(_05883_));
 sky130_fd_sc_hd__clkinv_4 _20504_ (.A(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__o21a_4 _20505_ (.A1(_05373_),
    .A2(_05881_),
    .B1(_05884_),
    .X(net126));
 sky130_fd_sc_hd__nor3b_1 _20506_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][1] ),
    .Y(_05885_));
 sky130_fd_sc_hd__and3_1 _20507_ (.A(_05203_),
    .B(\line_cache[203][1] ),
    .C(_05685_),
    .X(_05886_));
 sky130_fd_sc_hd__and3_1 _20508_ (.A(_05586_),
    .B(\line_cache[206][1] ),
    .C(_05685_),
    .X(_05887_));
 sky130_fd_sc_hd__and2b_1 _20509_ (.A_N(_05687_),
    .B(\line_cache[204][1] ),
    .X(_05888_));
 sky130_fd_sc_hd__a2111o_1 _20510_ (.A1(\line_cache[205][1] ),
    .A2(_05683_),
    .B1(_05886_),
    .C1(_05887_),
    .D1(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__a22o_1 _20511_ (.A1(_05484_),
    .A2(\line_cache[195][1] ),
    .B1(_05485_),
    .B2(\line_cache[196][1] ),
    .X(_05890_));
 sky130_fd_sc_hd__a221o_1 _20512_ (.A1(\line_cache[198][1] ),
    .A2(_05487_),
    .B1(\line_cache[197][1] ),
    .B2(_05489_),
    .C1(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__a22o_1 _20513_ (.A1(_05495_),
    .A2(\line_cache[200][1] ),
    .B1(_05493_),
    .B2(\line_cache[199][1] ),
    .X(_05892_));
 sky130_fd_sc_hd__a221o_1 _20514_ (.A1(\line_cache[202][1] ),
    .A2(_05492_),
    .B1(\line_cache[201][1] ),
    .B2(_05491_),
    .C1(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__and3_1 _20515_ (.A(_05470_),
    .B(\line_cache[193][1] ),
    .C(_05472_),
    .X(_05894_));
 sky130_fd_sc_hd__and3_1 _20516_ (.A(_05475_),
    .B(\line_cache[192][1] ),
    .C(_05472_),
    .X(_05895_));
 sky130_fd_sc_hd__and3_1 _20517_ (.A(_05409_),
    .B(\line_cache[194][1] ),
    .C(_05472_),
    .X(_05896_));
 sky130_fd_sc_hd__a2111o_1 _20518_ (.A1(_05630_),
    .A2(\line_cache[286][1] ),
    .B1(_05894_),
    .C1(_05895_),
    .D1(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__or4_1 _20519_ (.A(_05889_),
    .B(_05891_),
    .C(_05893_),
    .D(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__a22o_1 _20520_ (.A1(_05676_),
    .A2(\line_cache[283][1] ),
    .B1(_05678_),
    .B2(\line_cache[282][1] ),
    .X(_05899_));
 sky130_fd_sc_hd__a22o_1 _20521_ (.A1(_05674_),
    .A2(\line_cache[284][1] ),
    .B1(_05631_),
    .B2(\line_cache[285][1] ),
    .X(_05900_));
 sky130_fd_sc_hd__a32o_1 _20522_ (.A1(_05165_),
    .A2(_05151_),
    .A3(\line_cache[278][1] ),
    .B1(_05654_),
    .B2(\line_cache[279][1] ),
    .X(_05901_));
 sky130_fd_sc_hd__a221o_1 _20523_ (.A1(\line_cache[281][1] ),
    .A2(_05677_),
    .B1(\line_cache[280][1] ),
    .B2(_05144_),
    .C1(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__a22o_1 _20524_ (.A1(_05668_),
    .A2(\line_cache[270][1] ),
    .B1(\line_cache[269][1] ),
    .B2(_05670_),
    .X(_05903_));
 sky130_fd_sc_hd__a22o_1 _20525_ (.A1(_05659_),
    .A2(\line_cache[275][1] ),
    .B1(\line_cache[274][1] ),
    .B2(_05662_),
    .X(_05904_));
 sky130_fd_sc_hd__a22o_1 _20526_ (.A1(_05658_),
    .A2(\line_cache[276][1] ),
    .B1(\line_cache[277][1] ),
    .B2(_05655_),
    .X(_05905_));
 sky130_fd_sc_hd__a22o_1 _20527_ (.A1(_05666_),
    .A2(\line_cache[272][1] ),
    .B1(\line_cache[273][1] ),
    .B2(_05660_),
    .X(_05906_));
 sky130_fd_sc_hd__or4_1 _20528_ (.A(_05903_),
    .B(_05904_),
    .C(_05905_),
    .D(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__or4_1 _20529_ (.A(_05899_),
    .B(_05900_),
    .C(_05902_),
    .D(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__nor2_1 _20530_ (.A(_05898_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__and3_1 _20531_ (.A(_05058_),
    .B(_05059_),
    .C(\line_cache[302][1] ),
    .X(_05910_));
 sky130_fd_sc_hd__a22o_1 _20532_ (.A1(_05056_),
    .A2(\line_cache[301][1] ),
    .B1(\line_cache[300][1] ),
    .B2(_05053_),
    .X(_05911_));
 sky130_fd_sc_hd__a211o_1 _20533_ (.A1(\line_cache[256][1] ),
    .A2(_05777_),
    .B1(_05910_),
    .C1(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__and3_1 _20534_ (.A(_05779_),
    .B(_05176_),
    .C(\line_cache[258][1] ),
    .X(_05913_));
 sky130_fd_sc_hd__and3_1 _20535_ (.A(_05771_),
    .B(_05059_),
    .C(\line_cache[260][1] ),
    .X(_05914_));
 sky130_fd_sc_hd__and3_1 _20536_ (.A(_05778_),
    .B(_05059_),
    .C(\line_cache[259][1] ),
    .X(_05915_));
 sky130_fd_sc_hd__a2111o_1 _20537_ (.A1(\line_cache[257][1] ),
    .A2(_05776_),
    .B1(_05913_),
    .C1(_05914_),
    .D1(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__and3_1 _20538_ (.A(_05356_),
    .B(_05059_),
    .C(\line_cache[267][1] ),
    .X(_05917_));
 sky130_fd_sc_hd__a22o_1 _20539_ (.A1(_05760_),
    .A2(\line_cache[266][1] ),
    .B1(\line_cache[265][1] ),
    .B2(_05764_),
    .X(_05918_));
 sky130_fd_sc_hd__a311o_1 _20540_ (.A1(_05113_),
    .A2(\line_cache[268][1] ),
    .A3(_05364_),
    .B1(_05917_),
    .C1(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__nand2_1 _20541_ (.A(_05768_),
    .B(\line_cache[262][1] ),
    .Y(_05920_));
 sky130_fd_sc_hd__nand2_1 _20542_ (.A(_05773_),
    .B(\line_cache[261][1] ),
    .Y(_05921_));
 sky130_fd_sc_hd__nand2_1 _20543_ (.A(_05920_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__a221oi_2 _20544_ (.A1(_05763_),
    .A2(\line_cache[264][1] ),
    .B1(_05770_),
    .B2(\line_cache[263][1] ),
    .C1(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__or4b_1 _20545_ (.A(_05912_),
    .B(_05916_),
    .C(_05919_),
    .D_N(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__a22o_1 _20546_ (.A1(_05098_),
    .A2(\line_cache[308][1] ),
    .B1(\line_cache[309][1] ),
    .B2(_05093_),
    .X(_05925_));
 sky130_fd_sc_hd__a221o_1 _20547_ (.A1(\line_cache[311][1] ),
    .A2(_05097_),
    .B1(\line_cache[310][1] ),
    .B2(_05103_),
    .C1(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__a22o_1 _20548_ (.A1(_05046_),
    .A2(\line_cache[295][1] ),
    .B1(\line_cache[294][1] ),
    .B2(_05043_),
    .X(_05927_));
 sky130_fd_sc_hd__a221o_1 _20549_ (.A1(\line_cache[293][1] ),
    .A2(_05628_),
    .B1(\line_cache[292][1] ),
    .B2(_05627_),
    .C1(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__a22o_1 _20550_ (.A1(_05069_),
    .A2(\line_cache[296][1] ),
    .B1(\line_cache[297][1] ),
    .B2(_05076_),
    .X(_05929_));
 sky130_fd_sc_hd__a221o_1 _20551_ (.A1(\line_cache[299][1] ),
    .A2(_05073_),
    .B1(\line_cache[298][1] ),
    .B2(_05079_),
    .C1(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__a22o_1 _20552_ (.A1(_05632_),
    .A2(\line_cache[288][1] ),
    .B1(\line_cache[289][1] ),
    .B2(_05633_),
    .X(_05931_));
 sky130_fd_sc_hd__a221o_1 _20553_ (.A1(\line_cache[291][1] ),
    .A2(_05623_),
    .B1(\line_cache[290][1] ),
    .B2(_05624_),
    .C1(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__or4_2 _20554_ (.A(_05926_),
    .B(_05928_),
    .C(_05930_),
    .D(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__nor2_1 _20555_ (.A(_05924_),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__nand2_1 _20556_ (.A(_05909_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__and3_1 _20557_ (.A(_05454_),
    .B(\line_cache[239][1] ),
    .C(_05194_),
    .X(_05936_));
 sky130_fd_sc_hd__and3_1 _20558_ (.A(_05470_),
    .B(\line_cache[241][1] ),
    .C(_05206_),
    .X(_05937_));
 sky130_fd_sc_hd__and3_1 _20559_ (.A(_05409_),
    .B(\line_cache[242][1] ),
    .C(_05206_),
    .X(_05938_));
 sky130_fd_sc_hd__a2111o_1 _20560_ (.A1(_05233_),
    .A2(\line_cache[240][1] ),
    .B1(_05936_),
    .C1(_05937_),
    .D1(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__and2_1 _20561_ (.A(_05235_),
    .B(\line_cache[243][1] ),
    .X(_05940_));
 sky130_fd_sc_hd__a21o_1 _20562_ (.A1(\line_cache[244][1] ),
    .A2(_05224_),
    .B1(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__a221o_1 _20563_ (.A1(\line_cache[246][1] ),
    .A2(_05753_),
    .B1(\line_cache[245][1] ),
    .B2(_05226_),
    .C1(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__a22o_1 _20564_ (.A1(_05212_),
    .A2(\line_cache[252][1] ),
    .B1(_05205_),
    .B2(\line_cache[251][1] ),
    .X(_05943_));
 sky130_fd_sc_hd__a221o_1 _20565_ (.A1(\line_cache[254][1] ),
    .A2(_05217_),
    .B1(\line_cache[253][1] ),
    .B2(_05214_),
    .C1(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__a22o_1 _20566_ (.A1(_05750_),
    .A2(\line_cache[248][1] ),
    .B1(_05229_),
    .B2(\line_cache[247][1] ),
    .X(_05945_));
 sky130_fd_sc_hd__a221o_1 _20567_ (.A1(\line_cache[250][1] ),
    .A2(_05202_),
    .B1(\line_cache[249][1] ),
    .B2(_05209_),
    .C1(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__or4_1 _20568_ (.A(_05939_),
    .B(_05942_),
    .C(_05944_),
    .D(_05946_),
    .X(_05947_));
 sky130_fd_sc_hd__a22o_1 _20569_ (.A1(_05873_),
    .A2(\line_cache[68][1] ),
    .B1(_05872_),
    .B2(\line_cache[69][1] ),
    .X(_05948_));
 sky130_fd_sc_hd__a221o_1 _20570_ (.A1(\line_cache[71][1] ),
    .A2(_05868_),
    .B1(\line_cache[70][1] ),
    .B2(_05871_),
    .C1(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__and2_1 _20571_ (.A(_05860_),
    .B(\line_cache[65][1] ),
    .X(_05950_));
 sky130_fd_sc_hd__a21o_1 _20572_ (.A1(_05858_),
    .A2(\line_cache[64][1] ),
    .B1(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__a221o_1 _20573_ (.A1(\line_cache[67][1] ),
    .A2(_05875_),
    .B1(\line_cache[66][1] ),
    .B2(_05861_),
    .C1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__and3_1 _20574_ (.A(_05200_),
    .B(\line_cache[74][1] ),
    .C(_05536_),
    .X(_05953_));
 sky130_fd_sc_hd__a22o_1 _20575_ (.A1(_05867_),
    .A2(\line_cache[72][1] ),
    .B1(_05866_),
    .B2(\line_cache[73][1] ),
    .X(_05954_));
 sky130_fd_sc_hd__a32o_1 _20576_ (.A1(_05544_),
    .A2(\line_cache[77][1] ),
    .A3(_05536_),
    .B1(\line_cache[76][1] ),
    .B2(_05542_),
    .X(_05955_));
 sky130_fd_sc_hd__a221o_1 _20577_ (.A1(\line_cache[79][1] ),
    .A2(_05537_),
    .B1(\line_cache[78][1] ),
    .B2(_05545_),
    .C1(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__a2111oi_1 _20578_ (.A1(\line_cache[75][1] ),
    .A2(_05543_),
    .B1(_05953_),
    .C1(_05954_),
    .D1(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__or3b_2 _20579_ (.A(_05949_),
    .B(_05952_),
    .C_N(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__nor2_1 _20580_ (.A(_05947_),
    .B(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__a22o_1 _20581_ (.A1(_05746_),
    .A2(\line_cache[236][1] ),
    .B1(_05747_),
    .B2(\line_cache[235][1] ),
    .X(_05960_));
 sky130_fd_sc_hd__a221o_1 _20582_ (.A1(\line_cache[238][1] ),
    .A2(_05744_),
    .B1(\line_cache[237][1] ),
    .B2(_05745_),
    .C1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__and3_1 _20583_ (.A(_05470_),
    .B(\line_cache[225][1] ),
    .C(_05194_),
    .X(_05962_));
 sky130_fd_sc_hd__and3_1 _20584_ (.A(_05409_),
    .B(\line_cache[226][1] ),
    .C(_05194_),
    .X(_05963_));
 sky130_fd_sc_hd__and3_1 _20585_ (.A(_05475_),
    .B(\line_cache[224][1] ),
    .C(_05194_),
    .X(_05964_));
 sky130_fd_sc_hd__a2111o_1 _20586_ (.A1(\line_cache[223][1] ),
    .A2(_05720_),
    .B1(_05962_),
    .C1(_05963_),
    .D1(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__and3_1 _20587_ (.A(_05704_),
    .B(\line_cache[227][1] ),
    .C(_05721_),
    .X(_05966_));
 sky130_fd_sc_hd__and3_1 _20588_ (.A(_05611_),
    .B(\line_cache[228][1] ),
    .C(_05721_),
    .X(_05967_));
 sky130_fd_sc_hd__and3_1 _20589_ (.A(_05710_),
    .B(\line_cache[229][1] ),
    .C(_05721_),
    .X(_05968_));
 sky130_fd_sc_hd__and3_1 _20590_ (.A(_05708_),
    .B(\line_cache[230][1] ),
    .C(_05194_),
    .X(_05969_));
 sky130_fd_sc_hd__or4_1 _20591_ (.A(_05966_),
    .B(_05967_),
    .C(_05968_),
    .D(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__a22o_1 _20592_ (.A1(_05728_),
    .A2(\line_cache[232][1] ),
    .B1(_05729_),
    .B2(\line_cache[231][1] ),
    .X(_05971_));
 sky130_fd_sc_hd__a221o_1 _20593_ (.A1(\line_cache[234][1] ),
    .A2(_05726_),
    .B1(\line_cache[233][1] ),
    .B2(_05727_),
    .C1(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__or4_1 _20594_ (.A(_05961_),
    .B(_05965_),
    .C(_05970_),
    .D(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__a22o_1 _20595_ (.A1(_05716_),
    .A2(\line_cache[220][1] ),
    .B1(_05717_),
    .B2(\line_cache[219][1] ),
    .X(_05974_));
 sky130_fd_sc_hd__a221o_1 _20596_ (.A1(\line_cache[222][1] ),
    .A2(_05714_),
    .B1(\line_cache[221][1] ),
    .B2(_05715_),
    .C1(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__a22o_1 _20597_ (.A1(_05700_),
    .A2(\line_cache[209][1] ),
    .B1(\line_cache[210][1] ),
    .B2(_05701_),
    .X(_05976_));
 sky130_fd_sc_hd__a221o_1 _20598_ (.A1(\line_cache[208][1] ),
    .A2(_05698_),
    .B1(\line_cache[207][1] ),
    .B2(_05699_),
    .C1(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__and3_1 _20599_ (.A(_05704_),
    .B(\line_cache[211][1] ),
    .C(_05706_),
    .X(_05978_));
 sky130_fd_sc_hd__and3_1 _20600_ (.A(_05611_),
    .B(\line_cache[212][1] ),
    .C(_05706_),
    .X(_05979_));
 sky130_fd_sc_hd__and3_1 _20601_ (.A(_05710_),
    .B(\line_cache[213][1] ),
    .C(_05706_),
    .X(_05980_));
 sky130_fd_sc_hd__and3_1 _20602_ (.A(_05708_),
    .B(\line_cache[214][1] ),
    .C(_05706_),
    .X(_05981_));
 sky130_fd_sc_hd__or4_1 _20603_ (.A(_05978_),
    .B(_05979_),
    .C(_05980_),
    .D(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__nor2_2 _20604_ (.A(_05195_),
    .B(_05228_),
    .Y(_05983_));
 sky130_fd_sc_hd__a22o_1 _20605_ (.A1(_05692_),
    .A2(\line_cache[216][1] ),
    .B1(_05983_),
    .B2(\line_cache[215][1] ),
    .X(_05984_));
 sky130_fd_sc_hd__a221o_1 _20606_ (.A1(\line_cache[218][1] ),
    .A2(_05690_),
    .B1(\line_cache[217][1] ),
    .B2(_05691_),
    .C1(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__or4_2 _20607_ (.A(_05975_),
    .B(_05977_),
    .C(_05982_),
    .D(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__nor2_1 _20608_ (.A(_05973_),
    .B(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__nand2_1 _20609_ (.A(_05959_),
    .B(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__nor2_2 _20610_ (.A(_05935_),
    .B(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__and2_1 _20611_ (.A(_05797_),
    .B(\line_cache[1][1] ),
    .X(_05990_));
 sky130_fd_sc_hd__buf_4 _20612_ (.A(_05792_),
    .X(_05991_));
 sky130_fd_sc_hd__and3_1 _20613_ (.A(_05779_),
    .B(_05991_),
    .C(\line_cache[2][1] ),
    .X(_05992_));
 sky130_fd_sc_hd__a211o_1 _20614_ (.A1(\line_cache[15][1] ),
    .A2(_05798_),
    .B1(_05990_),
    .C1(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__and3_1 _20615_ (.A(_05778_),
    .B(_05792_),
    .C(\line_cache[3][1] ),
    .X(_05994_));
 sky130_fd_sc_hd__a31o_1 _20616_ (.A1(_05840_),
    .A2(\line_cache[4][1] ),
    .A3(_05771_),
    .B1(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__a221o_1 _20617_ (.A1(_05343_),
    .A2(\line_cache[5][1] ),
    .B1(\line_cache[6][1] ),
    .B2(_05348_),
    .C1(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__and3_1 _20618_ (.A(_05112_),
    .B(_05151_),
    .C(\line_cache[319][1] ),
    .X(_05997_));
 sky130_fd_sc_hd__inv_2 _20619_ (.A(_05288_),
    .Y(_05998_));
 sky130_fd_sc_hd__a32o_1 _20620_ (.A1(_05991_),
    .A2(_05180_),
    .A3(\line_cache[31][1] ),
    .B1(_05998_),
    .B2(\line_cache[47][1] ),
    .X(_05999_));
 sky130_fd_sc_hd__a311o_1 _20621_ (.A1(_05188_),
    .A2(\line_cache[63][1] ),
    .A3(_05112_),
    .B1(_05997_),
    .C1(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__nand2_1 _20622_ (.A(_05787_),
    .B(\line_cache[303][1] ),
    .Y(_06001_));
 sky130_fd_sc_hd__nand2_1 _20623_ (.A(_05791_),
    .B(\line_cache[271][1] ),
    .Y(_06002_));
 sky130_fd_sc_hd__nand2_1 _20624_ (.A(_06001_),
    .B(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__a221oi_4 _20625_ (.A1(\line_cache[255][1] ),
    .A2(_05220_),
    .B1(\line_cache[287][1] ),
    .B2(_05788_),
    .C1(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__or4b_1 _20626_ (.A(_05993_),
    .B(_05996_),
    .C(_06000_),
    .D_N(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__a22o_1 _20627_ (.A1(_05283_),
    .A2(\line_cache[45][1] ),
    .B1(\line_cache[46][1] ),
    .B2(_05285_),
    .X(_06006_));
 sky130_fd_sc_hd__a22o_1 _20628_ (.A1(_05298_),
    .A2(\line_cache[48][1] ),
    .B1(\line_cache[49][1] ),
    .B2(_05300_),
    .X(_06007_));
 sky130_fd_sc_hd__nand2_1 _20629_ (.A(_05279_),
    .B(\line_cache[41][1] ),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_1 _20630_ (.A(_05281_),
    .B(\line_cache[42][1] ),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2_1 _20631_ (.A(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__a221oi_1 _20632_ (.A1(_05277_),
    .A2(\line_cache[43][1] ),
    .B1(\line_cache[44][1] ),
    .B2(_05287_),
    .C1(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__or3b_1 _20633_ (.A(_06006_),
    .B(_06007_),
    .C_N(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__a22o_1 _20634_ (.A1(_05106_),
    .A2(\line_cache[317][1] ),
    .B1(\line_cache[316][1] ),
    .B2(_05108_),
    .X(_06013_));
 sky130_fd_sc_hd__a22o_1 _20635_ (.A1(_05292_),
    .A2(\line_cache[61][1] ),
    .B1(\line_cache[60][1] ),
    .B2(_05294_),
    .X(_06014_));
 sky130_fd_sc_hd__a22o_1 _20636_ (.A1(_05312_),
    .A2(\line_cache[58][1] ),
    .B1(_05317_),
    .B2(\line_cache[59][1] ),
    .X(_06015_));
 sky130_fd_sc_hd__and3_1 _20637_ (.A(_05109_),
    .B(_05021_),
    .C(\line_cache[318][1] ),
    .X(_06016_));
 sky130_fd_sc_hd__a21o_1 _20638_ (.A1(\line_cache[62][1] ),
    .A2(_05296_),
    .B1(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__or4_1 _20639_ (.A(_06013_),
    .B(_06014_),
    .C(_06015_),
    .D(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__a22o_1 _20640_ (.A1(_05129_),
    .A2(\line_cache[304][1] ),
    .B1(\line_cache[305][1] ),
    .B2(_05127_),
    .X(_06019_));
 sky130_fd_sc_hd__a22o_1 _20641_ (.A1(_05119_),
    .A2(\line_cache[312][1] ),
    .B1(\line_cache[313][1] ),
    .B2(_05121_),
    .X(_06020_));
 sky130_fd_sc_hd__a22o_1 _20642_ (.A1(_05123_),
    .A2(\line_cache[314][1] ),
    .B1(_05644_),
    .B2(\line_cache[315][1] ),
    .X(_06021_));
 sky130_fd_sc_hd__a22o_1 _20643_ (.A1(_05132_),
    .A2(\line_cache[306][1] ),
    .B1(\line_cache[307][1] ),
    .B2(_05136_),
    .X(_06022_));
 sky130_fd_sc_hd__or4_2 _20644_ (.A(_06019_),
    .B(_06020_),
    .C(_06021_),
    .D(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__a22o_1 _20645_ (.A1(_05314_),
    .A2(\line_cache[56][1] ),
    .B1(\line_cache[57][1] ),
    .B2(_05315_),
    .X(_06024_));
 sky130_fd_sc_hd__a22o_1 _20646_ (.A1(_05304_),
    .A2(\line_cache[52][1] ),
    .B1(\line_cache[53][1] ),
    .B2(_05306_),
    .X(_06025_));
 sky130_fd_sc_hd__a22o_1 _20647_ (.A1(_05301_),
    .A2(\line_cache[50][1] ),
    .B1(\line_cache[51][1] ),
    .B2(_05302_),
    .X(_06026_));
 sky130_fd_sc_hd__a22o_1 _20648_ (.A1(_05307_),
    .A2(\line_cache[54][1] ),
    .B1(_05309_),
    .B2(\line_cache[55][1] ),
    .X(_06027_));
 sky130_fd_sc_hd__or4_2 _20649_ (.A(_06024_),
    .B(_06025_),
    .C(_06026_),
    .D(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__or4_1 _20650_ (.A(_06012_),
    .B(_06018_),
    .C(_06023_),
    .D(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__or2b_1 _20651_ (.A(_05365_),
    .B_N(\line_cache[12][1] ),
    .X(_06030_));
 sky130_fd_sc_hd__nand2_1 _20652_ (.A(_05358_),
    .B(\line_cache[11][1] ),
    .Y(_06031_));
 sky130_fd_sc_hd__nand2_1 _20653_ (.A(_06030_),
    .B(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__a221oi_1 _20654_ (.A1(\line_cache[14][1] ),
    .A2(_05838_),
    .B1(\line_cache[13][1] ),
    .B2(_05839_),
    .C1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__nand2_1 _20655_ (.A(_05353_),
    .B(\line_cache[10][1] ),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _20656_ (.A(_05351_),
    .B(\line_cache[9][1] ),
    .Y(_06035_));
 sky130_fd_sc_hd__nand2_1 _20657_ (.A(_06034_),
    .B(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__a221oi_2 _20658_ (.A1(_05355_),
    .A2(\line_cache[8][1] ),
    .B1(_05346_),
    .B2(\line_cache[7][1] ),
    .C1(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__nand2_1 _20659_ (.A(_06033_),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__and3_1 _20660_ (.A(_05163_),
    .B(_05187_),
    .C(\line_cache[21][1] ),
    .X(_06039_));
 sky130_fd_sc_hd__and3_1 _20661_ (.A(_05167_),
    .B(_05812_),
    .C(\line_cache[20][1] ),
    .X(_06040_));
 sky130_fd_sc_hd__a22o_1 _20662_ (.A1(_05825_),
    .A2(\line_cache[23][1] ),
    .B1(\line_cache[22][1] ),
    .B2(_05826_),
    .X(_06041_));
 sky130_fd_sc_hd__a22o_1 _20663_ (.A1(_05329_),
    .A2(\line_cache[16][1] ),
    .B1(\line_cache[17][1] ),
    .B2(_05330_),
    .X(_06042_));
 sky130_fd_sc_hd__a221o_1 _20664_ (.A1(\line_cache[19][1] ),
    .A2(_05831_),
    .B1(\line_cache[18][1] ),
    .B2(_05832_),
    .C1(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__or4_2 _20665_ (.A(_06039_),
    .B(_06040_),
    .C(_06041_),
    .D(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__a22o_1 _20666_ (.A1(_05262_),
    .A2(\line_cache[33][1] ),
    .B1(\line_cache[34][1] ),
    .B2(_05263_),
    .X(_06045_));
 sky130_fd_sc_hd__a221o_1 _20667_ (.A1(\line_cache[36][1] ),
    .A2(_05266_),
    .B1(\line_cache[35][1] ),
    .B2(_05261_),
    .C1(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__and3_1 _20668_ (.A(_05146_),
    .B(_05792_),
    .C(\line_cache[25][1] ),
    .X(_06047_));
 sky130_fd_sc_hd__a31o_1 _20669_ (.A1(_05991_),
    .A2(\line_cache[24][1] ),
    .A3(_05320_),
    .B1(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__a221oi_4 _20670_ (.A1(\line_cache[27][1] ),
    .A2(_05817_),
    .B1(\line_cache[26][1] ),
    .B2(_05819_),
    .C1(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__a32o_1 _20671_ (.A1(_05175_),
    .A2(_05812_),
    .A3(\line_cache[30][1] ),
    .B1(_05260_),
    .B2(\line_cache[32][1] ),
    .X(_06050_));
 sky130_fd_sc_hd__inv_2 _20672_ (.A(_05335_),
    .Y(_06051_));
 sky130_fd_sc_hd__a32o_1 _20673_ (.A1(_05991_),
    .A2(_05173_),
    .A3(\line_cache[29][1] ),
    .B1(_06051_),
    .B2(\line_cache[28][1] ),
    .X(_06052_));
 sky130_fd_sc_hd__nor2_1 _20674_ (.A(_06050_),
    .B(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__nand2_1 _20675_ (.A(_05270_),
    .B(\line_cache[38][1] ),
    .Y(_06054_));
 sky130_fd_sc_hd__nand2_1 _20676_ (.A(_05272_),
    .B(\line_cache[37][1] ),
    .Y(_06055_));
 sky130_fd_sc_hd__nand2_1 _20677_ (.A(_06054_),
    .B(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__a221oi_1 _20678_ (.A1(_05268_),
    .A2(\line_cache[39][1] ),
    .B1(\line_cache[40][1] ),
    .B2(_05275_),
    .C1(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__and4b_1 _20679_ (.A_N(_06046_),
    .B(_06049_),
    .C(_06053_),
    .D(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__or3b_2 _20680_ (.A(_06038_),
    .B(_06044_),
    .C_N(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__nor3_2 _20681_ (.A(_06005_),
    .B(_06029_),
    .C(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__and3_1 _20682_ (.A(_05227_),
    .B(\line_cache[87][1] ),
    .C(_05518_),
    .X(_06061_));
 sky130_fd_sc_hd__a21o_1 _20683_ (.A1(\line_cache[86][1] ),
    .A2(_05529_),
    .B1(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__a221o_1 _20684_ (.A1(\line_cache[85][1] ),
    .A2(_05530_),
    .B1(\line_cache[84][1] ),
    .B2(_05532_),
    .C1(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__a22o_1 _20685_ (.A1(_05531_),
    .A2(\line_cache[83][1] ),
    .B1(_05539_),
    .B2(\line_cache[82][1] ),
    .X(_06064_));
 sky130_fd_sc_hd__a221o_1 _20686_ (.A1(\line_cache[81][1] ),
    .A2(_05538_),
    .B1(\line_cache[80][1] ),
    .B2(_05535_),
    .C1(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__a22o_1 _20687_ (.A1(_05524_),
    .A2(\line_cache[92][1] ),
    .B1(_05523_),
    .B2(\line_cache[93][1] ),
    .X(_06066_));
 sky130_fd_sc_hd__a221o_1 _20688_ (.A1(\line_cache[95][1] ),
    .A2(_05519_),
    .B1(\line_cache[94][1] ),
    .B2(_05522_),
    .C1(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__a22o_1 _20689_ (.A1(_05553_),
    .A2(\line_cache[88][1] ),
    .B1(_05549_),
    .B2(\line_cache[89][1] ),
    .X(_06068_));
 sky130_fd_sc_hd__a221o_1 _20690_ (.A1(\line_cache[91][1] ),
    .A2(_05525_),
    .B1(\line_cache[90][1] ),
    .B2(_05550_),
    .C1(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__or4_1 _20691_ (.A(_06063_),
    .B(_06065_),
    .C(_06067_),
    .D(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__a22o_1 _20692_ (.A1(_05510_),
    .A2(\line_cache[99][1] ),
    .B1(_05516_),
    .B2(\line_cache[98][1] ),
    .X(_06071_));
 sky130_fd_sc_hd__a221o_1 _20693_ (.A1(\line_cache[97][1] ),
    .A2(_05515_),
    .B1(\line_cache[96][1] ),
    .B2(_05520_),
    .C1(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__a22o_1 _20694_ (.A1(_05575_),
    .A2(\line_cache[108][1] ),
    .B1(_05574_),
    .B2(\line_cache[109][1] ),
    .X(_06073_));
 sky130_fd_sc_hd__a221o_1 _20695_ (.A1(\line_cache[111][1] ),
    .A2(_05580_),
    .B1(\line_cache[110][1] ),
    .B2(_05573_),
    .C1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__and2_1 _20696_ (.A(_05502_),
    .B(\line_cache[102][1] ),
    .X(_06075_));
 sky130_fd_sc_hd__a21o_1 _20697_ (.A1(\line_cache[103][1] ),
    .A2(_05504_),
    .B1(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__a221o_1 _20698_ (.A1(\line_cache[101][1] ),
    .A2(_05509_),
    .B1(\line_cache[100][1] ),
    .B2(_05511_),
    .C1(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__a22o_1 _20699_ (.A1(_05503_),
    .A2(\line_cache[104][1] ),
    .B1(_05508_),
    .B2(\line_cache[105][1] ),
    .X(_06078_));
 sky130_fd_sc_hd__a221o_1 _20700_ (.A1(\line_cache[107][1] ),
    .A2(_05576_),
    .B1(\line_cache[106][1] ),
    .B2(_05506_),
    .C1(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__or4_1 _20701_ (.A(_06072_),
    .B(_06074_),
    .C(_06077_),
    .D(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__nor2_1 _20702_ (.A(_06070_),
    .B(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__and3_1 _20703_ (.A(_05207_),
    .B(\line_cache[121][1] ),
    .C(_05562_),
    .X(_06082_));
 sky130_fd_sc_hd__a21o_1 _20704_ (.A1(\line_cache[120][1] ),
    .A2(_05561_),
    .B1(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__a221o_1 _20705_ (.A1(\line_cache[123][1] ),
    .A2(_05591_),
    .B1(\line_cache[122][1] ),
    .B2(_05559_),
    .C1(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__and3_1 _20706_ (.A(_05586_),
    .B(\line_cache[126][1] ),
    .C(_05562_),
    .X(_06085_));
 sky130_fd_sc_hd__a21o_1 _20707_ (.A1(\line_cache[127][1] ),
    .A2(_05596_),
    .B1(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__a221o_1 _20708_ (.A1(\line_cache[125][1] ),
    .A2(_05589_),
    .B1(\line_cache[124][1] ),
    .B2(_05590_),
    .C1(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__nor2_2 _20709_ (.A(_05246_),
    .B(_05228_),
    .Y(_06088_));
 sky130_fd_sc_hd__a22o_1 _20710_ (.A1(_05568_),
    .A2(\line_cache[116][1] ),
    .B1(_05567_),
    .B2(\line_cache[117][1] ),
    .X(_06089_));
 sky130_fd_sc_hd__a221o_1 _20711_ (.A1(\line_cache[119][1] ),
    .A2(_06088_),
    .B1(\line_cache[118][1] ),
    .B2(_05566_),
    .C1(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__a22o_1 _20712_ (.A1(_05569_),
    .A2(\line_cache[115][1] ),
    .B1(_05582_),
    .B2(\line_cache[114][1] ),
    .X(_06091_));
 sky130_fd_sc_hd__a221o_1 _20713_ (.A1(\line_cache[113][1] ),
    .A2(_05581_),
    .B1(\line_cache[112][1] ),
    .B2(_05579_),
    .C1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__or4_1 _20714_ (.A(_06084_),
    .B(_06087_),
    .C(_06090_),
    .D(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__and3_1 _20715_ (.A(_05207_),
    .B(\line_cache[137][1] ),
    .C(_05381_),
    .X(_06094_));
 sky130_fd_sc_hd__a21o_1 _20716_ (.A1(\line_cache[136][1] ),
    .A2(_05604_),
    .B1(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__a221o_1 _20717_ (.A1(\line_cache[139][1] ),
    .A2(_05377_),
    .B1(\line_cache[138][1] ),
    .B2(_05602_),
    .C1(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__a22o_1 _20718_ (.A1(_05376_),
    .A2(\line_cache[140][1] ),
    .B1(_05375_),
    .B2(\line_cache[141][1] ),
    .X(_06097_));
 sky130_fd_sc_hd__a221o_1 _20719_ (.A1(\line_cache[143][1] ),
    .A2(_05382_),
    .B1(\line_cache[142][1] ),
    .B2(_05374_),
    .C1(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__a22o_1 _20720_ (.A1(_05612_),
    .A2(\line_cache[131][1] ),
    .B1(_05598_),
    .B2(\line_cache[130][1] ),
    .X(_06099_));
 sky130_fd_sc_hd__a221o_1 _20721_ (.A1(\line_cache[129][1] ),
    .A2(_05597_),
    .B1(\line_cache[128][1] ),
    .B2(_05594_),
    .C1(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__and2_1 _20722_ (.A(_05609_),
    .B(\line_cache[133][1] ),
    .X(_06101_));
 sky130_fd_sc_hd__and3_1 _20723_ (.A(_05611_),
    .B(\line_cache[132][1] ),
    .C(_05381_),
    .X(_06102_));
 sky130_fd_sc_hd__or2_1 _20724_ (.A(_06101_),
    .B(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__a221o_1 _20725_ (.A1(\line_cache[135][1] ),
    .A2(_05605_),
    .B1(\line_cache[134][1] ),
    .B2(_05608_),
    .C1(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__or4_1 _20726_ (.A(_06096_),
    .B(_06098_),
    .C(_06100_),
    .D(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__nor2_1 _20727_ (.A(_06093_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__nor2_2 _20728_ (.A(_05252_),
    .B(_05201_),
    .Y(_06107_));
 sky130_fd_sc_hd__a22o_1 _20729_ (.A1(_05419_),
    .A2(\line_cache[155][1] ),
    .B1(\line_cache[154][1] ),
    .B2(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__a221o_1 _20730_ (.A1(\line_cache[153][1] ),
    .A2(_05399_),
    .B1(\line_cache[152][1] ),
    .B2(_05397_),
    .C1(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__a22o_1 _20731_ (.A1(_05392_),
    .A2(\line_cache[147][1] ),
    .B1(_05386_),
    .B2(\line_cache[146][1] ),
    .X(_06110_));
 sky130_fd_sc_hd__a221oi_2 _20732_ (.A1(\line_cache[145][1] ),
    .A2(_05384_),
    .B1(\line_cache[144][1] ),
    .B2(_05380_),
    .C1(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__a22o_1 _20733_ (.A1(_05393_),
    .A2(\line_cache[148][1] ),
    .B1(\line_cache[149][1] ),
    .B2(_05391_),
    .X(_06112_));
 sky130_fd_sc_hd__a221oi_2 _20734_ (.A1(\line_cache[151][1] ),
    .A2(_05398_),
    .B1(\line_cache[150][1] ),
    .B2(_05390_),
    .C1(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__a22o_1 _20735_ (.A1(_05418_),
    .A2(\line_cache[156][1] ),
    .B1(_05417_),
    .B2(\line_cache[157][1] ),
    .X(_06114_));
 sky130_fd_sc_hd__a221oi_1 _20736_ (.A1(\line_cache[159][1] ),
    .A2(_05413_),
    .B1(\line_cache[158][1] ),
    .B2(_05416_),
    .C1(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__and4b_1 _20737_ (.A_N(_06109_),
    .B(_06111_),
    .C(_06113_),
    .D(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__a22o_1 _20738_ (.A1(_05464_),
    .A2(\line_cache[171][1] ),
    .B1(\line_cache[170][1] ),
    .B2(_05424_),
    .X(_06117_));
 sky130_fd_sc_hd__a221o_1 _20739_ (.A1(\line_cache[169][1] ),
    .A2(_05423_),
    .B1(\line_cache[168][1] ),
    .B2(_05427_),
    .C1(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__a32o_1 _20740_ (.A1(_05409_),
    .A2(\line_cache[162][1] ),
    .A3(_05410_),
    .B1(\line_cache[163][1] ),
    .B2(_05433_),
    .X(_06119_));
 sky130_fd_sc_hd__a221oi_1 _20741_ (.A1(\line_cache[161][1] ),
    .A2(_05406_),
    .B1(\line_cache[160][1] ),
    .B2(_05414_),
    .C1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__a22o_1 _20742_ (.A1(_05434_),
    .A2(\line_cache[164][1] ),
    .B1(\line_cache[165][1] ),
    .B2(_05432_),
    .X(_06121_));
 sky130_fd_sc_hd__nand2_1 _20743_ (.A(_05431_),
    .B(\line_cache[166][1] ),
    .Y(_06122_));
 sky130_fd_sc_hd__nand2_1 _20744_ (.A(_05425_),
    .B(\line_cache[167][1] ),
    .Y(_06123_));
 sky130_fd_sc_hd__and3b_1 _20745_ (.A_N(_06121_),
    .B(_06122_),
    .C(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__nand2_1 _20746_ (.A(_05462_),
    .B(\line_cache[173][1] ),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_1 _20747_ (.A(_05463_),
    .B(\line_cache[172][1] ),
    .Y(_06126_));
 sky130_fd_sc_hd__nand2_1 _20748_ (.A(_06125_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__a221oi_2 _20749_ (.A1(_05461_),
    .A2(\line_cache[174][1] ),
    .B1(_05456_),
    .B2(\line_cache[175][1] ),
    .C1(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__and4b_1 _20750_ (.A_N(_06118_),
    .B(_06120_),
    .C(_06124_),
    .D(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__nand2_1 _20751_ (.A(_05200_),
    .B(_05441_),
    .Y(_06130_));
 sky130_fd_sc_hd__inv_2 _20752_ (.A(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__a22o_1 _20753_ (.A1(_05438_),
    .A2(\line_cache[184][1] ),
    .B1(_05440_),
    .B2(\line_cache[185][1] ),
    .X(_06132_));
 sky130_fd_sc_hd__a221o_1 _20754_ (.A1(\line_cache[187][1] ),
    .A2(_05481_),
    .B1(\line_cache[186][1] ),
    .B2(_06131_),
    .C1(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__a22o_1 _20755_ (.A1(_05449_),
    .A2(\line_cache[180][1] ),
    .B1(\line_cache[181][1] ),
    .B2(_05446_),
    .X(_06134_));
 sky130_fd_sc_hd__a221oi_1 _20756_ (.A1(\line_cache[183][1] ),
    .A2(_05439_),
    .B1(\line_cache[182][1] ),
    .B2(_05445_),
    .C1(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__a22o_1 _20757_ (.A1(_05447_),
    .A2(\line_cache[179][1] ),
    .B1(_05458_),
    .B2(\line_cache[178][1] ),
    .X(_06136_));
 sky130_fd_sc_hd__a221oi_1 _20758_ (.A1(\line_cache[177][1] ),
    .A2(_05457_),
    .B1(\line_cache[176][1] ),
    .B2(_05453_),
    .C1(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__a22o_1 _20759_ (.A1(_05480_),
    .A2(\line_cache[188][1] ),
    .B1(_05479_),
    .B2(\line_cache[189][1] ),
    .X(_06138_));
 sky130_fd_sc_hd__a221oi_2 _20760_ (.A1(\line_cache[191][1] ),
    .A2(_05468_),
    .B1(\line_cache[190][1] ),
    .B2(_05478_),
    .C1(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__and4b_1 _20761_ (.A_N(_06133_),
    .B(_06135_),
    .C(_06137_),
    .D(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__and3_1 _20762_ (.A(_06116_),
    .B(_06129_),
    .C(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__and3_2 _20763_ (.A(_06081_),
    .B(_06106_),
    .C(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__nand3_1 _20764_ (.A(_05989_),
    .B(_06060_),
    .C(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__o21a_4 _20765_ (.A1(_05885_),
    .A2(_06143_),
    .B1(_05884_),
    .X(net127));
 sky130_fd_sc_hd__nor3b_1 _20766_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][2] ),
    .Y(_06144_));
 sky130_fd_sc_hd__and2_1 _20767_ (.A(_05797_),
    .B(\line_cache[1][2] ),
    .X(_06145_));
 sky130_fd_sc_hd__and3_1 _20768_ (.A(_05779_),
    .B(_05840_),
    .C(\line_cache[2][2] ),
    .X(_06146_));
 sky130_fd_sc_hd__a211o_1 _20769_ (.A1(\line_cache[15][2] ),
    .A2(_05798_),
    .B1(_06145_),
    .C1(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__and3_1 _20770_ (.A(_05778_),
    .B(_05792_),
    .C(\line_cache[3][2] ),
    .X(_06148_));
 sky130_fd_sc_hd__a31o_1 _20771_ (.A1(_05188_),
    .A2(\line_cache[4][2] ),
    .A3(_05771_),
    .B1(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__a221o_1 _20772_ (.A1(_05343_),
    .A2(\line_cache[5][2] ),
    .B1(\line_cache[6][2] ),
    .B2(_05348_),
    .C1(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__and3_1 _20773_ (.A(_05112_),
    .B(_05151_),
    .C(\line_cache[319][2] ),
    .X(_06151_));
 sky130_fd_sc_hd__a32o_1 _20774_ (.A1(_05840_),
    .A2(_05180_),
    .A3(\line_cache[31][2] ),
    .B1(_05998_),
    .B2(\line_cache[47][2] ),
    .X(_06152_));
 sky130_fd_sc_hd__a311o_1 _20775_ (.A1(_05188_),
    .A2(\line_cache[63][2] ),
    .A3(_05112_),
    .B1(_06151_),
    .C1(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__nand2_1 _20776_ (.A(_05787_),
    .B(\line_cache[303][2] ),
    .Y(_06154_));
 sky130_fd_sc_hd__nand2_1 _20777_ (.A(_05791_),
    .B(\line_cache[271][2] ),
    .Y(_06155_));
 sky130_fd_sc_hd__nand2_1 _20778_ (.A(_06154_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__a221oi_2 _20779_ (.A1(\line_cache[255][2] ),
    .A2(_05220_),
    .B1(\line_cache[287][2] ),
    .B2(_05788_),
    .C1(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__or4b_1 _20780_ (.A(_06147_),
    .B(_06150_),
    .C(_06153_),
    .D_N(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__a22o_1 _20781_ (.A1(_05283_),
    .A2(\line_cache[45][2] ),
    .B1(\line_cache[46][2] ),
    .B2(_05285_),
    .X(_06159_));
 sky130_fd_sc_hd__a22o_1 _20782_ (.A1(_05298_),
    .A2(\line_cache[48][2] ),
    .B1(\line_cache[49][2] ),
    .B2(_05300_),
    .X(_06160_));
 sky130_fd_sc_hd__nand2_1 _20783_ (.A(_05279_),
    .B(\line_cache[41][2] ),
    .Y(_06161_));
 sky130_fd_sc_hd__nand2_1 _20784_ (.A(_05281_),
    .B(\line_cache[42][2] ),
    .Y(_06162_));
 sky130_fd_sc_hd__nand2_1 _20785_ (.A(_06161_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__a221oi_1 _20786_ (.A1(_05277_),
    .A2(\line_cache[43][2] ),
    .B1(\line_cache[44][2] ),
    .B2(_05287_),
    .C1(_06163_),
    .Y(_06164_));
 sky130_fd_sc_hd__or3b_2 _20787_ (.A(_06159_),
    .B(_06160_),
    .C_N(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__a22o_1 _20788_ (.A1(_05106_),
    .A2(\line_cache[317][2] ),
    .B1(\line_cache[316][2] ),
    .B2(_05108_),
    .X(_06166_));
 sky130_fd_sc_hd__a22o_1 _20789_ (.A1(_05292_),
    .A2(\line_cache[61][2] ),
    .B1(\line_cache[60][2] ),
    .B2(_05294_),
    .X(_06167_));
 sky130_fd_sc_hd__a22o_1 _20790_ (.A1(_05312_),
    .A2(\line_cache[58][2] ),
    .B1(_05317_),
    .B2(\line_cache[59][2] ),
    .X(_06168_));
 sky130_fd_sc_hd__and3_1 _20791_ (.A(_05109_),
    .B(_05021_),
    .C(\line_cache[318][2] ),
    .X(_06169_));
 sky130_fd_sc_hd__a21o_1 _20792_ (.A1(\line_cache[62][2] ),
    .A2(_05296_),
    .B1(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__or4_1 _20793_ (.A(_06166_),
    .B(_06167_),
    .C(_06168_),
    .D(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__a22o_1 _20794_ (.A1(_05129_),
    .A2(\line_cache[304][2] ),
    .B1(\line_cache[305][2] ),
    .B2(_05127_),
    .X(_06172_));
 sky130_fd_sc_hd__a22o_1 _20795_ (.A1(_05119_),
    .A2(\line_cache[312][2] ),
    .B1(\line_cache[313][2] ),
    .B2(_05121_),
    .X(_06173_));
 sky130_fd_sc_hd__a22o_1 _20796_ (.A1(_05123_),
    .A2(\line_cache[314][2] ),
    .B1(_05644_),
    .B2(\line_cache[315][2] ),
    .X(_06174_));
 sky130_fd_sc_hd__a22o_1 _20797_ (.A1(_05132_),
    .A2(\line_cache[306][2] ),
    .B1(\line_cache[307][2] ),
    .B2(_05136_),
    .X(_06175_));
 sky130_fd_sc_hd__or4_2 _20798_ (.A(_06172_),
    .B(_06173_),
    .C(_06174_),
    .D(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__a22o_1 _20799_ (.A1(_05314_),
    .A2(\line_cache[56][2] ),
    .B1(\line_cache[57][2] ),
    .B2(_05315_),
    .X(_06177_));
 sky130_fd_sc_hd__a22o_1 _20800_ (.A1(_05304_),
    .A2(\line_cache[52][2] ),
    .B1(\line_cache[53][2] ),
    .B2(_05306_),
    .X(_06178_));
 sky130_fd_sc_hd__a22o_1 _20801_ (.A1(_05301_),
    .A2(\line_cache[50][2] ),
    .B1(\line_cache[51][2] ),
    .B2(_05302_),
    .X(_06179_));
 sky130_fd_sc_hd__a22o_1 _20802_ (.A1(_05307_),
    .A2(\line_cache[54][2] ),
    .B1(_05309_),
    .B2(\line_cache[55][2] ),
    .X(_06180_));
 sky130_fd_sc_hd__or4_2 _20803_ (.A(_06177_),
    .B(_06178_),
    .C(_06179_),
    .D(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__or4_2 _20804_ (.A(_06165_),
    .B(_06171_),
    .C(_06176_),
    .D(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__or2b_1 _20805_ (.A(_05365_),
    .B_N(\line_cache[12][2] ),
    .X(_06183_));
 sky130_fd_sc_hd__nand2_1 _20806_ (.A(_05358_),
    .B(\line_cache[11][2] ),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _20807_ (.A(_06183_),
    .B(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__a221oi_1 _20808_ (.A1(\line_cache[14][2] ),
    .A2(_05838_),
    .B1(\line_cache[13][2] ),
    .B2(_05839_),
    .C1(_06185_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_1 _20809_ (.A(_05353_),
    .B(\line_cache[10][2] ),
    .Y(_06187_));
 sky130_fd_sc_hd__nand2_1 _20810_ (.A(_05351_),
    .B(\line_cache[9][2] ),
    .Y(_06188_));
 sky130_fd_sc_hd__nand2_1 _20811_ (.A(_06187_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__a221oi_2 _20812_ (.A1(_05355_),
    .A2(\line_cache[8][2] ),
    .B1(_05346_),
    .B2(\line_cache[7][2] ),
    .C1(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__nand2_1 _20813_ (.A(_06186_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__and3_1 _20814_ (.A(_05163_),
    .B(_05812_),
    .C(\line_cache[21][2] ),
    .X(_06192_));
 sky130_fd_sc_hd__and3_1 _20815_ (.A(_05167_),
    .B(_05812_),
    .C(\line_cache[20][2] ),
    .X(_06193_));
 sky130_fd_sc_hd__a22o_1 _20816_ (.A1(_05825_),
    .A2(\line_cache[23][2] ),
    .B1(\line_cache[22][2] ),
    .B2(_05826_),
    .X(_06194_));
 sky130_fd_sc_hd__a22o_1 _20817_ (.A1(_05329_),
    .A2(\line_cache[16][2] ),
    .B1(\line_cache[17][2] ),
    .B2(_05330_),
    .X(_06195_));
 sky130_fd_sc_hd__a221o_1 _20818_ (.A1(\line_cache[19][2] ),
    .A2(_05831_),
    .B1(\line_cache[18][2] ),
    .B2(_05832_),
    .C1(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__or4_1 _20819_ (.A(_06192_),
    .B(_06193_),
    .C(_06194_),
    .D(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__a22o_1 _20820_ (.A1(_05262_),
    .A2(\line_cache[33][2] ),
    .B1(\line_cache[34][2] ),
    .B2(_05263_),
    .X(_06198_));
 sky130_fd_sc_hd__a221o_1 _20821_ (.A1(\line_cache[36][2] ),
    .A2(_05266_),
    .B1(\line_cache[35][2] ),
    .B2(_05261_),
    .C1(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__and3_1 _20822_ (.A(_05146_),
    .B(_05792_),
    .C(\line_cache[25][2] ),
    .X(_06200_));
 sky130_fd_sc_hd__a31o_1 _20823_ (.A1(_05840_),
    .A2(\line_cache[24][2] ),
    .A3(_05320_),
    .B1(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__a221oi_4 _20824_ (.A1(\line_cache[27][2] ),
    .A2(_05817_),
    .B1(\line_cache[26][2] ),
    .B2(_05819_),
    .C1(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__a32o_1 _20825_ (.A1(_05175_),
    .A2(_05991_),
    .A3(\line_cache[30][2] ),
    .B1(_05260_),
    .B2(\line_cache[32][2] ),
    .X(_06203_));
 sky130_fd_sc_hd__a32o_1 _20826_ (.A1(_05188_),
    .A2(_05173_),
    .A3(\line_cache[29][2] ),
    .B1(_06051_),
    .B2(\line_cache[28][2] ),
    .X(_06204_));
 sky130_fd_sc_hd__nor2_1 _20827_ (.A(_06203_),
    .B(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__nand2_1 _20828_ (.A(_05270_),
    .B(\line_cache[38][2] ),
    .Y(_06206_));
 sky130_fd_sc_hd__nand2_1 _20829_ (.A(_05272_),
    .B(\line_cache[37][2] ),
    .Y(_06207_));
 sky130_fd_sc_hd__nand2_1 _20830_ (.A(_06206_),
    .B(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__a221oi_1 _20831_ (.A1(_05268_),
    .A2(\line_cache[39][2] ),
    .B1(\line_cache[40][2] ),
    .B2(_05275_),
    .C1(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__and4b_1 _20832_ (.A_N(_06199_),
    .B(_06202_),
    .C(_06205_),
    .D(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__or3b_2 _20833_ (.A(_06191_),
    .B(_06197_),
    .C_N(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__nor3_2 _20834_ (.A(_06158_),
    .B(_06182_),
    .C(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__and3_1 _20835_ (.A(_05058_),
    .B(_05176_),
    .C(\line_cache[302][2] ),
    .X(_06213_));
 sky130_fd_sc_hd__a22o_1 _20836_ (.A1(_05056_),
    .A2(\line_cache[301][2] ),
    .B1(\line_cache[300][2] ),
    .B2(_05053_),
    .X(_06214_));
 sky130_fd_sc_hd__a211o_1 _20837_ (.A1(\line_cache[256][2] ),
    .A2(_05777_),
    .B1(_06213_),
    .C1(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__and3_1 _20838_ (.A(_05779_),
    .B(_05034_),
    .C(\line_cache[258][2] ),
    .X(_06216_));
 sky130_fd_sc_hd__and3_1 _20839_ (.A(_05771_),
    .B(_05034_),
    .C(\line_cache[260][2] ),
    .X(_06217_));
 sky130_fd_sc_hd__and3_1 _20840_ (.A(_05778_),
    .B(_05176_),
    .C(\line_cache[259][2] ),
    .X(_06218_));
 sky130_fd_sc_hd__a2111o_1 _20841_ (.A1(\line_cache[257][2] ),
    .A2(_05776_),
    .B1(_06216_),
    .C1(_06217_),
    .D1(_06218_),
    .X(_06219_));
 sky130_fd_sc_hd__and3_1 _20842_ (.A(_05356_),
    .B(_05176_),
    .C(\line_cache[267][2] ),
    .X(_06220_));
 sky130_fd_sc_hd__a22o_1 _20843_ (.A1(_05760_),
    .A2(\line_cache[266][2] ),
    .B1(\line_cache[265][2] ),
    .B2(_05764_),
    .X(_06221_));
 sky130_fd_sc_hd__a311o_1 _20844_ (.A1(_05113_),
    .A2(\line_cache[268][2] ),
    .A3(_05364_),
    .B1(_06220_),
    .C1(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__nand2_1 _20845_ (.A(_05768_),
    .B(\line_cache[262][2] ),
    .Y(_06223_));
 sky130_fd_sc_hd__nand2_1 _20846_ (.A(_05773_),
    .B(\line_cache[261][2] ),
    .Y(_06224_));
 sky130_fd_sc_hd__nand2_1 _20847_ (.A(_06223_),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__a221oi_1 _20848_ (.A1(_05763_),
    .A2(\line_cache[264][2] ),
    .B1(_05770_),
    .B2(\line_cache[263][2] ),
    .C1(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__or4b_1 _20849_ (.A(_06215_),
    .B(_06219_),
    .C(_06222_),
    .D_N(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__a22o_1 _20850_ (.A1(_05098_),
    .A2(\line_cache[308][2] ),
    .B1(\line_cache[309][2] ),
    .B2(_05093_),
    .X(_06228_));
 sky130_fd_sc_hd__a221o_1 _20851_ (.A1(\line_cache[311][2] ),
    .A2(_05097_),
    .B1(\line_cache[310][2] ),
    .B2(_05103_),
    .C1(_06228_),
    .X(_06229_));
 sky130_fd_sc_hd__a22o_1 _20852_ (.A1(_05046_),
    .A2(\line_cache[295][2] ),
    .B1(\line_cache[294][2] ),
    .B2(_05043_),
    .X(_06230_));
 sky130_fd_sc_hd__a221o_1 _20853_ (.A1(\line_cache[293][2] ),
    .A2(_05628_),
    .B1(\line_cache[292][2] ),
    .B2(_05627_),
    .C1(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__a22o_1 _20854_ (.A1(_05069_),
    .A2(\line_cache[296][2] ),
    .B1(\line_cache[297][2] ),
    .B2(_05076_),
    .X(_06232_));
 sky130_fd_sc_hd__a221o_1 _20855_ (.A1(\line_cache[299][2] ),
    .A2(_05073_),
    .B1(\line_cache[298][2] ),
    .B2(_05079_),
    .C1(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__a22o_1 _20856_ (.A1(_05632_),
    .A2(\line_cache[288][2] ),
    .B1(\line_cache[289][2] ),
    .B2(_05633_),
    .X(_06234_));
 sky130_fd_sc_hd__a221o_1 _20857_ (.A1(\line_cache[291][2] ),
    .A2(_05623_),
    .B1(\line_cache[290][2] ),
    .B2(_05624_),
    .C1(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__or4_2 _20858_ (.A(_06229_),
    .B(_06231_),
    .C(_06233_),
    .D(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__nor2_1 _20859_ (.A(_06227_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__and3_1 _20860_ (.A(_05203_),
    .B(\line_cache[203][2] ),
    .C(_05471_),
    .X(_06238_));
 sky130_fd_sc_hd__and3_1 _20861_ (.A(_05586_),
    .B(\line_cache[206][2] ),
    .C(_05471_),
    .X(_06239_));
 sky130_fd_sc_hd__and2b_1 _20862_ (.A_N(_05687_),
    .B(\line_cache[204][2] ),
    .X(_06240_));
 sky130_fd_sc_hd__a2111o_1 _20863_ (.A1(\line_cache[205][2] ),
    .A2(_05683_),
    .B1(_06238_),
    .C1(_06239_),
    .D1(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__a22o_1 _20864_ (.A1(_05484_),
    .A2(\line_cache[195][2] ),
    .B1(_05485_),
    .B2(\line_cache[196][2] ),
    .X(_06242_));
 sky130_fd_sc_hd__a221o_1 _20865_ (.A1(\line_cache[198][2] ),
    .A2(_05487_),
    .B1(\line_cache[197][2] ),
    .B2(_05489_),
    .C1(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__a22o_1 _20866_ (.A1(_05495_),
    .A2(\line_cache[200][2] ),
    .B1(_05493_),
    .B2(\line_cache[199][2] ),
    .X(_06244_));
 sky130_fd_sc_hd__a221o_1 _20867_ (.A1(\line_cache[202][2] ),
    .A2(_05492_),
    .B1(\line_cache[201][2] ),
    .B2(_05491_),
    .C1(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__and3_1 _20868_ (.A(_05470_),
    .B(\line_cache[193][2] ),
    .C(_05685_),
    .X(_06246_));
 sky130_fd_sc_hd__and3_1 _20869_ (.A(_05475_),
    .B(\line_cache[192][2] ),
    .C(_05685_),
    .X(_06247_));
 sky130_fd_sc_hd__and3_1 _20870_ (.A(_05408_),
    .B(\line_cache[194][2] ),
    .C(_05472_),
    .X(_06248_));
 sky130_fd_sc_hd__a2111o_1 _20871_ (.A1(_05630_),
    .A2(\line_cache[286][2] ),
    .B1(_06246_),
    .C1(_06247_),
    .D1(_06248_),
    .X(_06249_));
 sky130_fd_sc_hd__or4_1 _20872_ (.A(_06241_),
    .B(_06243_),
    .C(_06245_),
    .D(_06249_),
    .X(_06250_));
 sky130_fd_sc_hd__a22o_1 _20873_ (.A1(_05659_),
    .A2(\line_cache[275][2] ),
    .B1(\line_cache[274][2] ),
    .B2(_05662_),
    .X(_06251_));
 sky130_fd_sc_hd__a22o_1 _20874_ (.A1(_05658_),
    .A2(\line_cache[276][2] ),
    .B1(\line_cache[277][2] ),
    .B2(_05655_),
    .X(_06252_));
 sky130_fd_sc_hd__a22o_1 _20875_ (.A1(_05668_),
    .A2(\line_cache[270][2] ),
    .B1(\line_cache[269][2] ),
    .B2(_05670_),
    .X(_06253_));
 sky130_fd_sc_hd__a221o_1 _20876_ (.A1(\line_cache[273][2] ),
    .A2(_05660_),
    .B1(\line_cache[272][2] ),
    .B2(_05666_),
    .C1(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__a22oi_1 _20877_ (.A1(_05676_),
    .A2(\line_cache[283][2] ),
    .B1(_05678_),
    .B2(\line_cache[282][2] ),
    .Y(_06255_));
 sky130_fd_sc_hd__a22oi_2 _20878_ (.A1(_05674_),
    .A2(\line_cache[284][2] ),
    .B1(_05631_),
    .B2(\line_cache[285][2] ),
    .Y(_06256_));
 sky130_fd_sc_hd__nand2_1 _20879_ (.A(_06255_),
    .B(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__a22o_1 _20880_ (.A1(_05144_),
    .A2(\line_cache[280][2] ),
    .B1(_05677_),
    .B2(\line_cache[281][2] ),
    .X(_06258_));
 sky130_fd_sc_hd__a32o_1 _20881_ (.A1(_05165_),
    .A2(_05151_),
    .A3(\line_cache[278][2] ),
    .B1(_05654_),
    .B2(\line_cache[279][2] ),
    .X(_06259_));
 sky130_fd_sc_hd__nor3_1 _20882_ (.A(_06257_),
    .B(_06258_),
    .C(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__or4b_2 _20883_ (.A(_06251_),
    .B(_06252_),
    .C(_06254_),
    .D_N(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__nor2_1 _20884_ (.A(_06250_),
    .B(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__a22o_1 _20885_ (.A1(_05746_),
    .A2(\line_cache[236][2] ),
    .B1(_05747_),
    .B2(\line_cache[235][2] ),
    .X(_06263_));
 sky130_fd_sc_hd__a221o_1 _20886_ (.A1(\line_cache[238][2] ),
    .A2(_05744_),
    .B1(\line_cache[237][2] ),
    .B2(_05745_),
    .C1(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__and3_1 _20887_ (.A(_05469_),
    .B(\line_cache[225][2] ),
    .C(_05732_),
    .X(_06265_));
 sky130_fd_sc_hd__and3_1 _20888_ (.A(_05408_),
    .B(\line_cache[226][2] ),
    .C(_05721_),
    .X(_06266_));
 sky130_fd_sc_hd__and3_1 _20889_ (.A(_05475_),
    .B(\line_cache[224][2] ),
    .C(_05721_),
    .X(_06267_));
 sky130_fd_sc_hd__a2111o_1 _20890_ (.A1(\line_cache[223][2] ),
    .A2(_05720_),
    .B1(_06265_),
    .C1(_06266_),
    .D1(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__and3_1 _20891_ (.A(_05704_),
    .B(\line_cache[227][2] ),
    .C(_05193_),
    .X(_06269_));
 sky130_fd_sc_hd__and3_1 _20892_ (.A(_05610_),
    .B(\line_cache[228][2] ),
    .C(_05193_),
    .X(_06270_));
 sky130_fd_sc_hd__and3_1 _20893_ (.A(_05710_),
    .B(\line_cache[229][2] ),
    .C(_05193_),
    .X(_06271_));
 sky130_fd_sc_hd__and3_1 _20894_ (.A(_05708_),
    .B(\line_cache[230][2] ),
    .C(_05732_),
    .X(_06272_));
 sky130_fd_sc_hd__or4_1 _20895_ (.A(_06269_),
    .B(_06270_),
    .C(_06271_),
    .D(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__a22o_1 _20896_ (.A1(_05728_),
    .A2(\line_cache[232][2] ),
    .B1(_05729_),
    .B2(\line_cache[231][2] ),
    .X(_06274_));
 sky130_fd_sc_hd__a221o_1 _20897_ (.A1(\line_cache[234][2] ),
    .A2(_05726_),
    .B1(\line_cache[233][2] ),
    .B2(_05727_),
    .C1(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__or4_1 _20898_ (.A(_06264_),
    .B(_06268_),
    .C(_06273_),
    .D(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__a22o_1 _20899_ (.A1(_05716_),
    .A2(\line_cache[220][2] ),
    .B1(_05717_),
    .B2(\line_cache[219][2] ),
    .X(_06277_));
 sky130_fd_sc_hd__a221o_1 _20900_ (.A1(\line_cache[222][2] ),
    .A2(_05714_),
    .B1(\line_cache[221][2] ),
    .B2(_05715_),
    .C1(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__a22o_1 _20901_ (.A1(_05700_),
    .A2(\line_cache[209][2] ),
    .B1(\line_cache[210][2] ),
    .B2(_05701_),
    .X(_06279_));
 sky130_fd_sc_hd__a221o_1 _20902_ (.A1(\line_cache[208][2] ),
    .A2(_05698_),
    .B1(\line_cache[207][2] ),
    .B2(_05699_),
    .C1(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__and3_1 _20903_ (.A(_05704_),
    .B(\line_cache[211][2] ),
    .C(_05694_),
    .X(_06281_));
 sky130_fd_sc_hd__and3_1 _20904_ (.A(_05611_),
    .B(\line_cache[212][2] ),
    .C(_05694_),
    .X(_06282_));
 sky130_fd_sc_hd__and3_1 _20905_ (.A(_05710_),
    .B(\line_cache[213][2] ),
    .C(_05694_),
    .X(_06283_));
 sky130_fd_sc_hd__and3_1 _20906_ (.A(_05708_),
    .B(\line_cache[214][2] ),
    .C(_05706_),
    .X(_06284_));
 sky130_fd_sc_hd__or4_2 _20907_ (.A(_06281_),
    .B(_06282_),
    .C(_06283_),
    .D(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__a22o_1 _20908_ (.A1(_05692_),
    .A2(\line_cache[216][2] ),
    .B1(_05983_),
    .B2(\line_cache[215][2] ),
    .X(_06286_));
 sky130_fd_sc_hd__a221o_1 _20909_ (.A1(\line_cache[218][2] ),
    .A2(_05690_),
    .B1(\line_cache[217][2] ),
    .B2(_05691_),
    .C1(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__or4_2 _20910_ (.A(_06278_),
    .B(_06280_),
    .C(_06285_),
    .D(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__nor2_1 _20911_ (.A(_06276_),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__and3_1 _20912_ (.A(_05454_),
    .B(\line_cache[239][2] ),
    .C(_05732_),
    .X(_06290_));
 sky130_fd_sc_hd__and3_1 _20913_ (.A(_05470_),
    .B(\line_cache[241][2] ),
    .C(_05206_),
    .X(_06291_));
 sky130_fd_sc_hd__and3_1 _20914_ (.A(_05408_),
    .B(\line_cache[242][2] ),
    .C(_05206_),
    .X(_06292_));
 sky130_fd_sc_hd__a2111o_1 _20915_ (.A1(_05233_),
    .A2(\line_cache[240][2] ),
    .B1(_06290_),
    .C1(_06291_),
    .D1(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__and2_1 _20916_ (.A(_05235_),
    .B(\line_cache[243][2] ),
    .X(_06294_));
 sky130_fd_sc_hd__a21o_1 _20917_ (.A1(\line_cache[244][2] ),
    .A2(_05224_),
    .B1(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__a221o_1 _20918_ (.A1(\line_cache[246][2] ),
    .A2(_05753_),
    .B1(\line_cache[245][2] ),
    .B2(_05226_),
    .C1(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__a22o_1 _20919_ (.A1(_05212_),
    .A2(\line_cache[252][2] ),
    .B1(_05205_),
    .B2(\line_cache[251][2] ),
    .X(_06297_));
 sky130_fd_sc_hd__a221o_1 _20920_ (.A1(\line_cache[254][2] ),
    .A2(_05217_),
    .B1(\line_cache[253][2] ),
    .B2(_05214_),
    .C1(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__a22o_1 _20921_ (.A1(_05750_),
    .A2(\line_cache[248][2] ),
    .B1(_05229_),
    .B2(\line_cache[247][2] ),
    .X(_06299_));
 sky130_fd_sc_hd__a221o_1 _20922_ (.A1(\line_cache[250][2] ),
    .A2(_05202_),
    .B1(\line_cache[249][2] ),
    .B2(_05209_),
    .C1(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__or4_1 _20923_ (.A(_06293_),
    .B(_06296_),
    .C(_06298_),
    .D(_06300_),
    .X(_06301_));
 sky130_fd_sc_hd__a22o_1 _20924_ (.A1(_05875_),
    .A2(\line_cache[67][2] ),
    .B1(_05861_),
    .B2(\line_cache[66][2] ),
    .X(_06302_));
 sky130_fd_sc_hd__a221o_1 _20925_ (.A1(\line_cache[65][2] ),
    .A2(_05860_),
    .B1(\line_cache[64][2] ),
    .B2(_05858_),
    .C1(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__a22o_1 _20926_ (.A1(_05867_),
    .A2(\line_cache[72][2] ),
    .B1(_05866_),
    .B2(\line_cache[73][2] ),
    .X(_06304_));
 sky130_fd_sc_hd__a221o_1 _20927_ (.A1(\line_cache[75][2] ),
    .A2(_05543_),
    .B1(\line_cache[74][2] ),
    .B2(_05865_),
    .C1(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__a22o_1 _20928_ (.A1(_05873_),
    .A2(\line_cache[68][2] ),
    .B1(_05872_),
    .B2(\line_cache[69][2] ),
    .X(_06306_));
 sky130_fd_sc_hd__a221o_1 _20929_ (.A1(\line_cache[71][2] ),
    .A2(_05868_),
    .B1(\line_cache[70][2] ),
    .B2(_05871_),
    .C1(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__and2_1 _20930_ (.A(_05542_),
    .B(\line_cache[76][2] ),
    .X(_06308_));
 sky130_fd_sc_hd__and3_1 _20931_ (.A(_05544_),
    .B(\line_cache[77][2] ),
    .C(_05536_),
    .X(_06309_));
 sky130_fd_sc_hd__or2_1 _20932_ (.A(_06308_),
    .B(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__a221o_1 _20933_ (.A1(\line_cache[79][2] ),
    .A2(_05537_),
    .B1(\line_cache[78][2] ),
    .B2(_05545_),
    .C1(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__or4_2 _20934_ (.A(_06303_),
    .B(_06305_),
    .C(_06307_),
    .D(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__nor2_1 _20935_ (.A(_06301_),
    .B(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__and4_1 _20936_ (.A(_06237_),
    .B(_06262_),
    .C(_06289_),
    .D(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__a22o_1 _20937_ (.A1(_05524_),
    .A2(\line_cache[92][2] ),
    .B1(_05523_),
    .B2(\line_cache[93][2] ),
    .X(_06315_));
 sky130_fd_sc_hd__a22o_1 _20938_ (.A1(_05522_),
    .A2(\line_cache[94][2] ),
    .B1(_05519_),
    .B2(\line_cache[95][2] ),
    .X(_06316_));
 sky130_fd_sc_hd__or2_1 _20939_ (.A(_06315_),
    .B(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__and3_1 _20940_ (.A(_05227_),
    .B(\line_cache[87][2] ),
    .C(_05518_),
    .X(_06318_));
 sky130_fd_sc_hd__a21o_1 _20941_ (.A1(\line_cache[86][2] ),
    .A2(_05529_),
    .B1(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__a221o_1 _20942_ (.A1(\line_cache[85][2] ),
    .A2(_05530_),
    .B1(\line_cache[84][2] ),
    .B2(_05532_),
    .C1(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__a22o_1 _20943_ (.A1(_05531_),
    .A2(\line_cache[83][2] ),
    .B1(_05539_),
    .B2(\line_cache[82][2] ),
    .X(_06321_));
 sky130_fd_sc_hd__a221o_2 _20944_ (.A1(\line_cache[81][2] ),
    .A2(_05538_),
    .B1(\line_cache[80][2] ),
    .B2(_05535_),
    .C1(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__a22o_1 _20945_ (.A1(_05553_),
    .A2(\line_cache[88][2] ),
    .B1(_05549_),
    .B2(\line_cache[89][2] ),
    .X(_06323_));
 sky130_fd_sc_hd__a221o_1 _20946_ (.A1(\line_cache[91][2] ),
    .A2(_05525_),
    .B1(\line_cache[90][2] ),
    .B2(_05550_),
    .C1(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__or4_1 _20947_ (.A(_06317_),
    .B(_06320_),
    .C(_06322_),
    .D(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__a22o_1 _20948_ (.A1(_05573_),
    .A2(\line_cache[110][2] ),
    .B1(_05580_),
    .B2(\line_cache[111][2] ),
    .X(_06326_));
 sky130_fd_sc_hd__a22o_1 _20949_ (.A1(_05575_),
    .A2(\line_cache[108][2] ),
    .B1(_05574_),
    .B2(\line_cache[109][2] ),
    .X(_06327_));
 sky130_fd_sc_hd__a22o_1 _20950_ (.A1(_05503_),
    .A2(\line_cache[104][2] ),
    .B1(_05508_),
    .B2(\line_cache[105][2] ),
    .X(_06328_));
 sky130_fd_sc_hd__a221o_1 _20951_ (.A1(\line_cache[107][2] ),
    .A2(_05576_),
    .B1(\line_cache[106][2] ),
    .B2(_05506_),
    .C1(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__a22o_1 _20952_ (.A1(\line_cache[97][2] ),
    .A2(_05515_),
    .B1(_05520_),
    .B2(\line_cache[96][2] ),
    .X(_06330_));
 sky130_fd_sc_hd__a22o_1 _20953_ (.A1(_05510_),
    .A2(\line_cache[99][2] ),
    .B1(_05516_),
    .B2(\line_cache[98][2] ),
    .X(_06331_));
 sky130_fd_sc_hd__and2_1 _20954_ (.A(_05502_),
    .B(\line_cache[102][2] ),
    .X(_06332_));
 sky130_fd_sc_hd__a21o_1 _20955_ (.A1(\line_cache[103][2] ),
    .A2(_05504_),
    .B1(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__a221o_1 _20956_ (.A1(\line_cache[101][2] ),
    .A2(_05509_),
    .B1(\line_cache[100][2] ),
    .B2(_05511_),
    .C1(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__or3_2 _20957_ (.A(_06330_),
    .B(_06331_),
    .C(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__or4_2 _20958_ (.A(_06326_),
    .B(_06327_),
    .C(_06329_),
    .D(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__nor2_1 _20959_ (.A(_06325_),
    .B(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__a22o_1 _20960_ (.A1(_05425_),
    .A2(\line_cache[167][2] ),
    .B1(\line_cache[166][2] ),
    .B2(_05431_),
    .X(_06338_));
 sky130_fd_sc_hd__a221o_1 _20961_ (.A1(\line_cache[165][2] ),
    .A2(_05432_),
    .B1(\line_cache[164][2] ),
    .B2(_05434_),
    .C1(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__a22o_1 _20962_ (.A1(\line_cache[161][2] ),
    .A2(_05406_),
    .B1(_05414_),
    .B2(\line_cache[160][2] ),
    .X(_06340_));
 sky130_fd_sc_hd__a32o_1 _20963_ (.A1(_05409_),
    .A2(\line_cache[162][2] ),
    .A3(_05410_),
    .B1(\line_cache[163][2] ),
    .B2(_05433_),
    .X(_06341_));
 sky130_fd_sc_hd__or2_1 _20964_ (.A(_06340_),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__a22o_1 _20965_ (.A1(_05427_),
    .A2(\line_cache[168][2] ),
    .B1(_05423_),
    .B2(\line_cache[169][2] ),
    .X(_06343_));
 sky130_fd_sc_hd__a22o_1 _20966_ (.A1(_05464_),
    .A2(\line_cache[171][2] ),
    .B1(\line_cache[170][2] ),
    .B2(_05424_),
    .X(_06344_));
 sky130_fd_sc_hd__a22o_1 _20967_ (.A1(_05463_),
    .A2(\line_cache[172][2] ),
    .B1(_05462_),
    .B2(\line_cache[173][2] ),
    .X(_06345_));
 sky130_fd_sc_hd__a221o_1 _20968_ (.A1(\line_cache[175][2] ),
    .A2(_05456_),
    .B1(\line_cache[174][2] ),
    .B2(_05461_),
    .C1(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__or3_1 _20969_ (.A(_06343_),
    .B(_06344_),
    .C(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__nor3_1 _20970_ (.A(_06339_),
    .B(_06342_),
    .C(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__a22o_1 _20971_ (.A1(_05419_),
    .A2(\line_cache[155][2] ),
    .B1(\line_cache[154][2] ),
    .B2(_06107_),
    .X(_06349_));
 sky130_fd_sc_hd__a221o_1 _20972_ (.A1(\line_cache[153][2] ),
    .A2(_05399_),
    .B1(\line_cache[152][2] ),
    .B2(_05397_),
    .C1(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__a22o_1 _20973_ (.A1(_05392_),
    .A2(\line_cache[147][2] ),
    .B1(_05386_),
    .B2(\line_cache[146][2] ),
    .X(_06351_));
 sky130_fd_sc_hd__a221oi_2 _20974_ (.A1(\line_cache[145][2] ),
    .A2(_05384_),
    .B1(\line_cache[144][2] ),
    .B2(_05380_),
    .C1(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__a22o_1 _20975_ (.A1(_05393_),
    .A2(\line_cache[148][2] ),
    .B1(\line_cache[149][2] ),
    .B2(_05391_),
    .X(_06353_));
 sky130_fd_sc_hd__a221oi_2 _20976_ (.A1(\line_cache[151][2] ),
    .A2(_05398_),
    .B1(\line_cache[150][2] ),
    .B2(_05390_),
    .C1(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__a22o_1 _20977_ (.A1(_05418_),
    .A2(\line_cache[156][2] ),
    .B1(_05417_),
    .B2(\line_cache[157][2] ),
    .X(_06355_));
 sky130_fd_sc_hd__a221oi_1 _20978_ (.A1(\line_cache[159][2] ),
    .A2(_05413_),
    .B1(\line_cache[158][2] ),
    .B2(_05416_),
    .C1(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__and4b_1 _20979_ (.A_N(_06350_),
    .B(_06352_),
    .C(_06354_),
    .D(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__a22o_1 _20980_ (.A1(_05449_),
    .A2(\line_cache[180][2] ),
    .B1(_05446_),
    .B2(\line_cache[181][2] ),
    .X(_06358_));
 sky130_fd_sc_hd__a221o_1 _20981_ (.A1(\line_cache[183][2] ),
    .A2(_05439_),
    .B1(\line_cache[182][2] ),
    .B2(_05445_),
    .C1(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__a22o_1 _20982_ (.A1(\line_cache[177][2] ),
    .A2(_05457_),
    .B1(_05453_),
    .B2(\line_cache[176][2] ),
    .X(_06360_));
 sky130_fd_sc_hd__a221o_1 _20983_ (.A1(\line_cache[179][2] ),
    .A2(_05447_),
    .B1(\line_cache[178][2] ),
    .B2(_05458_),
    .C1(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__a22o_1 _20984_ (.A1(_05438_),
    .A2(\line_cache[184][2] ),
    .B1(_05440_),
    .B2(\line_cache[185][2] ),
    .X(_06362_));
 sky130_fd_sc_hd__and2_1 _20985_ (.A(_05479_),
    .B(\line_cache[189][2] ),
    .X(_06363_));
 sky130_fd_sc_hd__a21o_1 _20986_ (.A1(\line_cache[188][2] ),
    .A2(_05480_),
    .B1(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__a22o_1 _20987_ (.A1(_05478_),
    .A2(\line_cache[190][2] ),
    .B1(_05468_),
    .B2(\line_cache[191][2] ),
    .X(_06365_));
 sky130_fd_sc_hd__a22o_1 _20988_ (.A1(_06131_),
    .A2(\line_cache[186][2] ),
    .B1(\line_cache[187][2] ),
    .B2(_05481_),
    .X(_06366_));
 sky130_fd_sc_hd__or4_1 _20989_ (.A(_06362_),
    .B(_06364_),
    .C(_06365_),
    .D(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nor3_1 _20990_ (.A(_06359_),
    .B(_06361_),
    .C(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__and3_1 _20991_ (.A(_06348_),
    .B(_06357_),
    .C(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__and3_1 _20992_ (.A(_05207_),
    .B(\line_cache[137][2] ),
    .C(_05381_),
    .X(_06370_));
 sky130_fd_sc_hd__a21o_1 _20993_ (.A1(\line_cache[136][2] ),
    .A2(_05604_),
    .B1(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__a221o_1 _20994_ (.A1(\line_cache[139][2] ),
    .A2(_05377_),
    .B1(\line_cache[138][2] ),
    .B2(_05602_),
    .C1(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__a22o_1 _20995_ (.A1(_05376_),
    .A2(\line_cache[140][2] ),
    .B1(_05375_),
    .B2(\line_cache[141][2] ),
    .X(_06373_));
 sky130_fd_sc_hd__a221o_1 _20996_ (.A1(\line_cache[143][2] ),
    .A2(_05382_),
    .B1(\line_cache[142][2] ),
    .B2(_05374_),
    .C1(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__a22o_1 _20997_ (.A1(_05612_),
    .A2(\line_cache[131][2] ),
    .B1(_05598_),
    .B2(\line_cache[130][2] ),
    .X(_06375_));
 sky130_fd_sc_hd__a221o_1 _20998_ (.A1(\line_cache[129][2] ),
    .A2(_05597_),
    .B1(\line_cache[128][2] ),
    .B2(_05594_),
    .C1(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__and2_1 _20999_ (.A(_05609_),
    .B(\line_cache[133][2] ),
    .X(_06377_));
 sky130_fd_sc_hd__and3_1 _21000_ (.A(_05611_),
    .B(\line_cache[132][2] ),
    .C(_05381_),
    .X(_06378_));
 sky130_fd_sc_hd__or2_1 _21001_ (.A(_06377_),
    .B(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__a221o_1 _21002_ (.A1(\line_cache[135][2] ),
    .A2(_05605_),
    .B1(\line_cache[134][2] ),
    .B2(_05608_),
    .C1(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__or4_1 _21003_ (.A(_06372_),
    .B(_06374_),
    .C(_06376_),
    .D(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__and3_1 _21004_ (.A(_05207_),
    .B(\line_cache[121][2] ),
    .C(_05562_),
    .X(_06382_));
 sky130_fd_sc_hd__a21o_1 _21005_ (.A1(\line_cache[120][2] ),
    .A2(_05561_),
    .B1(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__a221o_1 _21006_ (.A1(\line_cache[123][2] ),
    .A2(_05591_),
    .B1(\line_cache[122][2] ),
    .B2(_05559_),
    .C1(_06383_),
    .X(_06384_));
 sky130_fd_sc_hd__a22o_1 _21007_ (.A1(_05590_),
    .A2(\line_cache[124][2] ),
    .B1(_05589_),
    .B2(\line_cache[125][2] ),
    .X(_06385_));
 sky130_fd_sc_hd__a221o_1 _21008_ (.A1(\line_cache[127][2] ),
    .A2(_05596_),
    .B1(\line_cache[126][2] ),
    .B2(_05588_),
    .C1(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__a22o_1 _21009_ (.A1(_05568_),
    .A2(\line_cache[116][2] ),
    .B1(_05567_),
    .B2(\line_cache[117][2] ),
    .X(_06387_));
 sky130_fd_sc_hd__a221o_1 _21010_ (.A1(\line_cache[119][2] ),
    .A2(_06088_),
    .B1(\line_cache[118][2] ),
    .B2(_05566_),
    .C1(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__a22o_1 _21011_ (.A1(_05569_),
    .A2(\line_cache[115][2] ),
    .B1(_05582_),
    .B2(\line_cache[114][2] ),
    .X(_06389_));
 sky130_fd_sc_hd__a221o_1 _21012_ (.A1(\line_cache[113][2] ),
    .A2(_05581_),
    .B1(\line_cache[112][2] ),
    .B2(_05579_),
    .C1(_06389_),
    .X(_06390_));
 sky130_fd_sc_hd__or4_1 _21013_ (.A(_06384_),
    .B(_06386_),
    .C(_06388_),
    .D(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__nor2_1 _21014_ (.A(_06381_),
    .B(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__and3_2 _21015_ (.A(_06337_),
    .B(_06369_),
    .C(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__nand3_1 _21016_ (.A(_06212_),
    .B(_06314_),
    .C(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__o21a_4 _21017_ (.A1(_06144_),
    .A2(_06394_),
    .B1(_05884_),
    .X(net128));
 sky130_fd_sc_hd__nor3b_1 _21018_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][3] ),
    .Y(_06395_));
 sky130_fd_sc_hd__and3_1 _21019_ (.A(_05203_),
    .B(\line_cache[203][3] ),
    .C(_05685_),
    .X(_06396_));
 sky130_fd_sc_hd__and3_1 _21020_ (.A(_05586_),
    .B(\line_cache[206][3] ),
    .C(_05685_),
    .X(_06397_));
 sky130_fd_sc_hd__and2b_1 _21021_ (.A_N(_05687_),
    .B(\line_cache[204][3] ),
    .X(_06398_));
 sky130_fd_sc_hd__a2111o_1 _21022_ (.A1(\line_cache[205][3] ),
    .A2(_05683_),
    .B1(_06396_),
    .C1(_06397_),
    .D1(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__a22o_1 _21023_ (.A1(_05484_),
    .A2(\line_cache[195][3] ),
    .B1(_05485_),
    .B2(\line_cache[196][3] ),
    .X(_06400_));
 sky130_fd_sc_hd__a221o_1 _21024_ (.A1(\line_cache[198][3] ),
    .A2(_05487_),
    .B1(\line_cache[197][3] ),
    .B2(_05489_),
    .C1(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__a22o_1 _21025_ (.A1(_05495_),
    .A2(\line_cache[200][3] ),
    .B1(_05493_),
    .B2(\line_cache[199][3] ),
    .X(_06402_));
 sky130_fd_sc_hd__a221o_1 _21026_ (.A1(\line_cache[202][3] ),
    .A2(_05492_),
    .B1(\line_cache[201][3] ),
    .B2(_05491_),
    .C1(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__and3_1 _21027_ (.A(_05470_),
    .B(\line_cache[193][3] ),
    .C(_05472_),
    .X(_06404_));
 sky130_fd_sc_hd__and3_1 _21028_ (.A(_05475_),
    .B(\line_cache[192][3] ),
    .C(_05472_),
    .X(_06405_));
 sky130_fd_sc_hd__and3_1 _21029_ (.A(_05409_),
    .B(\line_cache[194][3] ),
    .C(_05472_),
    .X(_06406_));
 sky130_fd_sc_hd__a2111o_1 _21030_ (.A1(_05630_),
    .A2(\line_cache[286][3] ),
    .B1(_06404_),
    .C1(_06405_),
    .D1(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__or4_2 _21031_ (.A(_06399_),
    .B(_06401_),
    .C(_06403_),
    .D(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__a22o_1 _21032_ (.A1(_05676_),
    .A2(\line_cache[283][3] ),
    .B1(_05678_),
    .B2(\line_cache[282][3] ),
    .X(_06409_));
 sky130_fd_sc_hd__a22o_1 _21033_ (.A1(_05674_),
    .A2(\line_cache[284][3] ),
    .B1(_05631_),
    .B2(\line_cache[285][3] ),
    .X(_06410_));
 sky130_fd_sc_hd__a32o_1 _21034_ (.A1(_05165_),
    .A2(_05151_),
    .A3(\line_cache[278][3] ),
    .B1(_05654_),
    .B2(\line_cache[279][3] ),
    .X(_06411_));
 sky130_fd_sc_hd__a221o_1 _21035_ (.A1(\line_cache[281][3] ),
    .A2(_05677_),
    .B1(\line_cache[280][3] ),
    .B2(_05144_),
    .C1(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__a22o_1 _21036_ (.A1(_05668_),
    .A2(\line_cache[270][3] ),
    .B1(\line_cache[269][3] ),
    .B2(_05670_),
    .X(_06413_));
 sky130_fd_sc_hd__a22o_1 _21037_ (.A1(_05659_),
    .A2(\line_cache[275][3] ),
    .B1(\line_cache[274][3] ),
    .B2(_05662_),
    .X(_06414_));
 sky130_fd_sc_hd__a22o_1 _21038_ (.A1(_05658_),
    .A2(\line_cache[276][3] ),
    .B1(\line_cache[277][3] ),
    .B2(_05655_),
    .X(_06415_));
 sky130_fd_sc_hd__a22o_1 _21039_ (.A1(_05666_),
    .A2(\line_cache[272][3] ),
    .B1(\line_cache[273][3] ),
    .B2(_05660_),
    .X(_06416_));
 sky130_fd_sc_hd__or4_1 _21040_ (.A(_06413_),
    .B(_06414_),
    .C(_06415_),
    .D(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__or4_1 _21041_ (.A(_06409_),
    .B(_06410_),
    .C(_06412_),
    .D(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__nor2_1 _21042_ (.A(_06408_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__and3_1 _21043_ (.A(_05058_),
    .B(_05059_),
    .C(\line_cache[302][3] ),
    .X(_06420_));
 sky130_fd_sc_hd__a22o_1 _21044_ (.A1(_05056_),
    .A2(\line_cache[301][3] ),
    .B1(\line_cache[300][3] ),
    .B2(_05053_),
    .X(_06421_));
 sky130_fd_sc_hd__a211o_1 _21045_ (.A1(\line_cache[256][3] ),
    .A2(_05777_),
    .B1(_06420_),
    .C1(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__and3_1 _21046_ (.A(_05779_),
    .B(_05176_),
    .C(\line_cache[258][3] ),
    .X(_06423_));
 sky130_fd_sc_hd__and3_1 _21047_ (.A(_05771_),
    .B(_05059_),
    .C(\line_cache[260][3] ),
    .X(_06424_));
 sky130_fd_sc_hd__and3_1 _21048_ (.A(_05778_),
    .B(_05059_),
    .C(\line_cache[259][3] ),
    .X(_06425_));
 sky130_fd_sc_hd__a2111o_1 _21049_ (.A1(\line_cache[257][3] ),
    .A2(_05776_),
    .B1(_06423_),
    .C1(_06424_),
    .D1(_06425_),
    .X(_06426_));
 sky130_fd_sc_hd__and3_1 _21050_ (.A(_05356_),
    .B(_05059_),
    .C(\line_cache[267][3] ),
    .X(_06427_));
 sky130_fd_sc_hd__a22o_1 _21051_ (.A1(_05760_),
    .A2(\line_cache[266][3] ),
    .B1(\line_cache[265][3] ),
    .B2(_05764_),
    .X(_06428_));
 sky130_fd_sc_hd__a311o_1 _21052_ (.A1(_05113_),
    .A2(\line_cache[268][3] ),
    .A3(_05364_),
    .B1(_06427_),
    .C1(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__nand2_1 _21053_ (.A(_05768_),
    .B(\line_cache[262][3] ),
    .Y(_06430_));
 sky130_fd_sc_hd__nand2_1 _21054_ (.A(_05773_),
    .B(\line_cache[261][3] ),
    .Y(_06431_));
 sky130_fd_sc_hd__nand2_1 _21055_ (.A(_06430_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__a221oi_2 _21056_ (.A1(_05763_),
    .A2(\line_cache[264][3] ),
    .B1(_05770_),
    .B2(\line_cache[263][3] ),
    .C1(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__or4b_1 _21057_ (.A(_06422_),
    .B(_06426_),
    .C(_06429_),
    .D_N(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__a22o_1 _21058_ (.A1(_05098_),
    .A2(\line_cache[308][3] ),
    .B1(\line_cache[309][3] ),
    .B2(_05093_),
    .X(_06435_));
 sky130_fd_sc_hd__a221o_1 _21059_ (.A1(\line_cache[311][3] ),
    .A2(_05097_),
    .B1(\line_cache[310][3] ),
    .B2(_05103_),
    .C1(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__a22o_1 _21060_ (.A1(_05046_),
    .A2(\line_cache[295][3] ),
    .B1(\line_cache[294][3] ),
    .B2(_05043_),
    .X(_06437_));
 sky130_fd_sc_hd__a221o_1 _21061_ (.A1(\line_cache[293][3] ),
    .A2(_05628_),
    .B1(\line_cache[292][3] ),
    .B2(_05627_),
    .C1(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__a22o_1 _21062_ (.A1(_05069_),
    .A2(\line_cache[296][3] ),
    .B1(\line_cache[297][3] ),
    .B2(_05076_),
    .X(_06439_));
 sky130_fd_sc_hd__a221o_1 _21063_ (.A1(\line_cache[299][3] ),
    .A2(_05073_),
    .B1(\line_cache[298][3] ),
    .B2(_05079_),
    .C1(_06439_),
    .X(_06440_));
 sky130_fd_sc_hd__a22o_1 _21064_ (.A1(_05632_),
    .A2(\line_cache[288][3] ),
    .B1(\line_cache[289][3] ),
    .B2(_05633_),
    .X(_06441_));
 sky130_fd_sc_hd__a221o_1 _21065_ (.A1(\line_cache[291][3] ),
    .A2(_05623_),
    .B1(\line_cache[290][3] ),
    .B2(_05624_),
    .C1(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__or4_1 _21066_ (.A(_06436_),
    .B(_06438_),
    .C(_06440_),
    .D(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__nor2_1 _21067_ (.A(_06434_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__nand2_1 _21068_ (.A(_06419_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__and3_1 _21069_ (.A(_05454_),
    .B(\line_cache[239][3] ),
    .C(_05194_),
    .X(_06446_));
 sky130_fd_sc_hd__and3_1 _21070_ (.A(_05470_),
    .B(\line_cache[241][3] ),
    .C(_05206_),
    .X(_06447_));
 sky130_fd_sc_hd__and3_1 _21071_ (.A(_05409_),
    .B(\line_cache[242][3] ),
    .C(_05206_),
    .X(_06448_));
 sky130_fd_sc_hd__a2111o_1 _21072_ (.A1(_05233_),
    .A2(\line_cache[240][3] ),
    .B1(_06446_),
    .C1(_06447_),
    .D1(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__and2_1 _21073_ (.A(_05235_),
    .B(\line_cache[243][3] ),
    .X(_06450_));
 sky130_fd_sc_hd__a21o_1 _21074_ (.A1(\line_cache[244][3] ),
    .A2(_05224_),
    .B1(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__a221o_1 _21075_ (.A1(\line_cache[246][3] ),
    .A2(_05753_),
    .B1(\line_cache[245][3] ),
    .B2(_05226_),
    .C1(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__a22o_1 _21076_ (.A1(_05212_),
    .A2(\line_cache[252][3] ),
    .B1(_05205_),
    .B2(\line_cache[251][3] ),
    .X(_06453_));
 sky130_fd_sc_hd__a221o_1 _21077_ (.A1(\line_cache[254][3] ),
    .A2(_05217_),
    .B1(\line_cache[253][3] ),
    .B2(_05214_),
    .C1(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__a22o_1 _21078_ (.A1(_05750_),
    .A2(\line_cache[248][3] ),
    .B1(_05229_),
    .B2(\line_cache[247][3] ),
    .X(_06455_));
 sky130_fd_sc_hd__a221o_1 _21079_ (.A1(\line_cache[250][3] ),
    .A2(_05202_),
    .B1(\line_cache[249][3] ),
    .B2(_05209_),
    .C1(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__or4_1 _21080_ (.A(_06449_),
    .B(_06452_),
    .C(_06454_),
    .D(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__a22o_1 _21081_ (.A1(_05873_),
    .A2(\line_cache[68][3] ),
    .B1(_05872_),
    .B2(\line_cache[69][3] ),
    .X(_06458_));
 sky130_fd_sc_hd__a221o_1 _21082_ (.A1(\line_cache[71][3] ),
    .A2(_05868_),
    .B1(\line_cache[70][3] ),
    .B2(_05871_),
    .C1(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__and2_1 _21083_ (.A(_05860_),
    .B(\line_cache[65][3] ),
    .X(_06460_));
 sky130_fd_sc_hd__a21o_1 _21084_ (.A1(_05858_),
    .A2(\line_cache[64][3] ),
    .B1(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__a221o_1 _21085_ (.A1(\line_cache[67][3] ),
    .A2(_05875_),
    .B1(\line_cache[66][3] ),
    .B2(_05861_),
    .C1(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__and3_1 _21086_ (.A(_05200_),
    .B(\line_cache[74][3] ),
    .C(_05536_),
    .X(_06463_));
 sky130_fd_sc_hd__a22o_1 _21087_ (.A1(_05867_),
    .A2(\line_cache[72][3] ),
    .B1(_05866_),
    .B2(\line_cache[73][3] ),
    .X(_06464_));
 sky130_fd_sc_hd__a32o_1 _21088_ (.A1(_05544_),
    .A2(\line_cache[77][3] ),
    .A3(_05536_),
    .B1(\line_cache[76][3] ),
    .B2(_05542_),
    .X(_06465_));
 sky130_fd_sc_hd__a221o_1 _21089_ (.A1(\line_cache[79][3] ),
    .A2(_05537_),
    .B1(\line_cache[78][3] ),
    .B2(_05545_),
    .C1(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__a2111oi_1 _21090_ (.A1(\line_cache[75][3] ),
    .A2(_05543_),
    .B1(_06463_),
    .C1(_06464_),
    .D1(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__or3b_2 _21091_ (.A(_06459_),
    .B(_06462_),
    .C_N(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__nor2_1 _21092_ (.A(_06457_),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__a22o_1 _21093_ (.A1(_05746_),
    .A2(\line_cache[236][3] ),
    .B1(_05747_),
    .B2(\line_cache[235][3] ),
    .X(_06470_));
 sky130_fd_sc_hd__a221o_1 _21094_ (.A1(\line_cache[238][3] ),
    .A2(_05744_),
    .B1(\line_cache[237][3] ),
    .B2(_05745_),
    .C1(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__and3_1 _21095_ (.A(_05470_),
    .B(\line_cache[225][3] ),
    .C(_05194_),
    .X(_06472_));
 sky130_fd_sc_hd__and3_1 _21096_ (.A(_05408_),
    .B(\line_cache[226][3] ),
    .C(_05194_),
    .X(_06473_));
 sky130_fd_sc_hd__and3_1 _21097_ (.A(_05475_),
    .B(\line_cache[224][3] ),
    .C(_05194_),
    .X(_06474_));
 sky130_fd_sc_hd__a2111o_1 _21098_ (.A1(\line_cache[223][3] ),
    .A2(_05720_),
    .B1(_06472_),
    .C1(_06473_),
    .D1(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__and3_1 _21099_ (.A(_05704_),
    .B(\line_cache[227][3] ),
    .C(_05732_),
    .X(_06476_));
 sky130_fd_sc_hd__and3_1 _21100_ (.A(_05611_),
    .B(\line_cache[228][3] ),
    .C(_05721_),
    .X(_06477_));
 sky130_fd_sc_hd__and3_1 _21101_ (.A(_05710_),
    .B(\line_cache[229][3] ),
    .C(_05721_),
    .X(_06478_));
 sky130_fd_sc_hd__and3_1 _21102_ (.A(_05708_),
    .B(\line_cache[230][3] ),
    .C(_05194_),
    .X(_06479_));
 sky130_fd_sc_hd__or4_1 _21103_ (.A(_06476_),
    .B(_06477_),
    .C(_06478_),
    .D(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__a22o_1 _21104_ (.A1(_05728_),
    .A2(\line_cache[232][3] ),
    .B1(_05729_),
    .B2(\line_cache[231][3] ),
    .X(_06481_));
 sky130_fd_sc_hd__a221o_1 _21105_ (.A1(\line_cache[234][3] ),
    .A2(_05726_),
    .B1(\line_cache[233][3] ),
    .B2(_05727_),
    .C1(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__or4_1 _21106_ (.A(_06471_),
    .B(_06475_),
    .C(_06480_),
    .D(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__a22o_1 _21107_ (.A1(_05716_),
    .A2(\line_cache[220][3] ),
    .B1(_05717_),
    .B2(\line_cache[219][3] ),
    .X(_06484_));
 sky130_fd_sc_hd__a221o_1 _21108_ (.A1(\line_cache[222][3] ),
    .A2(_05714_),
    .B1(\line_cache[221][3] ),
    .B2(_05715_),
    .C1(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__a22o_1 _21109_ (.A1(_05700_),
    .A2(\line_cache[209][3] ),
    .B1(\line_cache[210][3] ),
    .B2(_05701_),
    .X(_06486_));
 sky130_fd_sc_hd__a221o_1 _21110_ (.A1(\line_cache[208][3] ),
    .A2(_05698_),
    .B1(\line_cache[207][3] ),
    .B2(_05699_),
    .C1(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__and3_1 _21111_ (.A(_05704_),
    .B(\line_cache[211][3] ),
    .C(_05706_),
    .X(_06488_));
 sky130_fd_sc_hd__and3_1 _21112_ (.A(_05611_),
    .B(\line_cache[212][3] ),
    .C(_05706_),
    .X(_06489_));
 sky130_fd_sc_hd__and3_1 _21113_ (.A(_05710_),
    .B(\line_cache[213][3] ),
    .C(_05706_),
    .X(_06490_));
 sky130_fd_sc_hd__and3_1 _21114_ (.A(_05708_),
    .B(\line_cache[214][3] ),
    .C(_05706_),
    .X(_06491_));
 sky130_fd_sc_hd__or4_2 _21115_ (.A(_06488_),
    .B(_06489_),
    .C(_06490_),
    .D(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__a22o_1 _21116_ (.A1(_05692_),
    .A2(\line_cache[216][3] ),
    .B1(_05983_),
    .B2(\line_cache[215][3] ),
    .X(_06493_));
 sky130_fd_sc_hd__a221o_1 _21117_ (.A1(\line_cache[218][3] ),
    .A2(_05690_),
    .B1(\line_cache[217][3] ),
    .B2(_05691_),
    .C1(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__or4_2 _21118_ (.A(_06485_),
    .B(_06487_),
    .C(_06492_),
    .D(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__nor2_1 _21119_ (.A(_06483_),
    .B(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__nand2_1 _21120_ (.A(_06469_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__nor2_1 _21121_ (.A(_06445_),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__and2_1 _21122_ (.A(_05797_),
    .B(\line_cache[1][3] ),
    .X(_06499_));
 sky130_fd_sc_hd__and3_1 _21123_ (.A(_05779_),
    .B(_05991_),
    .C(\line_cache[2][3] ),
    .X(_06500_));
 sky130_fd_sc_hd__a211o_1 _21124_ (.A1(\line_cache[15][3] ),
    .A2(_05798_),
    .B1(_06499_),
    .C1(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__and3_1 _21125_ (.A(_05778_),
    .B(_05792_),
    .C(\line_cache[3][3] ),
    .X(_06502_));
 sky130_fd_sc_hd__a31o_1 _21126_ (.A1(_05840_),
    .A2(\line_cache[4][3] ),
    .A3(_05771_),
    .B1(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__a221o_1 _21127_ (.A1(_05343_),
    .A2(\line_cache[5][3] ),
    .B1(\line_cache[6][3] ),
    .B2(_05348_),
    .C1(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__and3_1 _21128_ (.A(_05112_),
    .B(_05151_),
    .C(\line_cache[319][3] ),
    .X(_06505_));
 sky130_fd_sc_hd__a32o_1 _21129_ (.A1(_05991_),
    .A2(_05180_),
    .A3(\line_cache[31][3] ),
    .B1(_05998_),
    .B2(\line_cache[47][3] ),
    .X(_06506_));
 sky130_fd_sc_hd__a311o_1 _21130_ (.A1(_05188_),
    .A2(\line_cache[63][3] ),
    .A3(_05112_),
    .B1(_06505_),
    .C1(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__nand2_1 _21131_ (.A(_05787_),
    .B(\line_cache[303][3] ),
    .Y(_06508_));
 sky130_fd_sc_hd__nand2_1 _21132_ (.A(_05791_),
    .B(\line_cache[271][3] ),
    .Y(_06509_));
 sky130_fd_sc_hd__nand2_1 _21133_ (.A(_06508_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__a221oi_4 _21134_ (.A1(\line_cache[255][3] ),
    .A2(_05220_),
    .B1(\line_cache[287][3] ),
    .B2(_05788_),
    .C1(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__or4b_1 _21135_ (.A(_06501_),
    .B(_06504_),
    .C(_06507_),
    .D_N(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__a22o_1 _21136_ (.A1(_05283_),
    .A2(\line_cache[45][3] ),
    .B1(\line_cache[46][3] ),
    .B2(_05285_),
    .X(_06513_));
 sky130_fd_sc_hd__a22o_1 _21137_ (.A1(_05298_),
    .A2(\line_cache[48][3] ),
    .B1(\line_cache[49][3] ),
    .B2(_05300_),
    .X(_06514_));
 sky130_fd_sc_hd__nand2_1 _21138_ (.A(_05279_),
    .B(\line_cache[41][3] ),
    .Y(_06515_));
 sky130_fd_sc_hd__nand2_1 _21139_ (.A(_05281_),
    .B(\line_cache[42][3] ),
    .Y(_06516_));
 sky130_fd_sc_hd__nand2_1 _21140_ (.A(_06515_),
    .B(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__a221oi_1 _21141_ (.A1(_05277_),
    .A2(\line_cache[43][3] ),
    .B1(\line_cache[44][3] ),
    .B2(_05287_),
    .C1(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__or3b_2 _21142_ (.A(_06513_),
    .B(_06514_),
    .C_N(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__a22o_1 _21143_ (.A1(_05106_),
    .A2(\line_cache[317][3] ),
    .B1(\line_cache[316][3] ),
    .B2(_05108_),
    .X(_06520_));
 sky130_fd_sc_hd__a22o_1 _21144_ (.A1(_05292_),
    .A2(\line_cache[61][3] ),
    .B1(\line_cache[60][3] ),
    .B2(_05294_),
    .X(_06521_));
 sky130_fd_sc_hd__a22o_1 _21145_ (.A1(_05312_),
    .A2(\line_cache[58][3] ),
    .B1(_05317_),
    .B2(\line_cache[59][3] ),
    .X(_06522_));
 sky130_fd_sc_hd__and3_1 _21146_ (.A(_05109_),
    .B(_05021_),
    .C(\line_cache[318][3] ),
    .X(_06523_));
 sky130_fd_sc_hd__a21o_1 _21147_ (.A1(\line_cache[62][3] ),
    .A2(_05296_),
    .B1(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__or4_1 _21148_ (.A(_06520_),
    .B(_06521_),
    .C(_06522_),
    .D(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__a22o_1 _21149_ (.A1(_05129_),
    .A2(\line_cache[304][3] ),
    .B1(\line_cache[305][3] ),
    .B2(_05127_),
    .X(_06526_));
 sky130_fd_sc_hd__a22o_1 _21150_ (.A1(_05119_),
    .A2(\line_cache[312][3] ),
    .B1(\line_cache[313][3] ),
    .B2(_05121_),
    .X(_06527_));
 sky130_fd_sc_hd__a22o_1 _21151_ (.A1(_05123_),
    .A2(\line_cache[314][3] ),
    .B1(_05644_),
    .B2(\line_cache[315][3] ),
    .X(_06528_));
 sky130_fd_sc_hd__a22o_1 _21152_ (.A1(_05132_),
    .A2(\line_cache[306][3] ),
    .B1(\line_cache[307][3] ),
    .B2(_05136_),
    .X(_06529_));
 sky130_fd_sc_hd__or4_1 _21153_ (.A(_06526_),
    .B(_06527_),
    .C(_06528_),
    .D(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__a22o_1 _21154_ (.A1(_05314_),
    .A2(\line_cache[56][3] ),
    .B1(\line_cache[57][3] ),
    .B2(_05315_),
    .X(_06531_));
 sky130_fd_sc_hd__a22o_1 _21155_ (.A1(_05304_),
    .A2(\line_cache[52][3] ),
    .B1(\line_cache[53][3] ),
    .B2(_05306_),
    .X(_06532_));
 sky130_fd_sc_hd__a22o_1 _21156_ (.A1(_05301_),
    .A2(\line_cache[50][3] ),
    .B1(\line_cache[51][3] ),
    .B2(_05302_),
    .X(_06533_));
 sky130_fd_sc_hd__a22o_1 _21157_ (.A1(_05307_),
    .A2(\line_cache[54][3] ),
    .B1(_05309_),
    .B2(\line_cache[55][3] ),
    .X(_06534_));
 sky130_fd_sc_hd__or4_2 _21158_ (.A(_06531_),
    .B(_06532_),
    .C(_06533_),
    .D(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__or4_1 _21159_ (.A(_06519_),
    .B(_06525_),
    .C(_06530_),
    .D(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__or2b_1 _21160_ (.A(_05365_),
    .B_N(\line_cache[12][3] ),
    .X(_06537_));
 sky130_fd_sc_hd__nand2_1 _21161_ (.A(_05358_),
    .B(\line_cache[11][3] ),
    .Y(_06538_));
 sky130_fd_sc_hd__nand2_1 _21162_ (.A(_06537_),
    .B(_06538_),
    .Y(_06539_));
 sky130_fd_sc_hd__a221oi_1 _21163_ (.A1(\line_cache[14][3] ),
    .A2(_05838_),
    .B1(\line_cache[13][3] ),
    .B2(_05839_),
    .C1(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand2_1 _21164_ (.A(_05353_),
    .B(\line_cache[10][3] ),
    .Y(_06541_));
 sky130_fd_sc_hd__nand2_1 _21165_ (.A(_05351_),
    .B(\line_cache[9][3] ),
    .Y(_06542_));
 sky130_fd_sc_hd__nand2_1 _21166_ (.A(_06541_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__a221oi_2 _21167_ (.A1(_05355_),
    .A2(\line_cache[8][3] ),
    .B1(_05346_),
    .B2(\line_cache[7][3] ),
    .C1(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__nand2_1 _21168_ (.A(_06540_),
    .B(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__and3_1 _21169_ (.A(_05163_),
    .B(_05187_),
    .C(\line_cache[21][3] ),
    .X(_06546_));
 sky130_fd_sc_hd__and3_1 _21170_ (.A(_05167_),
    .B(_05187_),
    .C(\line_cache[20][3] ),
    .X(_06547_));
 sky130_fd_sc_hd__a22o_1 _21171_ (.A1(_05825_),
    .A2(\line_cache[23][3] ),
    .B1(\line_cache[22][3] ),
    .B2(_05826_),
    .X(_06548_));
 sky130_fd_sc_hd__a22o_1 _21172_ (.A1(_05329_),
    .A2(\line_cache[16][3] ),
    .B1(\line_cache[17][3] ),
    .B2(_05330_),
    .X(_06549_));
 sky130_fd_sc_hd__a221o_1 _21173_ (.A1(\line_cache[19][3] ),
    .A2(_05831_),
    .B1(\line_cache[18][3] ),
    .B2(_05832_),
    .C1(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__or4_2 _21174_ (.A(_06546_),
    .B(_06547_),
    .C(_06548_),
    .D(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__a22o_1 _21175_ (.A1(_05262_),
    .A2(\line_cache[33][3] ),
    .B1(\line_cache[34][3] ),
    .B2(_05263_),
    .X(_06552_));
 sky130_fd_sc_hd__a221o_1 _21176_ (.A1(\line_cache[36][3] ),
    .A2(_05266_),
    .B1(\line_cache[35][3] ),
    .B2(_05261_),
    .C1(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__and3_1 _21177_ (.A(_05146_),
    .B(_05792_),
    .C(\line_cache[25][3] ),
    .X(_06554_));
 sky130_fd_sc_hd__a31o_1 _21178_ (.A1(_05991_),
    .A2(\line_cache[24][3] ),
    .A3(_05320_),
    .B1(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__a221oi_4 _21179_ (.A1(\line_cache[27][3] ),
    .A2(_05817_),
    .B1(\line_cache[26][3] ),
    .B2(_05819_),
    .C1(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__a32o_1 _21180_ (.A1(_05175_),
    .A2(_05812_),
    .A3(\line_cache[30][3] ),
    .B1(_05260_),
    .B2(\line_cache[32][3] ),
    .X(_06557_));
 sky130_fd_sc_hd__a32o_1 _21181_ (.A1(_05991_),
    .A2(_05173_),
    .A3(\line_cache[29][3] ),
    .B1(_06051_),
    .B2(\line_cache[28][3] ),
    .X(_06558_));
 sky130_fd_sc_hd__nor2_1 _21182_ (.A(_06557_),
    .B(_06558_),
    .Y(_06559_));
 sky130_fd_sc_hd__nand2_1 _21183_ (.A(_05270_),
    .B(\line_cache[38][3] ),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_1 _21184_ (.A(_05272_),
    .B(\line_cache[37][3] ),
    .Y(_06561_));
 sky130_fd_sc_hd__nand2_1 _21185_ (.A(_06560_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__a221oi_1 _21186_ (.A1(_05268_),
    .A2(\line_cache[39][3] ),
    .B1(\line_cache[40][3] ),
    .B2(_05275_),
    .C1(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__and4b_1 _21187_ (.A_N(_06553_),
    .B(_06556_),
    .C(_06559_),
    .D(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__or3b_2 _21188_ (.A(_06545_),
    .B(_06551_),
    .C_N(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__nor3_2 _21189_ (.A(_06512_),
    .B(_06536_),
    .C(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__a22o_1 _21190_ (.A1(_05510_),
    .A2(\line_cache[99][3] ),
    .B1(_05516_),
    .B2(\line_cache[98][3] ),
    .X(_06567_));
 sky130_fd_sc_hd__a221o_1 _21191_ (.A1(\line_cache[97][3] ),
    .A2(_05515_),
    .B1(\line_cache[96][3] ),
    .B2(_05520_),
    .C1(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__a22o_1 _21192_ (.A1(_05575_),
    .A2(\line_cache[108][3] ),
    .B1(_05574_),
    .B2(\line_cache[109][3] ),
    .X(_06569_));
 sky130_fd_sc_hd__a221o_1 _21193_ (.A1(\line_cache[111][3] ),
    .A2(_05580_),
    .B1(\line_cache[110][3] ),
    .B2(_05573_),
    .C1(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__a22o_1 _21194_ (.A1(_05511_),
    .A2(\line_cache[100][3] ),
    .B1(\line_cache[101][3] ),
    .B2(_05509_),
    .X(_06571_));
 sky130_fd_sc_hd__a221o_1 _21195_ (.A1(\line_cache[103][3] ),
    .A2(_05504_),
    .B1(\line_cache[102][3] ),
    .B2(_05502_),
    .C1(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__and2_1 _21196_ (.A(_05503_),
    .B(\line_cache[104][3] ),
    .X(_06573_));
 sky130_fd_sc_hd__a21o_1 _21197_ (.A1(\line_cache[105][3] ),
    .A2(_05508_),
    .B1(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__a221o_1 _21198_ (.A1(\line_cache[107][3] ),
    .A2(_05576_),
    .B1(\line_cache[106][3] ),
    .B2(_05506_),
    .C1(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__or4_1 _21199_ (.A(_06568_),
    .B(_06570_),
    .C(_06572_),
    .D(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__a22o_1 _21200_ (.A1(_05531_),
    .A2(\line_cache[83][3] ),
    .B1(_05539_),
    .B2(\line_cache[82][3] ),
    .X(_06577_));
 sky130_fd_sc_hd__a221o_1 _21201_ (.A1(\line_cache[81][3] ),
    .A2(_05538_),
    .B1(\line_cache[80][3] ),
    .B2(_05535_),
    .C1(_06577_),
    .X(_06578_));
 sky130_fd_sc_hd__a22o_1 _21202_ (.A1(_05524_),
    .A2(\line_cache[92][3] ),
    .B1(_05523_),
    .B2(\line_cache[93][3] ),
    .X(_06579_));
 sky130_fd_sc_hd__a221o_1 _21203_ (.A1(\line_cache[95][3] ),
    .A2(_05519_),
    .B1(\line_cache[94][3] ),
    .B2(_05522_),
    .C1(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__a22o_1 _21204_ (.A1(_05532_),
    .A2(\line_cache[84][3] ),
    .B1(\line_cache[85][3] ),
    .B2(_05530_),
    .X(_06581_));
 sky130_fd_sc_hd__a221o_1 _21205_ (.A1(\line_cache[87][3] ),
    .A2(_05551_),
    .B1(\line_cache[86][3] ),
    .B2(_05529_),
    .C1(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__a22o_1 _21206_ (.A1(_05553_),
    .A2(\line_cache[88][3] ),
    .B1(_05549_),
    .B2(\line_cache[89][3] ),
    .X(_06583_));
 sky130_fd_sc_hd__a221o_1 _21207_ (.A1(\line_cache[91][3] ),
    .A2(_05525_),
    .B1(\line_cache[90][3] ),
    .B2(_05550_),
    .C1(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__or4_1 _21208_ (.A(_06578_),
    .B(_06580_),
    .C(_06582_),
    .D(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__nor2_1 _21209_ (.A(_06576_),
    .B(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__a22o_1 _21210_ (.A1(\line_cache[177][3] ),
    .A2(_05457_),
    .B1(_05453_),
    .B2(\line_cache[176][3] ),
    .X(_06587_));
 sky130_fd_sc_hd__a221o_1 _21211_ (.A1(\line_cache[179][3] ),
    .A2(_05447_),
    .B1(\line_cache[178][3] ),
    .B2(_05458_),
    .C1(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__a22o_1 _21212_ (.A1(_05478_),
    .A2(\line_cache[190][3] ),
    .B1(_05468_),
    .B2(\line_cache[191][3] ),
    .X(_06589_));
 sky130_fd_sc_hd__a221oi_2 _21213_ (.A1(\line_cache[189][3] ),
    .A2(_05479_),
    .B1(\line_cache[188][3] ),
    .B2(_05480_),
    .C1(_06589_),
    .Y(_06590_));
 sky130_fd_sc_hd__a22o_1 _21214_ (.A1(_05438_),
    .A2(\line_cache[184][3] ),
    .B1(_05440_),
    .B2(\line_cache[185][3] ),
    .X(_06591_));
 sky130_fd_sc_hd__a221oi_1 _21215_ (.A1(\line_cache[187][3] ),
    .A2(_05481_),
    .B1(\line_cache[186][3] ),
    .B2(_06131_),
    .C1(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__a22o_1 _21216_ (.A1(_05449_),
    .A2(\line_cache[180][3] ),
    .B1(_05446_),
    .B2(\line_cache[181][3] ),
    .X(_06593_));
 sky130_fd_sc_hd__a221oi_2 _21217_ (.A1(\line_cache[183][3] ),
    .A2(_05439_),
    .B1(\line_cache[182][3] ),
    .B2(_05445_),
    .C1(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__and4b_1 _21218_ (.A_N(_06588_),
    .B(_06590_),
    .C(_06592_),
    .D(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__a22o_1 _21219_ (.A1(_05397_),
    .A2(\line_cache[152][3] ),
    .B1(_05399_),
    .B2(\line_cache[153][3] ),
    .X(_06596_));
 sky130_fd_sc_hd__a221o_1 _21220_ (.A1(\line_cache[155][3] ),
    .A2(_05419_),
    .B1(\line_cache[154][3] ),
    .B2(_06107_),
    .C1(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__a22o_1 _21221_ (.A1(_05392_),
    .A2(\line_cache[147][3] ),
    .B1(_05386_),
    .B2(\line_cache[146][3] ),
    .X(_06598_));
 sky130_fd_sc_hd__a221oi_4 _21222_ (.A1(\line_cache[145][3] ),
    .A2(_05384_),
    .B1(\line_cache[144][3] ),
    .B2(_05380_),
    .C1(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__a22o_1 _21223_ (.A1(_05393_),
    .A2(\line_cache[148][3] ),
    .B1(\line_cache[149][3] ),
    .B2(_05391_),
    .X(_06600_));
 sky130_fd_sc_hd__a221oi_2 _21224_ (.A1(\line_cache[151][3] ),
    .A2(_05398_),
    .B1(\line_cache[150][3] ),
    .B2(_05390_),
    .C1(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__a22o_1 _21225_ (.A1(_05418_),
    .A2(\line_cache[156][3] ),
    .B1(_05417_),
    .B2(\line_cache[157][3] ),
    .X(_06602_));
 sky130_fd_sc_hd__a221oi_1 _21226_ (.A1(\line_cache[159][3] ),
    .A2(_05413_),
    .B1(\line_cache[158][3] ),
    .B2(_05416_),
    .C1(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__and4b_1 _21227_ (.A_N(_06597_),
    .B(_06599_),
    .C(_06601_),
    .D(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__a22o_1 _21228_ (.A1(_05464_),
    .A2(\line_cache[171][3] ),
    .B1(\line_cache[170][3] ),
    .B2(_05424_),
    .X(_06605_));
 sky130_fd_sc_hd__a221o_1 _21229_ (.A1(\line_cache[169][3] ),
    .A2(_05423_),
    .B1(\line_cache[168][3] ),
    .B2(_05427_),
    .C1(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__a32o_1 _21230_ (.A1(_05409_),
    .A2(\line_cache[162][3] ),
    .A3(_05410_),
    .B1(\line_cache[163][3] ),
    .B2(_05433_),
    .X(_06607_));
 sky130_fd_sc_hd__a221oi_1 _21231_ (.A1(\line_cache[161][3] ),
    .A2(_05406_),
    .B1(\line_cache[160][3] ),
    .B2(_05414_),
    .C1(_06607_),
    .Y(_06608_));
 sky130_fd_sc_hd__a22o_1 _21232_ (.A1(_05434_),
    .A2(\line_cache[164][3] ),
    .B1(\line_cache[165][3] ),
    .B2(_05432_),
    .X(_06609_));
 sky130_fd_sc_hd__nand2_1 _21233_ (.A(_05431_),
    .B(\line_cache[166][3] ),
    .Y(_06610_));
 sky130_fd_sc_hd__nand2_1 _21234_ (.A(_05425_),
    .B(\line_cache[167][3] ),
    .Y(_06611_));
 sky130_fd_sc_hd__and3b_1 _21235_ (.A_N(_06609_),
    .B(_06610_),
    .C(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__nand2_1 _21236_ (.A(_05462_),
    .B(\line_cache[173][3] ),
    .Y(_06613_));
 sky130_fd_sc_hd__nand2_1 _21237_ (.A(_05463_),
    .B(\line_cache[172][3] ),
    .Y(_06614_));
 sky130_fd_sc_hd__nand2_1 _21238_ (.A(_06613_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__a221oi_1 _21239_ (.A1(_05461_),
    .A2(\line_cache[174][3] ),
    .B1(_05456_),
    .B2(\line_cache[175][3] ),
    .C1(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__and4b_1 _21240_ (.A_N(_06606_),
    .B(_06608_),
    .C(_06612_),
    .D(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__and3_1 _21241_ (.A(_06595_),
    .B(_06604_),
    .C(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__and3_1 _21242_ (.A(_05586_),
    .B(\line_cache[126][3] ),
    .C(_05562_),
    .X(_06619_));
 sky130_fd_sc_hd__a21o_1 _21243_ (.A1(\line_cache[127][3] ),
    .A2(_05596_),
    .B1(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__a221o_1 _21244_ (.A1(\line_cache[125][3] ),
    .A2(_05589_),
    .B1(\line_cache[124][3] ),
    .B2(_05590_),
    .C1(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__a22o_1 _21245_ (.A1(_05569_),
    .A2(\line_cache[115][3] ),
    .B1(_05582_),
    .B2(\line_cache[114][3] ),
    .X(_06622_));
 sky130_fd_sc_hd__a221o_1 _21246_ (.A1(\line_cache[113][3] ),
    .A2(_05581_),
    .B1(\line_cache[112][3] ),
    .B2(_05579_),
    .C1(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__a22o_1 _21247_ (.A1(_05568_),
    .A2(\line_cache[116][3] ),
    .B1(_05567_),
    .B2(\line_cache[117][3] ),
    .X(_06624_));
 sky130_fd_sc_hd__a221o_1 _21248_ (.A1(\line_cache[119][3] ),
    .A2(_06088_),
    .B1(\line_cache[118][3] ),
    .B2(_05566_),
    .C1(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__a22o_1 _21249_ (.A1(_05561_),
    .A2(\line_cache[120][3] ),
    .B1(_05560_),
    .B2(\line_cache[121][3] ),
    .X(_06626_));
 sky130_fd_sc_hd__a221o_1 _21250_ (.A1(\line_cache[123][3] ),
    .A2(_05591_),
    .B1(\line_cache[122][3] ),
    .B2(_05559_),
    .C1(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__or4_1 _21251_ (.A(_06621_),
    .B(_06623_),
    .C(_06625_),
    .D(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__a22o_1 _21252_ (.A1(_05376_),
    .A2(\line_cache[140][3] ),
    .B1(_05375_),
    .B2(\line_cache[141][3] ),
    .X(_06629_));
 sky130_fd_sc_hd__a221o_1 _21253_ (.A1(\line_cache[143][3] ),
    .A2(_05382_),
    .B1(\line_cache[142][3] ),
    .B2(_05374_),
    .C1(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__a22o_1 _21254_ (.A1(_05612_),
    .A2(\line_cache[131][3] ),
    .B1(_05598_),
    .B2(\line_cache[130][3] ),
    .X(_06631_));
 sky130_fd_sc_hd__a221o_1 _21255_ (.A1(\line_cache[129][3] ),
    .A2(_05597_),
    .B1(\line_cache[128][3] ),
    .B2(_05594_),
    .C1(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__and2_1 _21256_ (.A(_05609_),
    .B(\line_cache[133][3] ),
    .X(_06633_));
 sky130_fd_sc_hd__and3_1 _21257_ (.A(_05611_),
    .B(\line_cache[132][3] ),
    .C(_05381_),
    .X(_06634_));
 sky130_fd_sc_hd__or2_1 _21258_ (.A(_06633_),
    .B(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__a221o_1 _21259_ (.A1(\line_cache[135][3] ),
    .A2(_05605_),
    .B1(\line_cache[134][3] ),
    .B2(_05608_),
    .C1(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__a22o_1 _21260_ (.A1(_05604_),
    .A2(\line_cache[136][3] ),
    .B1(_05603_),
    .B2(\line_cache[137][3] ),
    .X(_06637_));
 sky130_fd_sc_hd__a221o_1 _21261_ (.A1(\line_cache[139][3] ),
    .A2(_05377_),
    .B1(\line_cache[138][3] ),
    .B2(_05602_),
    .C1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__or4_1 _21262_ (.A(_06630_),
    .B(_06632_),
    .C(_06636_),
    .D(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__nor2_1 _21263_ (.A(_06628_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__and3_1 _21264_ (.A(_06586_),
    .B(_06618_),
    .C(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__nand3_1 _21265_ (.A(_06498_),
    .B(_06566_),
    .C(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__o21a_2 _21266_ (.A1(_06395_),
    .A2(_06642_),
    .B1(_05884_),
    .X(net129));
 sky130_fd_sc_hd__nor3b_1 _21267_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][4] ),
    .Y(_06643_));
 sky130_fd_sc_hd__and2_1 _21268_ (.A(_05797_),
    .B(\line_cache[1][4] ),
    .X(_06644_));
 sky130_fd_sc_hd__and3_1 _21269_ (.A(_05779_),
    .B(_05840_),
    .C(\line_cache[2][4] ),
    .X(_06645_));
 sky130_fd_sc_hd__a211o_1 _21270_ (.A1(\line_cache[15][4] ),
    .A2(_05798_),
    .B1(_06644_),
    .C1(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__and3_1 _21271_ (.A(_05778_),
    .B(_05792_),
    .C(\line_cache[3][4] ),
    .X(_06647_));
 sky130_fd_sc_hd__a31o_1 _21272_ (.A1(_05188_),
    .A2(\line_cache[4][4] ),
    .A3(_05771_),
    .B1(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__a221o_1 _21273_ (.A1(_05343_),
    .A2(\line_cache[5][4] ),
    .B1(\line_cache[6][4] ),
    .B2(_05348_),
    .C1(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__and3_1 _21274_ (.A(_05112_),
    .B(_05151_),
    .C(\line_cache[319][4] ),
    .X(_06650_));
 sky130_fd_sc_hd__a32o_1 _21275_ (.A1(_05991_),
    .A2(_05180_),
    .A3(\line_cache[31][4] ),
    .B1(_05998_),
    .B2(\line_cache[47][4] ),
    .X(_06651_));
 sky130_fd_sc_hd__a311o_1 _21276_ (.A1(_05188_),
    .A2(\line_cache[63][4] ),
    .A3(_05112_),
    .B1(_06650_),
    .C1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__nand2_1 _21277_ (.A(_05787_),
    .B(\line_cache[303][4] ),
    .Y(_06653_));
 sky130_fd_sc_hd__nand2_1 _21278_ (.A(_05791_),
    .B(\line_cache[271][4] ),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_1 _21279_ (.A(_06653_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__a221oi_4 _21280_ (.A1(\line_cache[255][4] ),
    .A2(_05220_),
    .B1(\line_cache[287][4] ),
    .B2(_05788_),
    .C1(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__or4b_1 _21281_ (.A(_06646_),
    .B(_06649_),
    .C(_06652_),
    .D_N(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__a22o_1 _21282_ (.A1(_05283_),
    .A2(\line_cache[45][4] ),
    .B1(\line_cache[46][4] ),
    .B2(_05285_),
    .X(_06658_));
 sky130_fd_sc_hd__a22o_1 _21283_ (.A1(_05298_),
    .A2(\line_cache[48][4] ),
    .B1(\line_cache[49][4] ),
    .B2(_05300_),
    .X(_06659_));
 sky130_fd_sc_hd__nand2_1 _21284_ (.A(_05279_),
    .B(\line_cache[41][4] ),
    .Y(_06660_));
 sky130_fd_sc_hd__nand2_1 _21285_ (.A(_05281_),
    .B(\line_cache[42][4] ),
    .Y(_06661_));
 sky130_fd_sc_hd__nand2_1 _21286_ (.A(_06660_),
    .B(_06661_),
    .Y(_06662_));
 sky130_fd_sc_hd__a221oi_1 _21287_ (.A1(_05277_),
    .A2(\line_cache[43][4] ),
    .B1(\line_cache[44][4] ),
    .B2(_05287_),
    .C1(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__or3b_2 _21288_ (.A(_06658_),
    .B(_06659_),
    .C_N(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__a22o_1 _21289_ (.A1(_05106_),
    .A2(\line_cache[317][4] ),
    .B1(\line_cache[316][4] ),
    .B2(_05108_),
    .X(_06665_));
 sky130_fd_sc_hd__a22o_1 _21290_ (.A1(_05292_),
    .A2(\line_cache[61][4] ),
    .B1(\line_cache[60][4] ),
    .B2(_05294_),
    .X(_06666_));
 sky130_fd_sc_hd__a22o_1 _21291_ (.A1(_05312_),
    .A2(\line_cache[58][4] ),
    .B1(_05317_),
    .B2(\line_cache[59][4] ),
    .X(_06667_));
 sky130_fd_sc_hd__and3_1 _21292_ (.A(_05109_),
    .B(_05021_),
    .C(\line_cache[318][4] ),
    .X(_06668_));
 sky130_fd_sc_hd__a21o_1 _21293_ (.A1(\line_cache[62][4] ),
    .A2(_05296_),
    .B1(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__or4_1 _21294_ (.A(_06665_),
    .B(_06666_),
    .C(_06667_),
    .D(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__a22o_1 _21295_ (.A1(_05129_),
    .A2(\line_cache[304][4] ),
    .B1(\line_cache[305][4] ),
    .B2(_05127_),
    .X(_06671_));
 sky130_fd_sc_hd__a22o_1 _21296_ (.A1(_05119_),
    .A2(\line_cache[312][4] ),
    .B1(\line_cache[313][4] ),
    .B2(_05121_),
    .X(_06672_));
 sky130_fd_sc_hd__a22o_1 _21297_ (.A1(_05123_),
    .A2(\line_cache[314][4] ),
    .B1(_05644_),
    .B2(\line_cache[315][4] ),
    .X(_06673_));
 sky130_fd_sc_hd__a22o_1 _21298_ (.A1(_05132_),
    .A2(\line_cache[306][4] ),
    .B1(\line_cache[307][4] ),
    .B2(_05136_),
    .X(_06674_));
 sky130_fd_sc_hd__or4_1 _21299_ (.A(_06671_),
    .B(_06672_),
    .C(_06673_),
    .D(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__a22o_1 _21300_ (.A1(_05314_),
    .A2(\line_cache[56][4] ),
    .B1(\line_cache[57][4] ),
    .B2(_05315_),
    .X(_06676_));
 sky130_fd_sc_hd__a22o_1 _21301_ (.A1(_05304_),
    .A2(\line_cache[52][4] ),
    .B1(\line_cache[53][4] ),
    .B2(_05306_),
    .X(_06677_));
 sky130_fd_sc_hd__a22o_1 _21302_ (.A1(_05301_),
    .A2(\line_cache[50][4] ),
    .B1(\line_cache[51][4] ),
    .B2(_05302_),
    .X(_06678_));
 sky130_fd_sc_hd__a22o_1 _21303_ (.A1(_05307_),
    .A2(\line_cache[54][4] ),
    .B1(_05309_),
    .B2(\line_cache[55][4] ),
    .X(_06679_));
 sky130_fd_sc_hd__or4_2 _21304_ (.A(_06676_),
    .B(_06677_),
    .C(_06678_),
    .D(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__or4_1 _21305_ (.A(_06664_),
    .B(_06670_),
    .C(_06675_),
    .D(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__or2b_1 _21306_ (.A(_05365_),
    .B_N(\line_cache[12][4] ),
    .X(_06682_));
 sky130_fd_sc_hd__nand2_1 _21307_ (.A(_05358_),
    .B(\line_cache[11][4] ),
    .Y(_06683_));
 sky130_fd_sc_hd__nand2_1 _21308_ (.A(_06682_),
    .B(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__a221oi_1 _21309_ (.A1(\line_cache[14][4] ),
    .A2(_05838_),
    .B1(\line_cache[13][4] ),
    .B2(_05839_),
    .C1(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__nand2_1 _21310_ (.A(_05353_),
    .B(\line_cache[10][4] ),
    .Y(_06686_));
 sky130_fd_sc_hd__nand2_1 _21311_ (.A(_05351_),
    .B(\line_cache[9][4] ),
    .Y(_06687_));
 sky130_fd_sc_hd__nand2_1 _21312_ (.A(_06686_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__a221oi_2 _21313_ (.A1(_05355_),
    .A2(\line_cache[8][4] ),
    .B1(_05346_),
    .B2(\line_cache[7][4] ),
    .C1(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__nand2_1 _21314_ (.A(_06685_),
    .B(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__and3_1 _21315_ (.A(_05163_),
    .B(_05812_),
    .C(\line_cache[21][4] ),
    .X(_06691_));
 sky130_fd_sc_hd__and3_1 _21316_ (.A(_05167_),
    .B(_05812_),
    .C(\line_cache[20][4] ),
    .X(_06692_));
 sky130_fd_sc_hd__a22o_1 _21317_ (.A1(_05825_),
    .A2(\line_cache[23][4] ),
    .B1(\line_cache[22][4] ),
    .B2(_05826_),
    .X(_06693_));
 sky130_fd_sc_hd__a22o_1 _21318_ (.A1(_05329_),
    .A2(\line_cache[16][4] ),
    .B1(\line_cache[17][4] ),
    .B2(_05330_),
    .X(_06694_));
 sky130_fd_sc_hd__a221o_1 _21319_ (.A1(\line_cache[19][4] ),
    .A2(_05831_),
    .B1(\line_cache[18][4] ),
    .B2(_05832_),
    .C1(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__or4_1 _21320_ (.A(_06691_),
    .B(_06692_),
    .C(_06693_),
    .D(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__a22o_1 _21321_ (.A1(_05262_),
    .A2(\line_cache[33][4] ),
    .B1(\line_cache[34][4] ),
    .B2(_05263_),
    .X(_06697_));
 sky130_fd_sc_hd__a221o_1 _21322_ (.A1(\line_cache[36][4] ),
    .A2(_05266_),
    .B1(\line_cache[35][4] ),
    .B2(_05261_),
    .C1(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__and3_1 _21323_ (.A(_05146_),
    .B(_05792_),
    .C(\line_cache[25][4] ),
    .X(_06699_));
 sky130_fd_sc_hd__a31o_1 _21324_ (.A1(_05840_),
    .A2(\line_cache[24][4] ),
    .A3(_05320_),
    .B1(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__a221oi_2 _21325_ (.A1(\line_cache[27][4] ),
    .A2(_05817_),
    .B1(\line_cache[26][4] ),
    .B2(_05819_),
    .C1(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__a32o_1 _21326_ (.A1(_05175_),
    .A2(_05812_),
    .A3(\line_cache[30][4] ),
    .B1(_05260_),
    .B2(\line_cache[32][4] ),
    .X(_06702_));
 sky130_fd_sc_hd__a32o_1 _21327_ (.A1(_05840_),
    .A2(_05173_),
    .A3(\line_cache[29][4] ),
    .B1(_06051_),
    .B2(\line_cache[28][4] ),
    .X(_06703_));
 sky130_fd_sc_hd__nor2_1 _21328_ (.A(_06702_),
    .B(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__nand2_1 _21329_ (.A(_05270_),
    .B(\line_cache[38][4] ),
    .Y(_06705_));
 sky130_fd_sc_hd__nand2_1 _21330_ (.A(_05272_),
    .B(\line_cache[37][4] ),
    .Y(_06706_));
 sky130_fd_sc_hd__nand2_1 _21331_ (.A(_06705_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__a221oi_1 _21332_ (.A1(_05268_),
    .A2(\line_cache[39][4] ),
    .B1(\line_cache[40][4] ),
    .B2(_05275_),
    .C1(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__and4b_1 _21333_ (.A_N(_06698_),
    .B(_06701_),
    .C(_06704_),
    .D(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__or3b_2 _21334_ (.A(_06690_),
    .B(_06696_),
    .C_N(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__nor3_2 _21335_ (.A(_06657_),
    .B(_06681_),
    .C(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__and3_1 _21336_ (.A(_05203_),
    .B(\line_cache[203][4] ),
    .C(_05685_),
    .X(_06712_));
 sky130_fd_sc_hd__and3_1 _21337_ (.A(_05586_),
    .B(\line_cache[206][4] ),
    .C(_05685_),
    .X(_06713_));
 sky130_fd_sc_hd__and2b_1 _21338_ (.A_N(_05687_),
    .B(\line_cache[204][4] ),
    .X(_06714_));
 sky130_fd_sc_hd__a2111o_1 _21339_ (.A1(\line_cache[205][4] ),
    .A2(_05683_),
    .B1(_06712_),
    .C1(_06713_),
    .D1(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__a22o_1 _21340_ (.A1(_05484_),
    .A2(\line_cache[195][4] ),
    .B1(_05485_),
    .B2(\line_cache[196][4] ),
    .X(_06716_));
 sky130_fd_sc_hd__a221o_1 _21341_ (.A1(\line_cache[198][4] ),
    .A2(_05487_),
    .B1(\line_cache[197][4] ),
    .B2(_05489_),
    .C1(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__a22o_1 _21342_ (.A1(_05495_),
    .A2(\line_cache[200][4] ),
    .B1(_05493_),
    .B2(\line_cache[199][4] ),
    .X(_06718_));
 sky130_fd_sc_hd__a221o_1 _21343_ (.A1(\line_cache[202][4] ),
    .A2(_05492_),
    .B1(\line_cache[201][4] ),
    .B2(_05491_),
    .C1(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__and3_1 _21344_ (.A(_05470_),
    .B(\line_cache[193][4] ),
    .C(_05685_),
    .X(_06720_));
 sky130_fd_sc_hd__and3_1 _21345_ (.A(_05475_),
    .B(\line_cache[192][4] ),
    .C(_05472_),
    .X(_06721_));
 sky130_fd_sc_hd__and3_1 _21346_ (.A(_05409_),
    .B(\line_cache[194][4] ),
    .C(_05472_),
    .X(_06722_));
 sky130_fd_sc_hd__a2111o_1 _21347_ (.A1(_05630_),
    .A2(\line_cache[286][4] ),
    .B1(_06720_),
    .C1(_06721_),
    .D1(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__or4_1 _21348_ (.A(_06715_),
    .B(_06717_),
    .C(_06719_),
    .D(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__a22o_1 _21349_ (.A1(_05676_),
    .A2(\line_cache[283][4] ),
    .B1(_05678_),
    .B2(\line_cache[282][4] ),
    .X(_06725_));
 sky130_fd_sc_hd__a22o_1 _21350_ (.A1(_05674_),
    .A2(\line_cache[284][4] ),
    .B1(_05631_),
    .B2(\line_cache[285][4] ),
    .X(_06726_));
 sky130_fd_sc_hd__a32o_1 _21351_ (.A1(_05165_),
    .A2(_05059_),
    .A3(\line_cache[278][4] ),
    .B1(_05654_),
    .B2(\line_cache[279][4] ),
    .X(_06727_));
 sky130_fd_sc_hd__a221o_1 _21352_ (.A1(\line_cache[281][4] ),
    .A2(_05677_),
    .B1(\line_cache[280][4] ),
    .B2(_05144_),
    .C1(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__a22o_1 _21353_ (.A1(_05668_),
    .A2(\line_cache[270][4] ),
    .B1(\line_cache[269][4] ),
    .B2(_05670_),
    .X(_06729_));
 sky130_fd_sc_hd__a22o_1 _21354_ (.A1(_05659_),
    .A2(\line_cache[275][4] ),
    .B1(\line_cache[274][4] ),
    .B2(_05662_),
    .X(_06730_));
 sky130_fd_sc_hd__a22o_1 _21355_ (.A1(_05658_),
    .A2(\line_cache[276][4] ),
    .B1(\line_cache[277][4] ),
    .B2(_05655_),
    .X(_06731_));
 sky130_fd_sc_hd__a22o_1 _21356_ (.A1(_05666_),
    .A2(\line_cache[272][4] ),
    .B1(\line_cache[273][4] ),
    .B2(_05660_),
    .X(_06732_));
 sky130_fd_sc_hd__or4_1 _21357_ (.A(_06729_),
    .B(_06730_),
    .C(_06731_),
    .D(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__or4_2 _21358_ (.A(_06725_),
    .B(_06726_),
    .C(_06728_),
    .D(_06733_),
    .X(_06734_));
 sky130_fd_sc_hd__nor2_1 _21359_ (.A(_06724_),
    .B(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__a22o_1 _21360_ (.A1(_05746_),
    .A2(\line_cache[236][4] ),
    .B1(_05747_),
    .B2(\line_cache[235][4] ),
    .X(_06736_));
 sky130_fd_sc_hd__a221o_1 _21361_ (.A1(\line_cache[238][4] ),
    .A2(_05744_),
    .B1(\line_cache[237][4] ),
    .B2(_05745_),
    .C1(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__and3_1 _21362_ (.A(_05469_),
    .B(\line_cache[225][4] ),
    .C(_05732_),
    .X(_06738_));
 sky130_fd_sc_hd__and3_1 _21363_ (.A(_05408_),
    .B(\line_cache[226][4] ),
    .C(_05721_),
    .X(_06739_));
 sky130_fd_sc_hd__and3_1 _21364_ (.A(_05475_),
    .B(\line_cache[224][4] ),
    .C(_05194_),
    .X(_06740_));
 sky130_fd_sc_hd__a2111o_1 _21365_ (.A1(\line_cache[223][4] ),
    .A2(_05720_),
    .B1(_06738_),
    .C1(_06739_),
    .D1(_06740_),
    .X(_06741_));
 sky130_fd_sc_hd__and3_1 _21366_ (.A(_05704_),
    .B(\line_cache[227][4] ),
    .C(_05193_),
    .X(_06742_));
 sky130_fd_sc_hd__and3_1 _21367_ (.A(_05610_),
    .B(\line_cache[228][4] ),
    .C(_05193_),
    .X(_06743_));
 sky130_fd_sc_hd__and3_1 _21368_ (.A(_05710_),
    .B(\line_cache[229][4] ),
    .C(_05193_),
    .X(_06744_));
 sky130_fd_sc_hd__and3_1 _21369_ (.A(_05708_),
    .B(\line_cache[230][4] ),
    .C(_05732_),
    .X(_06745_));
 sky130_fd_sc_hd__or4_1 _21370_ (.A(_06742_),
    .B(_06743_),
    .C(_06744_),
    .D(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__a22o_1 _21371_ (.A1(_05728_),
    .A2(\line_cache[232][4] ),
    .B1(_05729_),
    .B2(\line_cache[231][4] ),
    .X(_06747_));
 sky130_fd_sc_hd__a221o_1 _21372_ (.A1(\line_cache[234][4] ),
    .A2(_05726_),
    .B1(\line_cache[233][4] ),
    .B2(_05727_),
    .C1(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__or4_1 _21373_ (.A(_06737_),
    .B(_06741_),
    .C(_06746_),
    .D(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__a22o_1 _21374_ (.A1(_05716_),
    .A2(\line_cache[220][4] ),
    .B1(_05717_),
    .B2(\line_cache[219][4] ),
    .X(_06750_));
 sky130_fd_sc_hd__a221o_1 _21375_ (.A1(\line_cache[222][4] ),
    .A2(_05714_),
    .B1(\line_cache[221][4] ),
    .B2(_05715_),
    .C1(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__a22o_1 _21376_ (.A1(_05700_),
    .A2(\line_cache[209][4] ),
    .B1(\line_cache[210][4] ),
    .B2(_05701_),
    .X(_06752_));
 sky130_fd_sc_hd__a221o_1 _21377_ (.A1(\line_cache[208][4] ),
    .A2(_05698_),
    .B1(\line_cache[207][4] ),
    .B2(_05699_),
    .C1(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__and3_1 _21378_ (.A(_05704_),
    .B(\line_cache[211][4] ),
    .C(_05694_),
    .X(_06754_));
 sky130_fd_sc_hd__and3_1 _21379_ (.A(_05611_),
    .B(\line_cache[212][4] ),
    .C(_05694_),
    .X(_06755_));
 sky130_fd_sc_hd__and3_1 _21380_ (.A(_05710_),
    .B(\line_cache[213][4] ),
    .C(_05694_),
    .X(_06756_));
 sky130_fd_sc_hd__and3_1 _21381_ (.A(_05708_),
    .B(\line_cache[214][4] ),
    .C(_05706_),
    .X(_06757_));
 sky130_fd_sc_hd__or4_1 _21382_ (.A(_06754_),
    .B(_06755_),
    .C(_06756_),
    .D(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__a22o_1 _21383_ (.A1(_05692_),
    .A2(\line_cache[216][4] ),
    .B1(_05983_),
    .B2(\line_cache[215][4] ),
    .X(_06759_));
 sky130_fd_sc_hd__a221o_1 _21384_ (.A1(\line_cache[218][4] ),
    .A2(_05690_),
    .B1(\line_cache[217][4] ),
    .B2(_05691_),
    .C1(_06759_),
    .X(_06760_));
 sky130_fd_sc_hd__or4_2 _21385_ (.A(_06751_),
    .B(_06753_),
    .C(_06758_),
    .D(_06760_),
    .X(_06761_));
 sky130_fd_sc_hd__and3_1 _21386_ (.A(_05454_),
    .B(\line_cache[239][4] ),
    .C(_05192_),
    .X(_06762_));
 sky130_fd_sc_hd__and3_1 _21387_ (.A(_05469_),
    .B(\line_cache[241][4] ),
    .C(_05198_),
    .X(_06763_));
 sky130_fd_sc_hd__and3_1 _21388_ (.A(_05408_),
    .B(\line_cache[242][4] ),
    .C(_05198_),
    .X(_06764_));
 sky130_fd_sc_hd__a2111o_1 _21389_ (.A1(_05233_),
    .A2(\line_cache[240][4] ),
    .B1(_06762_),
    .C1(_06763_),
    .D1(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__and2_1 _21390_ (.A(_05235_),
    .B(\line_cache[243][4] ),
    .X(_06766_));
 sky130_fd_sc_hd__a21o_1 _21391_ (.A1(\line_cache[244][4] ),
    .A2(_05224_),
    .B1(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__a221o_1 _21392_ (.A1(\line_cache[246][4] ),
    .A2(_05753_),
    .B1(\line_cache[245][4] ),
    .B2(_05226_),
    .C1(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__a22o_1 _21393_ (.A1(_05212_),
    .A2(\line_cache[252][4] ),
    .B1(_05205_),
    .B2(\line_cache[251][4] ),
    .X(_06769_));
 sky130_fd_sc_hd__a221o_1 _21394_ (.A1(\line_cache[254][4] ),
    .A2(_05217_),
    .B1(\line_cache[253][4] ),
    .B2(_05214_),
    .C1(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__a22o_1 _21395_ (.A1(_05750_),
    .A2(\line_cache[248][4] ),
    .B1(_05229_),
    .B2(\line_cache[247][4] ),
    .X(_06771_));
 sky130_fd_sc_hd__a221o_1 _21396_ (.A1(\line_cache[250][4] ),
    .A2(_05202_),
    .B1(\line_cache[249][4] ),
    .B2(_05209_),
    .C1(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__or4_1 _21397_ (.A(_06765_),
    .B(_06768_),
    .C(_06770_),
    .D(_06772_),
    .X(_06773_));
 sky130_fd_sc_hd__a22o_1 _21398_ (.A1(_05545_),
    .A2(\line_cache[78][4] ),
    .B1(_05537_),
    .B2(\line_cache[79][4] ),
    .X(_06774_));
 sky130_fd_sc_hd__a32o_1 _21399_ (.A1(_05544_),
    .A2(\line_cache[77][4] ),
    .A3(_05536_),
    .B1(\line_cache[76][4] ),
    .B2(_05542_),
    .X(_06775_));
 sky130_fd_sc_hd__or2_1 _21400_ (.A(_06774_),
    .B(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__and2_1 _21401_ (.A(_05860_),
    .B(\line_cache[65][4] ),
    .X(_06777_));
 sky130_fd_sc_hd__a21o_1 _21402_ (.A1(_05858_),
    .A2(\line_cache[64][4] ),
    .B1(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__a221o_1 _21403_ (.A1(\line_cache[67][4] ),
    .A2(_05875_),
    .B1(\line_cache[66][4] ),
    .B2(_05861_),
    .C1(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__a22o_1 _21404_ (.A1(_05867_),
    .A2(\line_cache[72][4] ),
    .B1(_05866_),
    .B2(\line_cache[73][4] ),
    .X(_06780_));
 sky130_fd_sc_hd__a221o_1 _21405_ (.A1(\line_cache[75][4] ),
    .A2(_05543_),
    .B1(\line_cache[74][4] ),
    .B2(_05865_),
    .C1(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__a22o_1 _21406_ (.A1(_05873_),
    .A2(\line_cache[68][4] ),
    .B1(_05872_),
    .B2(\line_cache[69][4] ),
    .X(_06782_));
 sky130_fd_sc_hd__a221o_1 _21407_ (.A1(\line_cache[71][4] ),
    .A2(_05868_),
    .B1(\line_cache[70][4] ),
    .B2(_05871_),
    .C1(_06782_),
    .X(_06783_));
 sky130_fd_sc_hd__or4_4 _21408_ (.A(_06776_),
    .B(_06779_),
    .C(_06781_),
    .D(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__or2_1 _21409_ (.A(_06773_),
    .B(_06784_),
    .X(_06785_));
 sky130_fd_sc_hd__nor3_1 _21410_ (.A(_06749_),
    .B(_06761_),
    .C(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__and3_1 _21411_ (.A(_05058_),
    .B(_05034_),
    .C(\line_cache[302][4] ),
    .X(_06787_));
 sky130_fd_sc_hd__a22o_1 _21412_ (.A1(_05056_),
    .A2(\line_cache[301][4] ),
    .B1(\line_cache[300][4] ),
    .B2(_05053_),
    .X(_06788_));
 sky130_fd_sc_hd__a211o_1 _21413_ (.A1(\line_cache[256][4] ),
    .A2(_05777_),
    .B1(_06787_),
    .C1(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__and3_1 _21414_ (.A(_05779_),
    .B(_05021_),
    .C(\line_cache[258][4] ),
    .X(_06790_));
 sky130_fd_sc_hd__and3_1 _21415_ (.A(_05771_),
    .B(_05034_),
    .C(\line_cache[260][4] ),
    .X(_06791_));
 sky130_fd_sc_hd__and3_1 _21416_ (.A(_05778_),
    .B(_05034_),
    .C(\line_cache[259][4] ),
    .X(_06792_));
 sky130_fd_sc_hd__a2111o_1 _21417_ (.A1(\line_cache[257][4] ),
    .A2(_05776_),
    .B1(_06790_),
    .C1(_06791_),
    .D1(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__and3_1 _21418_ (.A(_05356_),
    .B(_05176_),
    .C(\line_cache[267][4] ),
    .X(_06794_));
 sky130_fd_sc_hd__a22o_1 _21419_ (.A1(_05760_),
    .A2(\line_cache[266][4] ),
    .B1(\line_cache[265][4] ),
    .B2(_05764_),
    .X(_06795_));
 sky130_fd_sc_hd__a311o_1 _21420_ (.A1(_05113_),
    .A2(\line_cache[268][4] ),
    .A3(_05364_),
    .B1(_06794_),
    .C1(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__nand2_1 _21421_ (.A(_05768_),
    .B(\line_cache[262][4] ),
    .Y(_06797_));
 sky130_fd_sc_hd__nand2_1 _21422_ (.A(_05773_),
    .B(\line_cache[261][4] ),
    .Y(_06798_));
 sky130_fd_sc_hd__nand2_1 _21423_ (.A(_06797_),
    .B(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__a221oi_2 _21424_ (.A1(_05763_),
    .A2(\line_cache[264][4] ),
    .B1(_05770_),
    .B2(\line_cache[263][4] ),
    .C1(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__or4b_1 _21425_ (.A(_06789_),
    .B(_06793_),
    .C(_06796_),
    .D_N(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__a22o_1 _21426_ (.A1(_05098_),
    .A2(\line_cache[308][4] ),
    .B1(\line_cache[309][4] ),
    .B2(_05093_),
    .X(_06802_));
 sky130_fd_sc_hd__a221o_1 _21427_ (.A1(\line_cache[311][4] ),
    .A2(_05097_),
    .B1(\line_cache[310][4] ),
    .B2(_05103_),
    .C1(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__a22o_1 _21428_ (.A1(_05046_),
    .A2(\line_cache[295][4] ),
    .B1(\line_cache[294][4] ),
    .B2(_05043_),
    .X(_06804_));
 sky130_fd_sc_hd__a221o_1 _21429_ (.A1(\line_cache[293][4] ),
    .A2(_05628_),
    .B1(\line_cache[292][4] ),
    .B2(_05627_),
    .C1(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__a22o_1 _21430_ (.A1(_05069_),
    .A2(\line_cache[296][4] ),
    .B1(\line_cache[297][4] ),
    .B2(_05076_),
    .X(_06806_));
 sky130_fd_sc_hd__a221o_1 _21431_ (.A1(\line_cache[299][4] ),
    .A2(_05073_),
    .B1(\line_cache[298][4] ),
    .B2(_05079_),
    .C1(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__a22o_1 _21432_ (.A1(_05632_),
    .A2(\line_cache[288][4] ),
    .B1(\line_cache[289][4] ),
    .B2(_05633_),
    .X(_06808_));
 sky130_fd_sc_hd__a221o_1 _21433_ (.A1(\line_cache[291][4] ),
    .A2(_05623_),
    .B1(\line_cache[290][4] ),
    .B2(_05624_),
    .C1(_06808_),
    .X(_06809_));
 sky130_fd_sc_hd__or4_1 _21434_ (.A(_06803_),
    .B(_06805_),
    .C(_06807_),
    .D(_06809_),
    .X(_06810_));
 sky130_fd_sc_hd__nor2_1 _21435_ (.A(_06801_),
    .B(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__and3_2 _21436_ (.A(_06735_),
    .B(_06786_),
    .C(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__a22o_1 _21437_ (.A1(_05425_),
    .A2(\line_cache[167][4] ),
    .B1(\line_cache[166][4] ),
    .B2(_05431_),
    .X(_06813_));
 sky130_fd_sc_hd__a221o_1 _21438_ (.A1(\line_cache[165][4] ),
    .A2(_05432_),
    .B1(\line_cache[164][4] ),
    .B2(_05434_),
    .C1(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__and3_1 _21439_ (.A(_05207_),
    .B(\line_cache[169][4] ),
    .C(_05410_),
    .X(_06815_));
 sky130_fd_sc_hd__a22o_1 _21440_ (.A1(_05464_),
    .A2(\line_cache[171][4] ),
    .B1(\line_cache[170][4] ),
    .B2(_05424_),
    .X(_06816_));
 sky130_fd_sc_hd__a22o_1 _21441_ (.A1(_05463_),
    .A2(\line_cache[172][4] ),
    .B1(_05462_),
    .B2(\line_cache[173][4] ),
    .X(_06817_));
 sky130_fd_sc_hd__a221o_1 _21442_ (.A1(\line_cache[175][4] ),
    .A2(_05456_),
    .B1(\line_cache[174][4] ),
    .B2(_05461_),
    .C1(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__a2111oi_1 _21443_ (.A1(\line_cache[168][4] ),
    .A2(_05427_),
    .B1(_06815_),
    .C1(_06816_),
    .D1(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__a32o_1 _21444_ (.A1(_05409_),
    .A2(\line_cache[162][4] ),
    .A3(_05410_),
    .B1(\line_cache[163][4] ),
    .B2(_05433_),
    .X(_06820_));
 sky130_fd_sc_hd__a221oi_1 _21445_ (.A1(\line_cache[161][4] ),
    .A2(_05406_),
    .B1(\line_cache[160][4] ),
    .B2(_05414_),
    .C1(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__and3b_1 _21446_ (.A_N(_06814_),
    .B(_06819_),
    .C(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__a22o_1 _21447_ (.A1(\line_cache[177][4] ),
    .A2(_05457_),
    .B1(_05453_),
    .B2(\line_cache[176][4] ),
    .X(_06823_));
 sky130_fd_sc_hd__a221o_1 _21448_ (.A1(\line_cache[179][4] ),
    .A2(_05447_),
    .B1(\line_cache[178][4] ),
    .B2(_05458_),
    .C1(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__a22o_1 _21449_ (.A1(_05478_),
    .A2(\line_cache[190][4] ),
    .B1(_05468_),
    .B2(\line_cache[191][4] ),
    .X(_06825_));
 sky130_fd_sc_hd__a221oi_2 _21450_ (.A1(\line_cache[189][4] ),
    .A2(_05479_),
    .B1(\line_cache[188][4] ),
    .B2(_05480_),
    .C1(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__a22o_1 _21451_ (.A1(_05438_),
    .A2(\line_cache[184][4] ),
    .B1(_05440_),
    .B2(\line_cache[185][4] ),
    .X(_06827_));
 sky130_fd_sc_hd__a221oi_1 _21452_ (.A1(\line_cache[187][4] ),
    .A2(_05481_),
    .B1(\line_cache[186][4] ),
    .B2(_06131_),
    .C1(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__a22o_1 _21453_ (.A1(_05449_),
    .A2(\line_cache[180][4] ),
    .B1(_05446_),
    .B2(\line_cache[181][4] ),
    .X(_06829_));
 sky130_fd_sc_hd__a221oi_2 _21454_ (.A1(\line_cache[183][4] ),
    .A2(_05439_),
    .B1(\line_cache[182][4] ),
    .B2(_05445_),
    .C1(_06829_),
    .Y(_06830_));
 sky130_fd_sc_hd__and4b_1 _21455_ (.A_N(_06824_),
    .B(_06826_),
    .C(_06828_),
    .D(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__a22o_1 _21456_ (.A1(_05419_),
    .A2(\line_cache[155][4] ),
    .B1(\line_cache[154][4] ),
    .B2(_06107_),
    .X(_06832_));
 sky130_fd_sc_hd__a221o_1 _21457_ (.A1(\line_cache[153][4] ),
    .A2(_05399_),
    .B1(\line_cache[152][4] ),
    .B2(_05397_),
    .C1(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__a22o_1 _21458_ (.A1(_05392_),
    .A2(\line_cache[147][4] ),
    .B1(_05386_),
    .B2(\line_cache[146][4] ),
    .X(_06834_));
 sky130_fd_sc_hd__a221oi_2 _21459_ (.A1(\line_cache[145][4] ),
    .A2(_05384_),
    .B1(\line_cache[144][4] ),
    .B2(_05380_),
    .C1(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__a22o_1 _21460_ (.A1(_05393_),
    .A2(\line_cache[148][4] ),
    .B1(\line_cache[149][4] ),
    .B2(_05391_),
    .X(_06836_));
 sky130_fd_sc_hd__a221oi_1 _21461_ (.A1(\line_cache[151][4] ),
    .A2(_05398_),
    .B1(\line_cache[150][4] ),
    .B2(_05390_),
    .C1(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__a22o_1 _21462_ (.A1(_05418_),
    .A2(\line_cache[156][4] ),
    .B1(_05417_),
    .B2(\line_cache[157][4] ),
    .X(_06838_));
 sky130_fd_sc_hd__a221oi_1 _21463_ (.A1(\line_cache[159][4] ),
    .A2(_05413_),
    .B1(\line_cache[158][4] ),
    .B2(_05416_),
    .C1(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__and4b_1 _21464_ (.A_N(_06833_),
    .B(_06835_),
    .C(_06837_),
    .D(_06839_),
    .X(_06840_));
 sky130_fd_sc_hd__and3_1 _21465_ (.A(_06822_),
    .B(_06831_),
    .C(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__a22o_1 _21466_ (.A1(_05510_),
    .A2(\line_cache[99][4] ),
    .B1(_05516_),
    .B2(\line_cache[98][4] ),
    .X(_06842_));
 sky130_fd_sc_hd__a221o_1 _21467_ (.A1(\line_cache[97][4] ),
    .A2(_05515_),
    .B1(\line_cache[96][4] ),
    .B2(_05520_),
    .C1(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__a22o_1 _21468_ (.A1(_05575_),
    .A2(\line_cache[108][4] ),
    .B1(_05574_),
    .B2(\line_cache[109][4] ),
    .X(_06844_));
 sky130_fd_sc_hd__a221o_1 _21469_ (.A1(\line_cache[111][4] ),
    .A2(_05580_),
    .B1(\line_cache[110][4] ),
    .B2(_05573_),
    .C1(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__and2_1 _21470_ (.A(_05502_),
    .B(\line_cache[102][4] ),
    .X(_06846_));
 sky130_fd_sc_hd__a21o_1 _21471_ (.A1(\line_cache[103][4] ),
    .A2(_05504_),
    .B1(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__a221o_1 _21472_ (.A1(\line_cache[101][4] ),
    .A2(_05509_),
    .B1(\line_cache[100][4] ),
    .B2(_05511_),
    .C1(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__and2_1 _21473_ (.A(_05503_),
    .B(\line_cache[104][4] ),
    .X(_06849_));
 sky130_fd_sc_hd__a21o_1 _21474_ (.A1(\line_cache[105][4] ),
    .A2(_05508_),
    .B1(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__a221o_1 _21475_ (.A1(\line_cache[107][4] ),
    .A2(_05576_),
    .B1(\line_cache[106][4] ),
    .B2(_05506_),
    .C1(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__or4_1 _21476_ (.A(_06843_),
    .B(_06845_),
    .C(_06848_),
    .D(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__a22o_1 _21477_ (.A1(_05531_),
    .A2(\line_cache[83][4] ),
    .B1(_05539_),
    .B2(\line_cache[82][4] ),
    .X(_06853_));
 sky130_fd_sc_hd__a221o_1 _21478_ (.A1(\line_cache[81][4] ),
    .A2(_05538_),
    .B1(\line_cache[80][4] ),
    .B2(_05535_),
    .C1(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__a22o_1 _21479_ (.A1(_05524_),
    .A2(\line_cache[92][4] ),
    .B1(_05523_),
    .B2(\line_cache[93][4] ),
    .X(_06855_));
 sky130_fd_sc_hd__a221o_1 _21480_ (.A1(\line_cache[95][4] ),
    .A2(_05519_),
    .B1(\line_cache[94][4] ),
    .B2(_05522_),
    .C1(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__a22o_1 _21481_ (.A1(_05532_),
    .A2(\line_cache[84][4] ),
    .B1(\line_cache[85][4] ),
    .B2(_05530_),
    .X(_06857_));
 sky130_fd_sc_hd__a221o_1 _21482_ (.A1(\line_cache[87][4] ),
    .A2(_05551_),
    .B1(\line_cache[86][4] ),
    .B2(_05529_),
    .C1(_06857_),
    .X(_06858_));
 sky130_fd_sc_hd__a22o_1 _21483_ (.A1(_05553_),
    .A2(\line_cache[88][4] ),
    .B1(_05549_),
    .B2(\line_cache[89][4] ),
    .X(_06859_));
 sky130_fd_sc_hd__a221o_1 _21484_ (.A1(\line_cache[91][4] ),
    .A2(_05525_),
    .B1(\line_cache[90][4] ),
    .B2(_05550_),
    .C1(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__or4_2 _21485_ (.A(_06854_),
    .B(_06856_),
    .C(_06858_),
    .D(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__nor2_1 _21486_ (.A(_06852_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__and3_1 _21487_ (.A(_05207_),
    .B(\line_cache[121][4] ),
    .C(_05562_),
    .X(_06863_));
 sky130_fd_sc_hd__a21o_1 _21488_ (.A1(\line_cache[120][4] ),
    .A2(_05561_),
    .B1(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__a221o_1 _21489_ (.A1(\line_cache[123][4] ),
    .A2(_05591_),
    .B1(\line_cache[122][4] ),
    .B2(_05559_),
    .C1(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__and3_1 _21490_ (.A(_05586_),
    .B(\line_cache[126][4] ),
    .C(_05562_),
    .X(_06866_));
 sky130_fd_sc_hd__a21o_1 _21491_ (.A1(\line_cache[127][4] ),
    .A2(_05596_),
    .B1(_06866_),
    .X(_06867_));
 sky130_fd_sc_hd__a221o_1 _21492_ (.A1(\line_cache[125][4] ),
    .A2(_05589_),
    .B1(\line_cache[124][4] ),
    .B2(_05590_),
    .C1(_06867_),
    .X(_06868_));
 sky130_fd_sc_hd__a22o_1 _21493_ (.A1(_05569_),
    .A2(\line_cache[115][4] ),
    .B1(_05582_),
    .B2(\line_cache[114][4] ),
    .X(_06869_));
 sky130_fd_sc_hd__a221o_1 _21494_ (.A1(\line_cache[113][4] ),
    .A2(_05581_),
    .B1(\line_cache[112][4] ),
    .B2(_05579_),
    .C1(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__a22o_1 _21495_ (.A1(_05568_),
    .A2(\line_cache[116][4] ),
    .B1(_05567_),
    .B2(\line_cache[117][4] ),
    .X(_06871_));
 sky130_fd_sc_hd__a221o_1 _21496_ (.A1(\line_cache[119][4] ),
    .A2(_06088_),
    .B1(\line_cache[118][4] ),
    .B2(_05566_),
    .C1(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__or4_1 _21497_ (.A(_06865_),
    .B(_06868_),
    .C(_06870_),
    .D(_06872_),
    .X(_06873_));
 sky130_fd_sc_hd__a22o_1 _21498_ (.A1(_05376_),
    .A2(\line_cache[140][4] ),
    .B1(_05375_),
    .B2(\line_cache[141][4] ),
    .X(_06874_));
 sky130_fd_sc_hd__a221o_1 _21499_ (.A1(\line_cache[143][4] ),
    .A2(_05382_),
    .B1(\line_cache[142][4] ),
    .B2(_05374_),
    .C1(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__a22o_1 _21500_ (.A1(_05612_),
    .A2(\line_cache[131][4] ),
    .B1(_05598_),
    .B2(\line_cache[130][4] ),
    .X(_06876_));
 sky130_fd_sc_hd__a221o_1 _21501_ (.A1(\line_cache[129][4] ),
    .A2(_05597_),
    .B1(\line_cache[128][4] ),
    .B2(_05594_),
    .C1(_06876_),
    .X(_06877_));
 sky130_fd_sc_hd__and2_1 _21502_ (.A(_05609_),
    .B(\line_cache[133][4] ),
    .X(_06878_));
 sky130_fd_sc_hd__and3_1 _21503_ (.A(_05611_),
    .B(\line_cache[132][4] ),
    .C(_05381_),
    .X(_06879_));
 sky130_fd_sc_hd__or2_1 _21504_ (.A(_06878_),
    .B(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__a221o_1 _21505_ (.A1(\line_cache[135][4] ),
    .A2(_05605_),
    .B1(\line_cache[134][4] ),
    .B2(_05608_),
    .C1(_06880_),
    .X(_06881_));
 sky130_fd_sc_hd__a22o_1 _21506_ (.A1(_05604_),
    .A2(\line_cache[136][4] ),
    .B1(_05603_),
    .B2(\line_cache[137][4] ),
    .X(_06882_));
 sky130_fd_sc_hd__a221o_1 _21507_ (.A1(\line_cache[139][4] ),
    .A2(_05377_),
    .B1(\line_cache[138][4] ),
    .B2(_05602_),
    .C1(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__or4_1 _21508_ (.A(_06875_),
    .B(_06877_),
    .C(_06881_),
    .D(_06883_),
    .X(_06884_));
 sky130_fd_sc_hd__nor2_1 _21509_ (.A(_06873_),
    .B(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__and3_2 _21510_ (.A(_06841_),
    .B(_06862_),
    .C(_06885_),
    .X(_06886_));
 sky130_fd_sc_hd__nand3_1 _21511_ (.A(_06711_),
    .B(_06812_),
    .C(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__o21a_4 _21512_ (.A1(_06643_),
    .A2(_06887_),
    .B1(_05884_),
    .X(net130));
 sky130_fd_sc_hd__nor3b_1 _21513_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][5] ),
    .Y(_06888_));
 sky130_fd_sc_hd__and2_1 _21514_ (.A(_05797_),
    .B(\line_cache[1][5] ),
    .X(_06889_));
 sky130_fd_sc_hd__and3_1 _21515_ (.A(_05779_),
    .B(_05840_),
    .C(\line_cache[2][5] ),
    .X(_06890_));
 sky130_fd_sc_hd__a211o_1 _21516_ (.A1(\line_cache[15][5] ),
    .A2(_05798_),
    .B1(_06889_),
    .C1(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__and3_1 _21517_ (.A(_05778_),
    .B(_05792_),
    .C(\line_cache[3][5] ),
    .X(_06892_));
 sky130_fd_sc_hd__a31o_1 _21518_ (.A1(_05188_),
    .A2(\line_cache[4][5] ),
    .A3(_05771_),
    .B1(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__a221o_1 _21519_ (.A1(_05343_),
    .A2(\line_cache[5][5] ),
    .B1(\line_cache[6][5] ),
    .B2(_05348_),
    .C1(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__and3_1 _21520_ (.A(_05112_),
    .B(_05151_),
    .C(\line_cache[319][5] ),
    .X(_06895_));
 sky130_fd_sc_hd__a32o_1 _21521_ (.A1(_05991_),
    .A2(_05180_),
    .A3(\line_cache[31][5] ),
    .B1(_05998_),
    .B2(\line_cache[47][5] ),
    .X(_06896_));
 sky130_fd_sc_hd__a311o_1 _21522_ (.A1(_05188_),
    .A2(\line_cache[63][5] ),
    .A3(_05112_),
    .B1(_06895_),
    .C1(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__nand2_1 _21523_ (.A(_05787_),
    .B(\line_cache[303][5] ),
    .Y(_06898_));
 sky130_fd_sc_hd__nand2_1 _21524_ (.A(_05791_),
    .B(\line_cache[271][5] ),
    .Y(_06899_));
 sky130_fd_sc_hd__nand2_1 _21525_ (.A(_06898_),
    .B(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__a221oi_4 _21526_ (.A1(\line_cache[255][5] ),
    .A2(_05220_),
    .B1(\line_cache[287][5] ),
    .B2(_05788_),
    .C1(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__or4b_1 _21527_ (.A(_06891_),
    .B(_06894_),
    .C(_06897_),
    .D_N(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__a22o_1 _21528_ (.A1(_05283_),
    .A2(\line_cache[45][5] ),
    .B1(\line_cache[46][5] ),
    .B2(_05285_),
    .X(_06903_));
 sky130_fd_sc_hd__a22o_1 _21529_ (.A1(_05298_),
    .A2(\line_cache[48][5] ),
    .B1(\line_cache[49][5] ),
    .B2(_05300_),
    .X(_06904_));
 sky130_fd_sc_hd__nand2_1 _21530_ (.A(_05279_),
    .B(\line_cache[41][5] ),
    .Y(_06905_));
 sky130_fd_sc_hd__nand2_1 _21531_ (.A(_05281_),
    .B(\line_cache[42][5] ),
    .Y(_06906_));
 sky130_fd_sc_hd__nand2_1 _21532_ (.A(_06905_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__a221oi_1 _21533_ (.A1(_05277_),
    .A2(\line_cache[43][5] ),
    .B1(\line_cache[44][5] ),
    .B2(_05287_),
    .C1(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__or3b_1 _21534_ (.A(_06903_),
    .B(_06904_),
    .C_N(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__a22o_1 _21535_ (.A1(_05106_),
    .A2(\line_cache[317][5] ),
    .B1(\line_cache[316][5] ),
    .B2(_05108_),
    .X(_06910_));
 sky130_fd_sc_hd__a22o_1 _21536_ (.A1(_05292_),
    .A2(\line_cache[61][5] ),
    .B1(\line_cache[60][5] ),
    .B2(_05294_),
    .X(_06911_));
 sky130_fd_sc_hd__a22o_1 _21537_ (.A1(_05312_),
    .A2(\line_cache[58][5] ),
    .B1(_05317_),
    .B2(\line_cache[59][5] ),
    .X(_06912_));
 sky130_fd_sc_hd__and3_1 _21538_ (.A(_05109_),
    .B(_05021_),
    .C(\line_cache[318][5] ),
    .X(_06913_));
 sky130_fd_sc_hd__a21o_1 _21539_ (.A1(\line_cache[62][5] ),
    .A2(_05296_),
    .B1(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__or4_1 _21540_ (.A(_06910_),
    .B(_06911_),
    .C(_06912_),
    .D(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__a22o_1 _21541_ (.A1(_05129_),
    .A2(\line_cache[304][5] ),
    .B1(\line_cache[305][5] ),
    .B2(_05127_),
    .X(_06916_));
 sky130_fd_sc_hd__a22o_1 _21542_ (.A1(_05119_),
    .A2(\line_cache[312][5] ),
    .B1(\line_cache[313][5] ),
    .B2(_05121_),
    .X(_06917_));
 sky130_fd_sc_hd__a22o_1 _21543_ (.A1(_05123_),
    .A2(\line_cache[314][5] ),
    .B1(_05644_),
    .B2(\line_cache[315][5] ),
    .X(_06918_));
 sky130_fd_sc_hd__a22o_1 _21544_ (.A1(_05132_),
    .A2(\line_cache[306][5] ),
    .B1(\line_cache[307][5] ),
    .B2(_05136_),
    .X(_06919_));
 sky130_fd_sc_hd__or4_1 _21545_ (.A(_06916_),
    .B(_06917_),
    .C(_06918_),
    .D(_06919_),
    .X(_06920_));
 sky130_fd_sc_hd__a22o_1 _21546_ (.A1(_05314_),
    .A2(\line_cache[56][5] ),
    .B1(\line_cache[57][5] ),
    .B2(_05315_),
    .X(_06921_));
 sky130_fd_sc_hd__a22o_1 _21547_ (.A1(_05304_),
    .A2(\line_cache[52][5] ),
    .B1(\line_cache[53][5] ),
    .B2(_05306_),
    .X(_06922_));
 sky130_fd_sc_hd__a22o_1 _21548_ (.A1(_05301_),
    .A2(\line_cache[50][5] ),
    .B1(\line_cache[51][5] ),
    .B2(_05302_),
    .X(_06923_));
 sky130_fd_sc_hd__a22o_1 _21549_ (.A1(_05307_),
    .A2(\line_cache[54][5] ),
    .B1(_05309_),
    .B2(\line_cache[55][5] ),
    .X(_06924_));
 sky130_fd_sc_hd__or4_2 _21550_ (.A(_06921_),
    .B(_06922_),
    .C(_06923_),
    .D(_06924_),
    .X(_06925_));
 sky130_fd_sc_hd__or4_1 _21551_ (.A(_06909_),
    .B(_06915_),
    .C(_06920_),
    .D(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__or2b_1 _21552_ (.A(_05365_),
    .B_N(\line_cache[12][5] ),
    .X(_06927_));
 sky130_fd_sc_hd__nand2_1 _21553_ (.A(_05358_),
    .B(\line_cache[11][5] ),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _21554_ (.A(_06927_),
    .B(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__a221oi_1 _21555_ (.A1(\line_cache[14][5] ),
    .A2(_05838_),
    .B1(\line_cache[13][5] ),
    .B2(_05839_),
    .C1(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__nand2_1 _21556_ (.A(_05353_),
    .B(\line_cache[10][5] ),
    .Y(_06931_));
 sky130_fd_sc_hd__nand2_1 _21557_ (.A(_05351_),
    .B(\line_cache[9][5] ),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_1 _21558_ (.A(_06931_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__a221oi_1 _21559_ (.A1(_05355_),
    .A2(\line_cache[8][5] ),
    .B1(_05346_),
    .B2(\line_cache[7][5] ),
    .C1(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__nand2_1 _21560_ (.A(_06930_),
    .B(_06934_),
    .Y(_06935_));
 sky130_fd_sc_hd__and3_1 _21561_ (.A(_05163_),
    .B(_05812_),
    .C(\line_cache[21][5] ),
    .X(_06936_));
 sky130_fd_sc_hd__and3_1 _21562_ (.A(_05167_),
    .B(_05812_),
    .C(\line_cache[20][5] ),
    .X(_06937_));
 sky130_fd_sc_hd__a22o_1 _21563_ (.A1(_05825_),
    .A2(\line_cache[23][5] ),
    .B1(\line_cache[22][5] ),
    .B2(_05826_),
    .X(_06938_));
 sky130_fd_sc_hd__a22o_1 _21564_ (.A1(_05329_),
    .A2(\line_cache[16][5] ),
    .B1(\line_cache[17][5] ),
    .B2(_05330_),
    .X(_06939_));
 sky130_fd_sc_hd__a221o_1 _21565_ (.A1(\line_cache[19][5] ),
    .A2(_05831_),
    .B1(\line_cache[18][5] ),
    .B2(_05832_),
    .C1(_06939_),
    .X(_06940_));
 sky130_fd_sc_hd__or4_1 _21566_ (.A(_06936_),
    .B(_06937_),
    .C(_06938_),
    .D(_06940_),
    .X(_06941_));
 sky130_fd_sc_hd__a22o_1 _21567_ (.A1(_05262_),
    .A2(\line_cache[33][5] ),
    .B1(\line_cache[34][5] ),
    .B2(_05263_),
    .X(_06942_));
 sky130_fd_sc_hd__a221o_1 _21568_ (.A1(\line_cache[36][5] ),
    .A2(_05266_),
    .B1(\line_cache[35][5] ),
    .B2(_05261_),
    .C1(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__and3_1 _21569_ (.A(_05146_),
    .B(_05792_),
    .C(\line_cache[25][5] ),
    .X(_06944_));
 sky130_fd_sc_hd__a31o_1 _21570_ (.A1(_05840_),
    .A2(\line_cache[24][5] ),
    .A3(_05320_),
    .B1(_06944_),
    .X(_06945_));
 sky130_fd_sc_hd__a221oi_2 _21571_ (.A1(\line_cache[27][5] ),
    .A2(_05817_),
    .B1(\line_cache[26][5] ),
    .B2(_05819_),
    .C1(_06945_),
    .Y(_06946_));
 sky130_fd_sc_hd__a32o_1 _21572_ (.A1(_05175_),
    .A2(_05812_),
    .A3(\line_cache[30][5] ),
    .B1(_05260_),
    .B2(\line_cache[32][5] ),
    .X(_06947_));
 sky130_fd_sc_hd__a32o_1 _21573_ (.A1(_05840_),
    .A2(_05173_),
    .A3(\line_cache[29][5] ),
    .B1(_06051_),
    .B2(\line_cache[28][5] ),
    .X(_06948_));
 sky130_fd_sc_hd__nor2_1 _21574_ (.A(_06947_),
    .B(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__nand2_1 _21575_ (.A(_05270_),
    .B(\line_cache[38][5] ),
    .Y(_06950_));
 sky130_fd_sc_hd__nand2_1 _21576_ (.A(_05272_),
    .B(\line_cache[37][5] ),
    .Y(_06951_));
 sky130_fd_sc_hd__nand2_1 _21577_ (.A(_06950_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__a221oi_2 _21578_ (.A1(_05268_),
    .A2(\line_cache[39][5] ),
    .B1(\line_cache[40][5] ),
    .B2(_05275_),
    .C1(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__and4b_1 _21579_ (.A_N(_06943_),
    .B(_06946_),
    .C(_06949_),
    .D(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__or3b_2 _21580_ (.A(_06935_),
    .B(_06941_),
    .C_N(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__nor3_2 _21581_ (.A(_06902_),
    .B(_06926_),
    .C(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__and3_1 _21582_ (.A(_05203_),
    .B(\line_cache[203][5] ),
    .C(_05471_),
    .X(_06957_));
 sky130_fd_sc_hd__and3_1 _21583_ (.A(_05586_),
    .B(\line_cache[206][5] ),
    .C(_05685_),
    .X(_06958_));
 sky130_fd_sc_hd__and2b_1 _21584_ (.A_N(_05687_),
    .B(\line_cache[204][5] ),
    .X(_06959_));
 sky130_fd_sc_hd__a2111o_1 _21585_ (.A1(\line_cache[205][5] ),
    .A2(_05683_),
    .B1(_06957_),
    .C1(_06958_),
    .D1(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__a22o_1 _21586_ (.A1(_05484_),
    .A2(\line_cache[195][5] ),
    .B1(_05485_),
    .B2(\line_cache[196][5] ),
    .X(_06961_));
 sky130_fd_sc_hd__a221o_1 _21587_ (.A1(\line_cache[198][5] ),
    .A2(_05487_),
    .B1(\line_cache[197][5] ),
    .B2(_05489_),
    .C1(_06961_),
    .X(_06962_));
 sky130_fd_sc_hd__a22o_1 _21588_ (.A1(_05495_),
    .A2(\line_cache[200][5] ),
    .B1(_05493_),
    .B2(\line_cache[199][5] ),
    .X(_06963_));
 sky130_fd_sc_hd__a221o_1 _21589_ (.A1(\line_cache[202][5] ),
    .A2(_05492_),
    .B1(\line_cache[201][5] ),
    .B2(_05491_),
    .C1(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__and3_1 _21590_ (.A(_05470_),
    .B(\line_cache[193][5] ),
    .C(_05685_),
    .X(_06965_));
 sky130_fd_sc_hd__and3_1 _21591_ (.A(_05475_),
    .B(\line_cache[192][5] ),
    .C(_05472_),
    .X(_06966_));
 sky130_fd_sc_hd__and3_1 _21592_ (.A(_05409_),
    .B(\line_cache[194][5] ),
    .C(_05472_),
    .X(_06967_));
 sky130_fd_sc_hd__a2111o_1 _21593_ (.A1(_05630_),
    .A2(\line_cache[286][5] ),
    .B1(_06965_),
    .C1(_06966_),
    .D1(_06967_),
    .X(_06968_));
 sky130_fd_sc_hd__or4_1 _21594_ (.A(_06960_),
    .B(_06962_),
    .C(_06964_),
    .D(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__a22o_1 _21595_ (.A1(_05676_),
    .A2(\line_cache[283][5] ),
    .B1(_05678_),
    .B2(\line_cache[282][5] ),
    .X(_06970_));
 sky130_fd_sc_hd__a22o_1 _21596_ (.A1(_05674_),
    .A2(\line_cache[284][5] ),
    .B1(_05631_),
    .B2(\line_cache[285][5] ),
    .X(_06971_));
 sky130_fd_sc_hd__a32o_1 _21597_ (.A1(_05165_),
    .A2(_05059_),
    .A3(\line_cache[278][5] ),
    .B1(_05654_),
    .B2(\line_cache[279][5] ),
    .X(_06972_));
 sky130_fd_sc_hd__a221o_1 _21598_ (.A1(\line_cache[281][5] ),
    .A2(_05677_),
    .B1(\line_cache[280][5] ),
    .B2(_05144_),
    .C1(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__a22o_1 _21599_ (.A1(_05668_),
    .A2(\line_cache[270][5] ),
    .B1(\line_cache[269][5] ),
    .B2(_05670_),
    .X(_06974_));
 sky130_fd_sc_hd__a22o_1 _21600_ (.A1(_05659_),
    .A2(\line_cache[275][5] ),
    .B1(\line_cache[274][5] ),
    .B2(_05662_),
    .X(_06975_));
 sky130_fd_sc_hd__a22o_1 _21601_ (.A1(_05658_),
    .A2(\line_cache[276][5] ),
    .B1(\line_cache[277][5] ),
    .B2(_05655_),
    .X(_06976_));
 sky130_fd_sc_hd__a22o_1 _21602_ (.A1(_05666_),
    .A2(\line_cache[272][5] ),
    .B1(\line_cache[273][5] ),
    .B2(_05660_),
    .X(_06977_));
 sky130_fd_sc_hd__or4_1 _21603_ (.A(_06974_),
    .B(_06975_),
    .C(_06976_),
    .D(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__or4_1 _21604_ (.A(_06970_),
    .B(_06971_),
    .C(_06973_),
    .D(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__nor2_1 _21605_ (.A(_06969_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__a22o_1 _21606_ (.A1(_05746_),
    .A2(\line_cache[236][5] ),
    .B1(_05747_),
    .B2(\line_cache[235][5] ),
    .X(_06981_));
 sky130_fd_sc_hd__a221o_1 _21607_ (.A1(\line_cache[238][5] ),
    .A2(_05744_),
    .B1(\line_cache[237][5] ),
    .B2(_05745_),
    .C1(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__and3_1 _21608_ (.A(_05469_),
    .B(\line_cache[225][5] ),
    .C(_05732_),
    .X(_06983_));
 sky130_fd_sc_hd__and3_1 _21609_ (.A(_05408_),
    .B(\line_cache[226][5] ),
    .C(_05721_),
    .X(_06984_));
 sky130_fd_sc_hd__and3_1 _21610_ (.A(_05475_),
    .B(\line_cache[224][5] ),
    .C(_05194_),
    .X(_06985_));
 sky130_fd_sc_hd__a2111o_1 _21611_ (.A1(\line_cache[223][5] ),
    .A2(_05720_),
    .B1(_06983_),
    .C1(_06984_),
    .D1(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__and3_1 _21612_ (.A(_05704_),
    .B(\line_cache[227][5] ),
    .C(_05193_),
    .X(_06987_));
 sky130_fd_sc_hd__and3_1 _21613_ (.A(_05610_),
    .B(\line_cache[228][5] ),
    .C(_05193_),
    .X(_06988_));
 sky130_fd_sc_hd__and3_1 _21614_ (.A(_05710_),
    .B(\line_cache[229][5] ),
    .C(_05193_),
    .X(_06989_));
 sky130_fd_sc_hd__and3_1 _21615_ (.A(_05708_),
    .B(\line_cache[230][5] ),
    .C(_05732_),
    .X(_06990_));
 sky130_fd_sc_hd__or4_1 _21616_ (.A(_06987_),
    .B(_06988_),
    .C(_06989_),
    .D(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__a22o_1 _21617_ (.A1(_05728_),
    .A2(\line_cache[232][5] ),
    .B1(_05729_),
    .B2(\line_cache[231][5] ),
    .X(_06992_));
 sky130_fd_sc_hd__a221o_1 _21618_ (.A1(\line_cache[234][5] ),
    .A2(_05726_),
    .B1(\line_cache[233][5] ),
    .B2(_05727_),
    .C1(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__or4_1 _21619_ (.A(_06982_),
    .B(_06986_),
    .C(_06991_),
    .D(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__a22o_1 _21620_ (.A1(_05716_),
    .A2(\line_cache[220][5] ),
    .B1(_05717_),
    .B2(\line_cache[219][5] ),
    .X(_06995_));
 sky130_fd_sc_hd__a221o_1 _21621_ (.A1(\line_cache[222][5] ),
    .A2(_05714_),
    .B1(\line_cache[221][5] ),
    .B2(_05715_),
    .C1(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__a22o_1 _21622_ (.A1(_05700_),
    .A2(\line_cache[209][5] ),
    .B1(\line_cache[210][5] ),
    .B2(_05701_),
    .X(_06997_));
 sky130_fd_sc_hd__a221o_1 _21623_ (.A1(\line_cache[208][5] ),
    .A2(_05698_),
    .B1(\line_cache[207][5] ),
    .B2(_05699_),
    .C1(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__and3_1 _21624_ (.A(_05704_),
    .B(\line_cache[211][5] ),
    .C(_05693_),
    .X(_06999_));
 sky130_fd_sc_hd__and3_1 _21625_ (.A(_05610_),
    .B(\line_cache[212][5] ),
    .C(_05694_),
    .X(_07000_));
 sky130_fd_sc_hd__and3_1 _21626_ (.A(_05710_),
    .B(\line_cache[213][5] ),
    .C(_05694_),
    .X(_07001_));
 sky130_fd_sc_hd__and3_1 _21627_ (.A(_05708_),
    .B(\line_cache[214][5] ),
    .C(_05706_),
    .X(_07002_));
 sky130_fd_sc_hd__or4_2 _21628_ (.A(_06999_),
    .B(_07000_),
    .C(_07001_),
    .D(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__a22o_1 _21629_ (.A1(_05692_),
    .A2(\line_cache[216][5] ),
    .B1(_05983_),
    .B2(\line_cache[215][5] ),
    .X(_07004_));
 sky130_fd_sc_hd__a221o_1 _21630_ (.A1(\line_cache[218][5] ),
    .A2(_05690_),
    .B1(\line_cache[217][5] ),
    .B2(_05691_),
    .C1(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__or4_2 _21631_ (.A(_06996_),
    .B(_06998_),
    .C(_07003_),
    .D(_07005_),
    .X(_07006_));
 sky130_fd_sc_hd__and3_1 _21632_ (.A(_05454_),
    .B(\line_cache[239][5] ),
    .C(_05192_),
    .X(_07007_));
 sky130_fd_sc_hd__and3_1 _21633_ (.A(_05469_),
    .B(\line_cache[241][5] ),
    .C(_05198_),
    .X(_07008_));
 sky130_fd_sc_hd__and3_1 _21634_ (.A(_05407_),
    .B(\line_cache[242][5] ),
    .C(_05198_),
    .X(_07009_));
 sky130_fd_sc_hd__a2111o_1 _21635_ (.A1(_05233_),
    .A2(\line_cache[240][5] ),
    .B1(_07007_),
    .C1(_07008_),
    .D1(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__and2_1 _21636_ (.A(_05235_),
    .B(\line_cache[243][5] ),
    .X(_07011_));
 sky130_fd_sc_hd__a21o_1 _21637_ (.A1(\line_cache[244][5] ),
    .A2(_05224_),
    .B1(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__a221o_1 _21638_ (.A1(\line_cache[246][5] ),
    .A2(_05753_),
    .B1(\line_cache[245][5] ),
    .B2(_05226_),
    .C1(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__a22o_1 _21639_ (.A1(_05212_),
    .A2(\line_cache[252][5] ),
    .B1(_05205_),
    .B2(\line_cache[251][5] ),
    .X(_07014_));
 sky130_fd_sc_hd__a221o_1 _21640_ (.A1(\line_cache[254][5] ),
    .A2(_05217_),
    .B1(\line_cache[253][5] ),
    .B2(_05214_),
    .C1(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__a22o_1 _21641_ (.A1(_05750_),
    .A2(\line_cache[248][5] ),
    .B1(_05229_),
    .B2(\line_cache[247][5] ),
    .X(_07016_));
 sky130_fd_sc_hd__a221o_1 _21642_ (.A1(\line_cache[250][5] ),
    .A2(_05202_),
    .B1(\line_cache[249][5] ),
    .B2(_05209_),
    .C1(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__or4_1 _21643_ (.A(_07010_),
    .B(_07013_),
    .C(_07015_),
    .D(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__a22o_1 _21644_ (.A1(_05545_),
    .A2(\line_cache[78][5] ),
    .B1(_05537_),
    .B2(\line_cache[79][5] ),
    .X(_07019_));
 sky130_fd_sc_hd__a32o_1 _21645_ (.A1(_05544_),
    .A2(\line_cache[77][5] ),
    .A3(_05536_),
    .B1(\line_cache[76][5] ),
    .B2(_05542_),
    .X(_07020_));
 sky130_fd_sc_hd__or2_1 _21646_ (.A(_07019_),
    .B(_07020_),
    .X(_07021_));
 sky130_fd_sc_hd__and2_1 _21647_ (.A(_05860_),
    .B(\line_cache[65][5] ),
    .X(_07022_));
 sky130_fd_sc_hd__a21o_1 _21648_ (.A1(_05858_),
    .A2(\line_cache[64][5] ),
    .B1(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__a221o_1 _21649_ (.A1(\line_cache[67][5] ),
    .A2(_05875_),
    .B1(\line_cache[66][5] ),
    .B2(_05861_),
    .C1(_07023_),
    .X(_07024_));
 sky130_fd_sc_hd__a22o_1 _21650_ (.A1(_05867_),
    .A2(\line_cache[72][5] ),
    .B1(_05866_),
    .B2(\line_cache[73][5] ),
    .X(_07025_));
 sky130_fd_sc_hd__a221o_1 _21651_ (.A1(\line_cache[75][5] ),
    .A2(_05543_),
    .B1(\line_cache[74][5] ),
    .B2(_05865_),
    .C1(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__a22o_1 _21652_ (.A1(_05873_),
    .A2(\line_cache[68][5] ),
    .B1(_05872_),
    .B2(\line_cache[69][5] ),
    .X(_07027_));
 sky130_fd_sc_hd__a221o_1 _21653_ (.A1(\line_cache[71][5] ),
    .A2(_05868_),
    .B1(\line_cache[70][5] ),
    .B2(_05871_),
    .C1(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__or4_4 _21654_ (.A(_07021_),
    .B(_07024_),
    .C(_07026_),
    .D(_07028_),
    .X(_07029_));
 sky130_fd_sc_hd__or2_1 _21655_ (.A(_07018_),
    .B(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__nor3_1 _21656_ (.A(_06994_),
    .B(_07006_),
    .C(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__and3_1 _21657_ (.A(_05058_),
    .B(_05034_),
    .C(\line_cache[302][5] ),
    .X(_07032_));
 sky130_fd_sc_hd__a22o_1 _21658_ (.A1(_05056_),
    .A2(\line_cache[301][5] ),
    .B1(\line_cache[300][5] ),
    .B2(_05053_),
    .X(_07033_));
 sky130_fd_sc_hd__a211o_1 _21659_ (.A1(\line_cache[256][5] ),
    .A2(_05777_),
    .B1(_07032_),
    .C1(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__and3_1 _21660_ (.A(_05779_),
    .B(_05021_),
    .C(\line_cache[258][5] ),
    .X(_07035_));
 sky130_fd_sc_hd__and3_1 _21661_ (.A(_05771_),
    .B(_05034_),
    .C(\line_cache[260][5] ),
    .X(_07036_));
 sky130_fd_sc_hd__and3_1 _21662_ (.A(_05778_),
    .B(_05034_),
    .C(\line_cache[259][5] ),
    .X(_07037_));
 sky130_fd_sc_hd__a2111o_1 _21663_ (.A1(\line_cache[257][5] ),
    .A2(_05776_),
    .B1(_07035_),
    .C1(_07036_),
    .D1(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__and3_1 _21664_ (.A(_05356_),
    .B(_05034_),
    .C(\line_cache[267][5] ),
    .X(_07039_));
 sky130_fd_sc_hd__a22o_1 _21665_ (.A1(_05760_),
    .A2(\line_cache[266][5] ),
    .B1(\line_cache[265][5] ),
    .B2(_05764_),
    .X(_07040_));
 sky130_fd_sc_hd__a311o_1 _21666_ (.A1(_05113_),
    .A2(\line_cache[268][5] ),
    .A3(_05364_),
    .B1(_07039_),
    .C1(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__nand2_1 _21667_ (.A(_05768_),
    .B(\line_cache[262][5] ),
    .Y(_07042_));
 sky130_fd_sc_hd__nand2_1 _21668_ (.A(_05773_),
    .B(\line_cache[261][5] ),
    .Y(_07043_));
 sky130_fd_sc_hd__nand2_1 _21669_ (.A(_07042_),
    .B(_07043_),
    .Y(_07044_));
 sky130_fd_sc_hd__a221oi_1 _21670_ (.A1(_05763_),
    .A2(\line_cache[264][5] ),
    .B1(_05770_),
    .B2(\line_cache[263][5] ),
    .C1(_07044_),
    .Y(_07045_));
 sky130_fd_sc_hd__or4b_1 _21671_ (.A(_07034_),
    .B(_07038_),
    .C(_07041_),
    .D_N(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__a22o_1 _21672_ (.A1(_05098_),
    .A2(\line_cache[308][5] ),
    .B1(\line_cache[309][5] ),
    .B2(_05093_),
    .X(_07047_));
 sky130_fd_sc_hd__a221o_1 _21673_ (.A1(\line_cache[311][5] ),
    .A2(_05097_),
    .B1(\line_cache[310][5] ),
    .B2(_05103_),
    .C1(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__a22o_1 _21674_ (.A1(_05046_),
    .A2(\line_cache[295][5] ),
    .B1(\line_cache[294][5] ),
    .B2(_05043_),
    .X(_07049_));
 sky130_fd_sc_hd__a221o_1 _21675_ (.A1(\line_cache[293][5] ),
    .A2(_05628_),
    .B1(\line_cache[292][5] ),
    .B2(_05627_),
    .C1(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__a22o_1 _21676_ (.A1(_05069_),
    .A2(\line_cache[296][5] ),
    .B1(\line_cache[297][5] ),
    .B2(_05076_),
    .X(_07051_));
 sky130_fd_sc_hd__a221o_1 _21677_ (.A1(\line_cache[299][5] ),
    .A2(_05073_),
    .B1(\line_cache[298][5] ),
    .B2(_05079_),
    .C1(_07051_),
    .X(_07052_));
 sky130_fd_sc_hd__a22o_1 _21678_ (.A1(_05632_),
    .A2(\line_cache[288][5] ),
    .B1(\line_cache[289][5] ),
    .B2(_05633_),
    .X(_07053_));
 sky130_fd_sc_hd__a221o_1 _21679_ (.A1(\line_cache[291][5] ),
    .A2(_05623_),
    .B1(\line_cache[290][5] ),
    .B2(_05624_),
    .C1(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__or4_2 _21680_ (.A(_07048_),
    .B(_07050_),
    .C(_07052_),
    .D(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__nor2_1 _21681_ (.A(_07046_),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__and3_2 _21682_ (.A(_06980_),
    .B(_07031_),
    .C(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__and3_1 _21683_ (.A(_05227_),
    .B(\line_cache[87][5] ),
    .C(_05518_),
    .X(_07058_));
 sky130_fd_sc_hd__a21o_1 _21684_ (.A1(\line_cache[86][5] ),
    .A2(_05529_),
    .B1(_07058_),
    .X(_07059_));
 sky130_fd_sc_hd__a221o_1 _21685_ (.A1(\line_cache[85][5] ),
    .A2(_05530_),
    .B1(\line_cache[84][5] ),
    .B2(_05532_),
    .C1(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__a22o_1 _21686_ (.A1(_05531_),
    .A2(\line_cache[83][5] ),
    .B1(_05539_),
    .B2(\line_cache[82][5] ),
    .X(_07061_));
 sky130_fd_sc_hd__a221o_1 _21687_ (.A1(\line_cache[81][5] ),
    .A2(_05538_),
    .B1(\line_cache[80][5] ),
    .B2(_05535_),
    .C1(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__a22o_1 _21688_ (.A1(_05524_),
    .A2(\line_cache[92][5] ),
    .B1(_05523_),
    .B2(\line_cache[93][5] ),
    .X(_07063_));
 sky130_fd_sc_hd__a221o_1 _21689_ (.A1(\line_cache[95][5] ),
    .A2(_05519_),
    .B1(\line_cache[94][5] ),
    .B2(_05522_),
    .C1(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__a22o_1 _21690_ (.A1(_05553_),
    .A2(\line_cache[88][5] ),
    .B1(_05549_),
    .B2(\line_cache[89][5] ),
    .X(_07065_));
 sky130_fd_sc_hd__a221o_1 _21691_ (.A1(\line_cache[91][5] ),
    .A2(_05525_),
    .B1(\line_cache[90][5] ),
    .B2(_05550_),
    .C1(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__or4_1 _21692_ (.A(_07060_),
    .B(_07062_),
    .C(_07064_),
    .D(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__a22o_1 _21693_ (.A1(_05510_),
    .A2(\line_cache[99][5] ),
    .B1(_05516_),
    .B2(\line_cache[98][5] ),
    .X(_07068_));
 sky130_fd_sc_hd__a221o_1 _21694_ (.A1(\line_cache[97][5] ),
    .A2(_05515_),
    .B1(\line_cache[96][5] ),
    .B2(_05520_),
    .C1(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__a22o_1 _21695_ (.A1(_05575_),
    .A2(\line_cache[108][5] ),
    .B1(_05574_),
    .B2(\line_cache[109][5] ),
    .X(_07070_));
 sky130_fd_sc_hd__a221o_1 _21696_ (.A1(\line_cache[111][5] ),
    .A2(_05580_),
    .B1(\line_cache[110][5] ),
    .B2(_05573_),
    .C1(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__and2_1 _21697_ (.A(_05502_),
    .B(\line_cache[102][5] ),
    .X(_07072_));
 sky130_fd_sc_hd__a21o_1 _21698_ (.A1(\line_cache[103][5] ),
    .A2(_05504_),
    .B1(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__a221o_1 _21699_ (.A1(\line_cache[101][5] ),
    .A2(_05509_),
    .B1(\line_cache[100][5] ),
    .B2(_05511_),
    .C1(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__a22o_1 _21700_ (.A1(_05503_),
    .A2(\line_cache[104][5] ),
    .B1(_05508_),
    .B2(\line_cache[105][5] ),
    .X(_07075_));
 sky130_fd_sc_hd__a221o_1 _21701_ (.A1(\line_cache[107][5] ),
    .A2(_05576_),
    .B1(\line_cache[106][5] ),
    .B2(_05506_),
    .C1(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__or4_1 _21702_ (.A(_07069_),
    .B(_07071_),
    .C(_07074_),
    .D(_07076_),
    .X(_07077_));
 sky130_fd_sc_hd__nor2_1 _21703_ (.A(_07067_),
    .B(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__and3_1 _21704_ (.A(_05207_),
    .B(\line_cache[137][5] ),
    .C(_05381_),
    .X(_07079_));
 sky130_fd_sc_hd__a21o_1 _21705_ (.A1(\line_cache[136][5] ),
    .A2(_05604_),
    .B1(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__a221o_1 _21706_ (.A1(\line_cache[139][5] ),
    .A2(_05377_),
    .B1(\line_cache[138][5] ),
    .B2(_05602_),
    .C1(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__a22o_1 _21707_ (.A1(_05376_),
    .A2(\line_cache[140][5] ),
    .B1(_05375_),
    .B2(\line_cache[141][5] ),
    .X(_07082_));
 sky130_fd_sc_hd__a221o_1 _21708_ (.A1(\line_cache[143][5] ),
    .A2(_05382_),
    .B1(\line_cache[142][5] ),
    .B2(_05374_),
    .C1(_07082_),
    .X(_07083_));
 sky130_fd_sc_hd__a22o_1 _21709_ (.A1(_05612_),
    .A2(\line_cache[131][5] ),
    .B1(_05598_),
    .B2(\line_cache[130][5] ),
    .X(_07084_));
 sky130_fd_sc_hd__a221o_1 _21710_ (.A1(\line_cache[129][5] ),
    .A2(_05597_),
    .B1(\line_cache[128][5] ),
    .B2(_05594_),
    .C1(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__and2_1 _21711_ (.A(_05609_),
    .B(\line_cache[133][5] ),
    .X(_07086_));
 sky130_fd_sc_hd__and3_1 _21712_ (.A(_05611_),
    .B(\line_cache[132][5] ),
    .C(_05381_),
    .X(_07087_));
 sky130_fd_sc_hd__or2_1 _21713_ (.A(_07086_),
    .B(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__a221o_1 _21714_ (.A1(\line_cache[135][5] ),
    .A2(_05605_),
    .B1(\line_cache[134][5] ),
    .B2(_05608_),
    .C1(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__or4_1 _21715_ (.A(_07081_),
    .B(_07083_),
    .C(_07085_),
    .D(_07089_),
    .X(_07090_));
 sky130_fd_sc_hd__and3_1 _21716_ (.A(_05586_),
    .B(\line_cache[126][5] ),
    .C(_05562_),
    .X(_07091_));
 sky130_fd_sc_hd__a21o_1 _21717_ (.A1(\line_cache[127][5] ),
    .A2(_05596_),
    .B1(_07091_),
    .X(_07092_));
 sky130_fd_sc_hd__a221o_1 _21718_ (.A1(\line_cache[125][5] ),
    .A2(_05589_),
    .B1(\line_cache[124][5] ),
    .B2(_05590_),
    .C1(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__a22o_1 _21719_ (.A1(_05569_),
    .A2(\line_cache[115][5] ),
    .B1(_05582_),
    .B2(\line_cache[114][5] ),
    .X(_07094_));
 sky130_fd_sc_hd__a221o_1 _21720_ (.A1(\line_cache[113][5] ),
    .A2(_05581_),
    .B1(\line_cache[112][5] ),
    .B2(_05579_),
    .C1(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__a22o_1 _21721_ (.A1(_05568_),
    .A2(\line_cache[116][5] ),
    .B1(_05567_),
    .B2(\line_cache[117][5] ),
    .X(_07096_));
 sky130_fd_sc_hd__a221o_1 _21722_ (.A1(\line_cache[119][5] ),
    .A2(_06088_),
    .B1(\line_cache[118][5] ),
    .B2(_05566_),
    .C1(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__a22o_1 _21723_ (.A1(_05561_),
    .A2(\line_cache[120][5] ),
    .B1(_05560_),
    .B2(\line_cache[121][5] ),
    .X(_07098_));
 sky130_fd_sc_hd__a221o_1 _21724_ (.A1(\line_cache[123][5] ),
    .A2(_05591_),
    .B1(\line_cache[122][5] ),
    .B2(_05559_),
    .C1(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__or4_1 _21725_ (.A(_07093_),
    .B(_07095_),
    .C(_07097_),
    .D(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__nor2_1 _21726_ (.A(_07090_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__a22o_1 _21727_ (.A1(_05419_),
    .A2(\line_cache[155][5] ),
    .B1(\line_cache[154][5] ),
    .B2(_06107_),
    .X(_07102_));
 sky130_fd_sc_hd__a221o_1 _21728_ (.A1(\line_cache[153][5] ),
    .A2(_05399_),
    .B1(\line_cache[152][5] ),
    .B2(_05397_),
    .C1(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__a22o_1 _21729_ (.A1(_05392_),
    .A2(\line_cache[147][5] ),
    .B1(_05386_),
    .B2(\line_cache[146][5] ),
    .X(_07104_));
 sky130_fd_sc_hd__a221oi_2 _21730_ (.A1(\line_cache[145][5] ),
    .A2(_05384_),
    .B1(\line_cache[144][5] ),
    .B2(_05380_),
    .C1(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__a22o_1 _21731_ (.A1(_05393_),
    .A2(\line_cache[148][5] ),
    .B1(\line_cache[149][5] ),
    .B2(_05391_),
    .X(_07106_));
 sky130_fd_sc_hd__a221oi_2 _21732_ (.A1(\line_cache[151][5] ),
    .A2(_05398_),
    .B1(\line_cache[150][5] ),
    .B2(_05390_),
    .C1(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__a22o_1 _21733_ (.A1(_05418_),
    .A2(\line_cache[156][5] ),
    .B1(_05417_),
    .B2(\line_cache[157][5] ),
    .X(_07108_));
 sky130_fd_sc_hd__a221oi_1 _21734_ (.A1(\line_cache[159][5] ),
    .A2(_05413_),
    .B1(\line_cache[158][5] ),
    .B2(_05416_),
    .C1(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__and4b_1 _21735_ (.A_N(_07103_),
    .B(_07105_),
    .C(_07107_),
    .D(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__a22o_1 _21736_ (.A1(_05438_),
    .A2(\line_cache[184][5] ),
    .B1(_05440_),
    .B2(\line_cache[185][5] ),
    .X(_07111_));
 sky130_fd_sc_hd__a221o_1 _21737_ (.A1(\line_cache[187][5] ),
    .A2(_05481_),
    .B1(\line_cache[186][5] ),
    .B2(_06131_),
    .C1(_07111_),
    .X(_07112_));
 sky130_fd_sc_hd__a22o_1 _21738_ (.A1(_05449_),
    .A2(\line_cache[180][5] ),
    .B1(_05446_),
    .B2(\line_cache[181][5] ),
    .X(_07113_));
 sky130_fd_sc_hd__a221oi_4 _21739_ (.A1(\line_cache[183][5] ),
    .A2(_05439_),
    .B1(\line_cache[182][5] ),
    .B2(_05445_),
    .C1(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__a22o_1 _21740_ (.A1(_05447_),
    .A2(\line_cache[179][5] ),
    .B1(\line_cache[178][5] ),
    .B2(_05458_),
    .X(_07115_));
 sky130_fd_sc_hd__a221oi_1 _21741_ (.A1(\line_cache[177][5] ),
    .A2(_05457_),
    .B1(\line_cache[176][5] ),
    .B2(_05453_),
    .C1(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__a22o_1 _21742_ (.A1(_05480_),
    .A2(\line_cache[188][5] ),
    .B1(_05479_),
    .B2(\line_cache[189][5] ),
    .X(_07117_));
 sky130_fd_sc_hd__a221oi_2 _21743_ (.A1(\line_cache[191][5] ),
    .A2(_05468_),
    .B1(\line_cache[190][5] ),
    .B2(_05478_),
    .C1(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__and4b_1 _21744_ (.A_N(_07112_),
    .B(_07114_),
    .C(_07116_),
    .D(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__a32o_1 _21745_ (.A1(_05409_),
    .A2(\line_cache[162][5] ),
    .A3(_05410_),
    .B1(\line_cache[163][5] ),
    .B2(_05433_),
    .X(_07120_));
 sky130_fd_sc_hd__a221oi_1 _21746_ (.A1(\line_cache[161][5] ),
    .A2(_05406_),
    .B1(\line_cache[160][5] ),
    .B2(_05414_),
    .C1(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__a22o_1 _21747_ (.A1(_05434_),
    .A2(\line_cache[164][5] ),
    .B1(\line_cache[165][5] ),
    .B2(_05432_),
    .X(_07122_));
 sky130_fd_sc_hd__a221oi_2 _21748_ (.A1(\line_cache[167][5] ),
    .A2(_05425_),
    .B1(\line_cache[166][5] ),
    .B2(_05431_),
    .C1(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__a22o_1 _21749_ (.A1(_05427_),
    .A2(\line_cache[168][5] ),
    .B1(_05423_),
    .B2(\line_cache[169][5] ),
    .X(_07124_));
 sky130_fd_sc_hd__a221oi_2 _21750_ (.A1(\line_cache[171][5] ),
    .A2(_05464_),
    .B1(\line_cache[170][5] ),
    .B2(_05424_),
    .C1(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__nand2_1 _21751_ (.A(_05462_),
    .B(\line_cache[173][5] ),
    .Y(_07126_));
 sky130_fd_sc_hd__nand2_1 _21752_ (.A(_05463_),
    .B(\line_cache[172][5] ),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_1 _21753_ (.A(_07126_),
    .B(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__a221oi_1 _21754_ (.A1(_05461_),
    .A2(\line_cache[174][5] ),
    .B1(_05456_),
    .B2(\line_cache[175][5] ),
    .C1(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__and4_2 _21755_ (.A(_07121_),
    .B(_07123_),
    .C(_07125_),
    .D(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__and3_1 _21756_ (.A(_07110_),
    .B(_07119_),
    .C(_07130_),
    .X(_07131_));
 sky130_fd_sc_hd__and3_1 _21757_ (.A(_07078_),
    .B(_07101_),
    .C(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__nand3_1 _21758_ (.A(_06956_),
    .B(_07057_),
    .C(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__o21a_4 _21759_ (.A1(_06888_),
    .A2(_07133_),
    .B1(_05884_),
    .X(net131));
 sky130_fd_sc_hd__nor3b_1 _21760_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][6] ),
    .Y(_07134_));
 sky130_fd_sc_hd__and2_1 _21761_ (.A(_05797_),
    .B(\line_cache[1][6] ),
    .X(_07135_));
 sky130_fd_sc_hd__and3_1 _21762_ (.A(_05779_),
    .B(_05840_),
    .C(\line_cache[2][6] ),
    .X(_07136_));
 sky130_fd_sc_hd__a211o_1 _21763_ (.A1(\line_cache[15][6] ),
    .A2(_05798_),
    .B1(_07135_),
    .C1(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__and3_1 _21764_ (.A(_05778_),
    .B(_05792_),
    .C(\line_cache[3][6] ),
    .X(_07138_));
 sky130_fd_sc_hd__a31o_1 _21765_ (.A1(_05188_),
    .A2(\line_cache[4][6] ),
    .A3(_05771_),
    .B1(_07138_),
    .X(_07139_));
 sky130_fd_sc_hd__a221o_1 _21766_ (.A1(_05343_),
    .A2(\line_cache[5][6] ),
    .B1(\line_cache[6][6] ),
    .B2(_05348_),
    .C1(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__and3_1 _21767_ (.A(_05112_),
    .B(_05151_),
    .C(\line_cache[319][6] ),
    .X(_07141_));
 sky130_fd_sc_hd__a32o_1 _21768_ (.A1(_05991_),
    .A2(_05180_),
    .A3(\line_cache[31][6] ),
    .B1(_05998_),
    .B2(\line_cache[47][6] ),
    .X(_07142_));
 sky130_fd_sc_hd__a311o_1 _21769_ (.A1(_05188_),
    .A2(\line_cache[63][6] ),
    .A3(_05112_),
    .B1(_07141_),
    .C1(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__nand2_1 _21770_ (.A(_05787_),
    .B(\line_cache[303][6] ),
    .Y(_07144_));
 sky130_fd_sc_hd__nand2_1 _21771_ (.A(_05791_),
    .B(\line_cache[271][6] ),
    .Y(_07145_));
 sky130_fd_sc_hd__nand2_1 _21772_ (.A(_07144_),
    .B(_07145_),
    .Y(_07146_));
 sky130_fd_sc_hd__a221oi_4 _21773_ (.A1(\line_cache[255][6] ),
    .A2(_05220_),
    .B1(\line_cache[287][6] ),
    .B2(_05788_),
    .C1(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__or4b_1 _21774_ (.A(_07137_),
    .B(_07140_),
    .C(_07143_),
    .D_N(_07147_),
    .X(_07148_));
 sky130_fd_sc_hd__a22o_1 _21775_ (.A1(_05283_),
    .A2(\line_cache[45][6] ),
    .B1(\line_cache[46][6] ),
    .B2(_05285_),
    .X(_07149_));
 sky130_fd_sc_hd__a22o_1 _21776_ (.A1(_05298_),
    .A2(\line_cache[48][6] ),
    .B1(\line_cache[49][6] ),
    .B2(_05300_),
    .X(_07150_));
 sky130_fd_sc_hd__nand2_1 _21777_ (.A(_05279_),
    .B(\line_cache[41][6] ),
    .Y(_07151_));
 sky130_fd_sc_hd__nand2_1 _21778_ (.A(_05281_),
    .B(\line_cache[42][6] ),
    .Y(_07152_));
 sky130_fd_sc_hd__nand2_1 _21779_ (.A(_07151_),
    .B(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__a221oi_1 _21780_ (.A1(_05277_),
    .A2(\line_cache[43][6] ),
    .B1(\line_cache[44][6] ),
    .B2(_05287_),
    .C1(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__or3b_1 _21781_ (.A(_07149_),
    .B(_07150_),
    .C_N(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__a22o_1 _21782_ (.A1(_05106_),
    .A2(\line_cache[317][6] ),
    .B1(\line_cache[316][6] ),
    .B2(_05108_),
    .X(_07156_));
 sky130_fd_sc_hd__a22o_1 _21783_ (.A1(_05292_),
    .A2(\line_cache[61][6] ),
    .B1(\line_cache[60][6] ),
    .B2(_05294_),
    .X(_07157_));
 sky130_fd_sc_hd__a22o_1 _21784_ (.A1(_05312_),
    .A2(\line_cache[58][6] ),
    .B1(_05317_),
    .B2(\line_cache[59][6] ),
    .X(_07158_));
 sky130_fd_sc_hd__and3_1 _21785_ (.A(_05109_),
    .B(_05021_),
    .C(\line_cache[318][6] ),
    .X(_07159_));
 sky130_fd_sc_hd__a21o_1 _21786_ (.A1(\line_cache[62][6] ),
    .A2(_05296_),
    .B1(_07159_),
    .X(_07160_));
 sky130_fd_sc_hd__or4_1 _21787_ (.A(_07156_),
    .B(_07157_),
    .C(_07158_),
    .D(_07160_),
    .X(_07161_));
 sky130_fd_sc_hd__a22o_1 _21788_ (.A1(_05129_),
    .A2(\line_cache[304][6] ),
    .B1(\line_cache[305][6] ),
    .B2(_05127_),
    .X(_07162_));
 sky130_fd_sc_hd__a22o_1 _21789_ (.A1(_05119_),
    .A2(\line_cache[312][6] ),
    .B1(\line_cache[313][6] ),
    .B2(_05121_),
    .X(_07163_));
 sky130_fd_sc_hd__a22o_1 _21790_ (.A1(_05123_),
    .A2(\line_cache[314][6] ),
    .B1(_05644_),
    .B2(\line_cache[315][6] ),
    .X(_07164_));
 sky130_fd_sc_hd__a22o_1 _21791_ (.A1(_05132_),
    .A2(\line_cache[306][6] ),
    .B1(\line_cache[307][6] ),
    .B2(_05136_),
    .X(_07165_));
 sky130_fd_sc_hd__or4_2 _21792_ (.A(_07162_),
    .B(_07163_),
    .C(_07164_),
    .D(_07165_),
    .X(_07166_));
 sky130_fd_sc_hd__a22o_1 _21793_ (.A1(_05314_),
    .A2(\line_cache[56][6] ),
    .B1(\line_cache[57][6] ),
    .B2(_05315_),
    .X(_07167_));
 sky130_fd_sc_hd__a22o_1 _21794_ (.A1(_05304_),
    .A2(\line_cache[52][6] ),
    .B1(\line_cache[53][6] ),
    .B2(_05306_),
    .X(_07168_));
 sky130_fd_sc_hd__a22o_1 _21795_ (.A1(_05301_),
    .A2(\line_cache[50][6] ),
    .B1(\line_cache[51][6] ),
    .B2(_05302_),
    .X(_07169_));
 sky130_fd_sc_hd__a22o_1 _21796_ (.A1(_05307_),
    .A2(\line_cache[54][6] ),
    .B1(_05309_),
    .B2(\line_cache[55][6] ),
    .X(_07170_));
 sky130_fd_sc_hd__or4_1 _21797_ (.A(_07167_),
    .B(_07168_),
    .C(_07169_),
    .D(_07170_),
    .X(_07171_));
 sky130_fd_sc_hd__or4_1 _21798_ (.A(_07155_),
    .B(_07161_),
    .C(_07166_),
    .D(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__or2b_1 _21799_ (.A(_05365_),
    .B_N(\line_cache[12][6] ),
    .X(_07173_));
 sky130_fd_sc_hd__nand2_1 _21800_ (.A(_05358_),
    .B(\line_cache[11][6] ),
    .Y(_07174_));
 sky130_fd_sc_hd__nand2_1 _21801_ (.A(_07173_),
    .B(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__a221oi_1 _21802_ (.A1(\line_cache[14][6] ),
    .A2(_05838_),
    .B1(\line_cache[13][6] ),
    .B2(_05839_),
    .C1(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__nand2_1 _21803_ (.A(_05353_),
    .B(\line_cache[10][6] ),
    .Y(_07177_));
 sky130_fd_sc_hd__nand2_1 _21804_ (.A(_05351_),
    .B(\line_cache[9][6] ),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_1 _21805_ (.A(_07177_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__a221oi_2 _21806_ (.A1(_05355_),
    .A2(\line_cache[8][6] ),
    .B1(_05346_),
    .B2(\line_cache[7][6] ),
    .C1(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__nand2_1 _21807_ (.A(_07176_),
    .B(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__and3_1 _21808_ (.A(_05163_),
    .B(_05812_),
    .C(\line_cache[21][6] ),
    .X(_07182_));
 sky130_fd_sc_hd__and3_1 _21809_ (.A(_05167_),
    .B(_05812_),
    .C(\line_cache[20][6] ),
    .X(_07183_));
 sky130_fd_sc_hd__a22o_1 _21810_ (.A1(_05825_),
    .A2(\line_cache[23][6] ),
    .B1(\line_cache[22][6] ),
    .B2(_05826_),
    .X(_07184_));
 sky130_fd_sc_hd__a22o_1 _21811_ (.A1(_05329_),
    .A2(\line_cache[16][6] ),
    .B1(\line_cache[17][6] ),
    .B2(_05330_),
    .X(_07185_));
 sky130_fd_sc_hd__a221o_1 _21812_ (.A1(\line_cache[19][6] ),
    .A2(_05831_),
    .B1(\line_cache[18][6] ),
    .B2(_05832_),
    .C1(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__or4_1 _21813_ (.A(_07182_),
    .B(_07183_),
    .C(_07184_),
    .D(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__a22o_1 _21814_ (.A1(_05262_),
    .A2(\line_cache[33][6] ),
    .B1(\line_cache[34][6] ),
    .B2(_05263_),
    .X(_07188_));
 sky130_fd_sc_hd__a221o_1 _21815_ (.A1(\line_cache[36][6] ),
    .A2(_05266_),
    .B1(\line_cache[35][6] ),
    .B2(_05261_),
    .C1(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__and3_1 _21816_ (.A(_05146_),
    .B(_05792_),
    .C(\line_cache[25][6] ),
    .X(_07190_));
 sky130_fd_sc_hd__a31o_1 _21817_ (.A1(_05840_),
    .A2(\line_cache[24][6] ),
    .A3(_05320_),
    .B1(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__a221oi_2 _21818_ (.A1(\line_cache[27][6] ),
    .A2(_05817_),
    .B1(\line_cache[26][6] ),
    .B2(_05819_),
    .C1(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__a32o_1 _21819_ (.A1(_05175_),
    .A2(_05812_),
    .A3(\line_cache[30][6] ),
    .B1(_05260_),
    .B2(\line_cache[32][6] ),
    .X(_07193_));
 sky130_fd_sc_hd__a32o_1 _21820_ (.A1(_05840_),
    .A2(_05173_),
    .A3(\line_cache[29][6] ),
    .B1(_06051_),
    .B2(\line_cache[28][6] ),
    .X(_07194_));
 sky130_fd_sc_hd__nor2_1 _21821_ (.A(_07193_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__nand2_1 _21822_ (.A(_05270_),
    .B(\line_cache[38][6] ),
    .Y(_07196_));
 sky130_fd_sc_hd__nand2_1 _21823_ (.A(_05272_),
    .B(\line_cache[37][6] ),
    .Y(_07197_));
 sky130_fd_sc_hd__nand2_1 _21824_ (.A(_07196_),
    .B(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__a221oi_2 _21825_ (.A1(_05268_),
    .A2(\line_cache[39][6] ),
    .B1(\line_cache[40][6] ),
    .B2(_05275_),
    .C1(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__and4b_1 _21826_ (.A_N(_07189_),
    .B(_07192_),
    .C(_07195_),
    .D(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__or3b_2 _21827_ (.A(_07181_),
    .B(_07187_),
    .C_N(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__nor3_2 _21828_ (.A(_07148_),
    .B(_07172_),
    .C(_07201_),
    .Y(_07202_));
 sky130_fd_sc_hd__and3_1 _21829_ (.A(_05058_),
    .B(_05176_),
    .C(\line_cache[302][6] ),
    .X(_07203_));
 sky130_fd_sc_hd__a22o_1 _21830_ (.A1(_05056_),
    .A2(\line_cache[301][6] ),
    .B1(\line_cache[300][6] ),
    .B2(_05053_),
    .X(_07204_));
 sky130_fd_sc_hd__a211o_1 _21831_ (.A1(\line_cache[256][6] ),
    .A2(_05777_),
    .B1(_07203_),
    .C1(_07204_),
    .X(_07205_));
 sky130_fd_sc_hd__and3_1 _21832_ (.A(_05779_),
    .B(_05021_),
    .C(\line_cache[258][6] ),
    .X(_07206_));
 sky130_fd_sc_hd__and3_1 _21833_ (.A(_05771_),
    .B(_05034_),
    .C(\line_cache[260][6] ),
    .X(_07207_));
 sky130_fd_sc_hd__and3_1 _21834_ (.A(_05778_),
    .B(_05176_),
    .C(\line_cache[259][6] ),
    .X(_07208_));
 sky130_fd_sc_hd__a2111o_1 _21835_ (.A1(\line_cache[257][6] ),
    .A2(_05776_),
    .B1(_07206_),
    .C1(_07207_),
    .D1(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__and3_1 _21836_ (.A(_05356_),
    .B(_05176_),
    .C(\line_cache[267][6] ),
    .X(_07210_));
 sky130_fd_sc_hd__a22o_1 _21837_ (.A1(_05760_),
    .A2(\line_cache[266][6] ),
    .B1(\line_cache[265][6] ),
    .B2(_05764_),
    .X(_07211_));
 sky130_fd_sc_hd__a311o_1 _21838_ (.A1(_05113_),
    .A2(\line_cache[268][6] ),
    .A3(_05364_),
    .B1(_07210_),
    .C1(_07211_),
    .X(_07212_));
 sky130_fd_sc_hd__nand2_1 _21839_ (.A(_05768_),
    .B(\line_cache[262][6] ),
    .Y(_07213_));
 sky130_fd_sc_hd__nand2_1 _21840_ (.A(_05773_),
    .B(\line_cache[261][6] ),
    .Y(_07214_));
 sky130_fd_sc_hd__nand2_1 _21841_ (.A(_07213_),
    .B(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__a221oi_1 _21842_ (.A1(_05763_),
    .A2(\line_cache[264][6] ),
    .B1(_05770_),
    .B2(\line_cache[263][6] ),
    .C1(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__or4b_1 _21843_ (.A(_07205_),
    .B(_07209_),
    .C(_07212_),
    .D_N(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__a22o_1 _21844_ (.A1(_05098_),
    .A2(\line_cache[308][6] ),
    .B1(\line_cache[309][6] ),
    .B2(_05093_),
    .X(_07218_));
 sky130_fd_sc_hd__a221o_1 _21845_ (.A1(\line_cache[311][6] ),
    .A2(_05097_),
    .B1(\line_cache[310][6] ),
    .B2(_05103_),
    .C1(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__a22o_1 _21846_ (.A1(_05046_),
    .A2(\line_cache[295][6] ),
    .B1(\line_cache[294][6] ),
    .B2(_05043_),
    .X(_07220_));
 sky130_fd_sc_hd__a221o_1 _21847_ (.A1(\line_cache[293][6] ),
    .A2(_05628_),
    .B1(\line_cache[292][6] ),
    .B2(_05627_),
    .C1(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__a22o_1 _21848_ (.A1(_05069_),
    .A2(\line_cache[296][6] ),
    .B1(\line_cache[297][6] ),
    .B2(_05076_),
    .X(_07222_));
 sky130_fd_sc_hd__a221o_1 _21849_ (.A1(\line_cache[299][6] ),
    .A2(_05073_),
    .B1(\line_cache[298][6] ),
    .B2(_05079_),
    .C1(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__a22o_1 _21850_ (.A1(_05632_),
    .A2(\line_cache[288][6] ),
    .B1(\line_cache[289][6] ),
    .B2(_05633_),
    .X(_07224_));
 sky130_fd_sc_hd__a221o_1 _21851_ (.A1(\line_cache[291][6] ),
    .A2(_05623_),
    .B1(\line_cache[290][6] ),
    .B2(_05624_),
    .C1(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__or4_2 _21852_ (.A(_07219_),
    .B(_07221_),
    .C(_07223_),
    .D(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__nor2_1 _21853_ (.A(_07217_),
    .B(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__and3_1 _21854_ (.A(_05203_),
    .B(\line_cache[203][6] ),
    .C(_05471_),
    .X(_07228_));
 sky130_fd_sc_hd__and3_1 _21855_ (.A(_05586_),
    .B(\line_cache[206][6] ),
    .C(_05471_),
    .X(_07229_));
 sky130_fd_sc_hd__and2b_1 _21856_ (.A_N(_05687_),
    .B(\line_cache[204][6] ),
    .X(_07230_));
 sky130_fd_sc_hd__a2111o_1 _21857_ (.A1(\line_cache[205][6] ),
    .A2(_05683_),
    .B1(_07228_),
    .C1(_07229_),
    .D1(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__a22o_1 _21858_ (.A1(_05484_),
    .A2(\line_cache[195][6] ),
    .B1(_05485_),
    .B2(\line_cache[196][6] ),
    .X(_07232_));
 sky130_fd_sc_hd__a221o_1 _21859_ (.A1(\line_cache[198][6] ),
    .A2(_05487_),
    .B1(\line_cache[197][6] ),
    .B2(_05489_),
    .C1(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__a22o_1 _21860_ (.A1(_05495_),
    .A2(\line_cache[200][6] ),
    .B1(_05493_),
    .B2(\line_cache[199][6] ),
    .X(_07234_));
 sky130_fd_sc_hd__a221o_1 _21861_ (.A1(\line_cache[202][6] ),
    .A2(_05492_),
    .B1(\line_cache[201][6] ),
    .B2(_05491_),
    .C1(_07234_),
    .X(_07235_));
 sky130_fd_sc_hd__and3_1 _21862_ (.A(_05470_),
    .B(\line_cache[193][6] ),
    .C(_05685_),
    .X(_07236_));
 sky130_fd_sc_hd__and3_1 _21863_ (.A(_05475_),
    .B(\line_cache[192][6] ),
    .C(_05685_),
    .X(_07237_));
 sky130_fd_sc_hd__and3_1 _21864_ (.A(_05408_),
    .B(\line_cache[194][6] ),
    .C(_05472_),
    .X(_07238_));
 sky130_fd_sc_hd__a2111o_1 _21865_ (.A1(_05630_),
    .A2(\line_cache[286][6] ),
    .B1(_07236_),
    .C1(_07237_),
    .D1(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__or4_1 _21866_ (.A(_07231_),
    .B(_07233_),
    .C(_07235_),
    .D(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__a22o_1 _21867_ (.A1(_05659_),
    .A2(\line_cache[275][6] ),
    .B1(\line_cache[274][6] ),
    .B2(_05662_),
    .X(_07241_));
 sky130_fd_sc_hd__a22o_1 _21868_ (.A1(_05658_),
    .A2(\line_cache[276][6] ),
    .B1(\line_cache[277][6] ),
    .B2(_05655_),
    .X(_07242_));
 sky130_fd_sc_hd__a22o_1 _21869_ (.A1(_05668_),
    .A2(\line_cache[270][6] ),
    .B1(\line_cache[269][6] ),
    .B2(_05670_),
    .X(_07243_));
 sky130_fd_sc_hd__a221o_1 _21870_ (.A1(\line_cache[273][6] ),
    .A2(_05660_),
    .B1(\line_cache[272][6] ),
    .B2(_05666_),
    .C1(_07243_),
    .X(_07244_));
 sky130_fd_sc_hd__a22oi_1 _21871_ (.A1(_05676_),
    .A2(\line_cache[283][6] ),
    .B1(_05678_),
    .B2(\line_cache[282][6] ),
    .Y(_07245_));
 sky130_fd_sc_hd__a22oi_1 _21872_ (.A1(_05674_),
    .A2(\line_cache[284][6] ),
    .B1(_05631_),
    .B2(\line_cache[285][6] ),
    .Y(_07246_));
 sky130_fd_sc_hd__nand2_1 _21873_ (.A(_07245_),
    .B(_07246_),
    .Y(_07247_));
 sky130_fd_sc_hd__a22o_1 _21874_ (.A1(_05144_),
    .A2(\line_cache[280][6] ),
    .B1(_05677_),
    .B2(\line_cache[281][6] ),
    .X(_07248_));
 sky130_fd_sc_hd__a32o_1 _21875_ (.A1(_05165_),
    .A2(_05151_),
    .A3(\line_cache[278][6] ),
    .B1(_05654_),
    .B2(\line_cache[279][6] ),
    .X(_07249_));
 sky130_fd_sc_hd__nor3_1 _21876_ (.A(_07247_),
    .B(_07248_),
    .C(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__or4b_2 _21877_ (.A(_07241_),
    .B(_07242_),
    .C(_07244_),
    .D_N(_07250_),
    .X(_07251_));
 sky130_fd_sc_hd__nor2_1 _21878_ (.A(_07240_),
    .B(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__a22o_1 _21879_ (.A1(_05746_),
    .A2(\line_cache[236][6] ),
    .B1(_05747_),
    .B2(\line_cache[235][6] ),
    .X(_07253_));
 sky130_fd_sc_hd__a221o_1 _21880_ (.A1(\line_cache[238][6] ),
    .A2(_05744_),
    .B1(\line_cache[237][6] ),
    .B2(_05745_),
    .C1(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__and3_1 _21881_ (.A(_05469_),
    .B(\line_cache[225][6] ),
    .C(_05732_),
    .X(_07255_));
 sky130_fd_sc_hd__and3_1 _21882_ (.A(_05408_),
    .B(\line_cache[226][6] ),
    .C(_05721_),
    .X(_07256_));
 sky130_fd_sc_hd__and3_1 _21883_ (.A(_05475_),
    .B(\line_cache[224][6] ),
    .C(_05721_),
    .X(_07257_));
 sky130_fd_sc_hd__a2111o_1 _21884_ (.A1(\line_cache[223][6] ),
    .A2(_05720_),
    .B1(_07255_),
    .C1(_07256_),
    .D1(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__and3_1 _21885_ (.A(_05704_),
    .B(\line_cache[227][6] ),
    .C(_05193_),
    .X(_07259_));
 sky130_fd_sc_hd__and3_1 _21886_ (.A(_05610_),
    .B(\line_cache[228][6] ),
    .C(_05193_),
    .X(_07260_));
 sky130_fd_sc_hd__and3_1 _21887_ (.A(_05710_),
    .B(\line_cache[229][6] ),
    .C(_05193_),
    .X(_07261_));
 sky130_fd_sc_hd__and3_1 _21888_ (.A(_05708_),
    .B(\line_cache[230][6] ),
    .C(_05732_),
    .X(_07262_));
 sky130_fd_sc_hd__or4_1 _21889_ (.A(_07259_),
    .B(_07260_),
    .C(_07261_),
    .D(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__a22o_1 _21890_ (.A1(_05728_),
    .A2(\line_cache[232][6] ),
    .B1(_05729_),
    .B2(\line_cache[231][6] ),
    .X(_07264_));
 sky130_fd_sc_hd__a221o_1 _21891_ (.A1(\line_cache[234][6] ),
    .A2(_05726_),
    .B1(\line_cache[233][6] ),
    .B2(_05727_),
    .C1(_07264_),
    .X(_07265_));
 sky130_fd_sc_hd__or4_1 _21892_ (.A(_07254_),
    .B(_07258_),
    .C(_07263_),
    .D(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__a22o_1 _21893_ (.A1(_05716_),
    .A2(\line_cache[220][6] ),
    .B1(_05717_),
    .B2(\line_cache[219][6] ),
    .X(_07267_));
 sky130_fd_sc_hd__a221o_1 _21894_ (.A1(\line_cache[222][6] ),
    .A2(_05714_),
    .B1(\line_cache[221][6] ),
    .B2(_05715_),
    .C1(_07267_),
    .X(_07268_));
 sky130_fd_sc_hd__a22o_1 _21895_ (.A1(_05700_),
    .A2(\line_cache[209][6] ),
    .B1(\line_cache[210][6] ),
    .B2(_05701_),
    .X(_07269_));
 sky130_fd_sc_hd__a221o_1 _21896_ (.A1(\line_cache[208][6] ),
    .A2(_05698_),
    .B1(\line_cache[207][6] ),
    .B2(_05699_),
    .C1(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__and3_1 _21897_ (.A(_05704_),
    .B(\line_cache[211][6] ),
    .C(_05694_),
    .X(_07271_));
 sky130_fd_sc_hd__and3_1 _21898_ (.A(_05611_),
    .B(\line_cache[212][6] ),
    .C(_05694_),
    .X(_07272_));
 sky130_fd_sc_hd__and3_1 _21899_ (.A(_05710_),
    .B(\line_cache[213][6] ),
    .C(_05694_),
    .X(_07273_));
 sky130_fd_sc_hd__and3_1 _21900_ (.A(_05708_),
    .B(\line_cache[214][6] ),
    .C(_05706_),
    .X(_07274_));
 sky130_fd_sc_hd__or4_1 _21901_ (.A(_07271_),
    .B(_07272_),
    .C(_07273_),
    .D(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__a22o_1 _21902_ (.A1(_05692_),
    .A2(\line_cache[216][6] ),
    .B1(_05983_),
    .B2(\line_cache[215][6] ),
    .X(_07276_));
 sky130_fd_sc_hd__a221o_1 _21903_ (.A1(\line_cache[218][6] ),
    .A2(_05690_),
    .B1(\line_cache[217][6] ),
    .B2(_05691_),
    .C1(_07276_),
    .X(_07277_));
 sky130_fd_sc_hd__or4_2 _21904_ (.A(_07268_),
    .B(_07270_),
    .C(_07275_),
    .D(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__nor2_1 _21905_ (.A(_07266_),
    .B(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__and3_1 _21906_ (.A(_05454_),
    .B(\line_cache[239][6] ),
    .C(_05732_),
    .X(_07280_));
 sky130_fd_sc_hd__and3_1 _21907_ (.A(_05470_),
    .B(\line_cache[241][6] ),
    .C(_05206_),
    .X(_07281_));
 sky130_fd_sc_hd__and3_1 _21908_ (.A(_05408_),
    .B(\line_cache[242][6] ),
    .C(_05206_),
    .X(_07282_));
 sky130_fd_sc_hd__a2111o_1 _21909_ (.A1(_05233_),
    .A2(\line_cache[240][6] ),
    .B1(_07280_),
    .C1(_07281_),
    .D1(_07282_),
    .X(_07283_));
 sky130_fd_sc_hd__and2_1 _21910_ (.A(_05235_),
    .B(\line_cache[243][6] ),
    .X(_07284_));
 sky130_fd_sc_hd__a21o_1 _21911_ (.A1(\line_cache[244][6] ),
    .A2(_05224_),
    .B1(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__a221o_1 _21912_ (.A1(\line_cache[246][6] ),
    .A2(_05753_),
    .B1(\line_cache[245][6] ),
    .B2(_05226_),
    .C1(_07285_),
    .X(_07286_));
 sky130_fd_sc_hd__a22o_1 _21913_ (.A1(_05212_),
    .A2(\line_cache[252][6] ),
    .B1(_05205_),
    .B2(\line_cache[251][6] ),
    .X(_07287_));
 sky130_fd_sc_hd__a221o_1 _21914_ (.A1(\line_cache[254][6] ),
    .A2(_05217_),
    .B1(\line_cache[253][6] ),
    .B2(_05214_),
    .C1(_07287_),
    .X(_07288_));
 sky130_fd_sc_hd__a22o_1 _21915_ (.A1(_05750_),
    .A2(\line_cache[248][6] ),
    .B1(_05229_),
    .B2(\line_cache[247][6] ),
    .X(_07289_));
 sky130_fd_sc_hd__a221o_1 _21916_ (.A1(\line_cache[250][6] ),
    .A2(_05202_),
    .B1(\line_cache[249][6] ),
    .B2(_05209_),
    .C1(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__or4_1 _21917_ (.A(_07283_),
    .B(_07286_),
    .C(_07288_),
    .D(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__a22o_1 _21918_ (.A1(_05875_),
    .A2(\line_cache[67][6] ),
    .B1(_05861_),
    .B2(\line_cache[66][6] ),
    .X(_07292_));
 sky130_fd_sc_hd__a221o_1 _21919_ (.A1(\line_cache[65][6] ),
    .A2(_05860_),
    .B1(\line_cache[64][6] ),
    .B2(_05858_),
    .C1(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__a22o_1 _21920_ (.A1(_05867_),
    .A2(\line_cache[72][6] ),
    .B1(_05866_),
    .B2(\line_cache[73][6] ),
    .X(_07294_));
 sky130_fd_sc_hd__a221o_1 _21921_ (.A1(\line_cache[75][6] ),
    .A2(_05543_),
    .B1(\line_cache[74][6] ),
    .B2(_05865_),
    .C1(_07294_),
    .X(_07295_));
 sky130_fd_sc_hd__a22o_1 _21922_ (.A1(_05873_),
    .A2(\line_cache[68][6] ),
    .B1(_05872_),
    .B2(\line_cache[69][6] ),
    .X(_07296_));
 sky130_fd_sc_hd__a221o_1 _21923_ (.A1(\line_cache[71][6] ),
    .A2(_05868_),
    .B1(\line_cache[70][6] ),
    .B2(_05871_),
    .C1(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__and2_1 _21924_ (.A(_05542_),
    .B(\line_cache[76][6] ),
    .X(_07298_));
 sky130_fd_sc_hd__and3_1 _21925_ (.A(_05544_),
    .B(\line_cache[77][6] ),
    .C(_05536_),
    .X(_07299_));
 sky130_fd_sc_hd__or2_1 _21926_ (.A(_07298_),
    .B(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__a221o_1 _21927_ (.A1(\line_cache[79][6] ),
    .A2(_05537_),
    .B1(\line_cache[78][6] ),
    .B2(_05545_),
    .C1(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__or4_4 _21928_ (.A(_07293_),
    .B(_07295_),
    .C(_07297_),
    .D(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__nor2_1 _21929_ (.A(_07291_),
    .B(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__and4_1 _21930_ (.A(_07227_),
    .B(_07252_),
    .C(_07279_),
    .D(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__and3_1 _21931_ (.A(_05207_),
    .B(\line_cache[89][6] ),
    .C(_05518_),
    .X(_07305_));
 sky130_fd_sc_hd__a21o_1 _21932_ (.A1(\line_cache[88][6] ),
    .A2(_05553_),
    .B1(_07305_),
    .X(_07306_));
 sky130_fd_sc_hd__a221o_1 _21933_ (.A1(\line_cache[91][6] ),
    .A2(_05525_),
    .B1(\line_cache[90][6] ),
    .B2(_05550_),
    .C1(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__a22o_1 _21934_ (.A1(_05531_),
    .A2(\line_cache[83][6] ),
    .B1(_05539_),
    .B2(\line_cache[82][6] ),
    .X(_07308_));
 sky130_fd_sc_hd__a221o_1 _21935_ (.A1(\line_cache[81][6] ),
    .A2(_05538_),
    .B1(\line_cache[80][6] ),
    .B2(_05535_),
    .C1(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__a22o_1 _21936_ (.A1(_05532_),
    .A2(\line_cache[84][6] ),
    .B1(\line_cache[85][6] ),
    .B2(_05530_),
    .X(_07310_));
 sky130_fd_sc_hd__a221o_1 _21937_ (.A1(\line_cache[87][6] ),
    .A2(_05551_),
    .B1(\line_cache[86][6] ),
    .B2(_05529_),
    .C1(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__a22o_1 _21938_ (.A1(_05524_),
    .A2(\line_cache[92][6] ),
    .B1(_05523_),
    .B2(\line_cache[93][6] ),
    .X(_07312_));
 sky130_fd_sc_hd__a221o_1 _21939_ (.A1(\line_cache[95][6] ),
    .A2(_05519_),
    .B1(\line_cache[94][6] ),
    .B2(_05522_),
    .C1(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__or4_1 _21940_ (.A(_07307_),
    .B(_07309_),
    .C(_07311_),
    .D(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__a22o_1 _21941_ (.A1(_05510_),
    .A2(\line_cache[99][6] ),
    .B1(_05516_),
    .B2(\line_cache[98][6] ),
    .X(_07315_));
 sky130_fd_sc_hd__a221o_1 _21942_ (.A1(\line_cache[97][6] ),
    .A2(_05515_),
    .B1(\line_cache[96][6] ),
    .B2(_05520_),
    .C1(_07315_),
    .X(_07316_));
 sky130_fd_sc_hd__a22o_1 _21943_ (.A1(_05575_),
    .A2(\line_cache[108][6] ),
    .B1(_05574_),
    .B2(\line_cache[109][6] ),
    .X(_07317_));
 sky130_fd_sc_hd__a221o_1 _21944_ (.A1(\line_cache[111][6] ),
    .A2(_05580_),
    .B1(\line_cache[110][6] ),
    .B2(_05573_),
    .C1(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__a22o_1 _21945_ (.A1(_05511_),
    .A2(\line_cache[100][6] ),
    .B1(\line_cache[101][6] ),
    .B2(_05509_),
    .X(_07319_));
 sky130_fd_sc_hd__a221o_1 _21946_ (.A1(\line_cache[103][6] ),
    .A2(_05504_),
    .B1(\line_cache[102][6] ),
    .B2(_05502_),
    .C1(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__a22o_1 _21947_ (.A1(_05503_),
    .A2(\line_cache[104][6] ),
    .B1(_05508_),
    .B2(\line_cache[105][6] ),
    .X(_07321_));
 sky130_fd_sc_hd__a221o_1 _21948_ (.A1(\line_cache[107][6] ),
    .A2(_05576_),
    .B1(\line_cache[106][6] ),
    .B2(_05506_),
    .C1(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__or4_1 _21949_ (.A(_07316_),
    .B(_07318_),
    .C(_07320_),
    .D(_07322_),
    .X(_07323_));
 sky130_fd_sc_hd__nor2_1 _21950_ (.A(_07314_),
    .B(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__and3_1 _21951_ (.A(_05586_),
    .B(\line_cache[126][6] ),
    .C(_05562_),
    .X(_07325_));
 sky130_fd_sc_hd__a21o_1 _21952_ (.A1(\line_cache[127][6] ),
    .A2(_05596_),
    .B1(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__a221o_1 _21953_ (.A1(\line_cache[125][6] ),
    .A2(_05589_),
    .B1(\line_cache[124][6] ),
    .B2(_05590_),
    .C1(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__a22o_1 _21954_ (.A1(_05569_),
    .A2(\line_cache[115][6] ),
    .B1(_05582_),
    .B2(\line_cache[114][6] ),
    .X(_07328_));
 sky130_fd_sc_hd__a221o_1 _21955_ (.A1(\line_cache[113][6] ),
    .A2(_05581_),
    .B1(\line_cache[112][6] ),
    .B2(_05579_),
    .C1(_07328_),
    .X(_07329_));
 sky130_fd_sc_hd__a22o_1 _21956_ (.A1(_05591_),
    .A2(\line_cache[123][6] ),
    .B1(\line_cache[122][6] ),
    .B2(_05559_),
    .X(_07330_));
 sky130_fd_sc_hd__a221o_1 _21957_ (.A1(\line_cache[121][6] ),
    .A2(_05560_),
    .B1(\line_cache[120][6] ),
    .B2(_05561_),
    .C1(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__a22o_1 _21958_ (.A1(_05568_),
    .A2(\line_cache[116][6] ),
    .B1(_05567_),
    .B2(\line_cache[117][6] ),
    .X(_07332_));
 sky130_fd_sc_hd__a221o_1 _21959_ (.A1(\line_cache[119][6] ),
    .A2(_06088_),
    .B1(\line_cache[118][6] ),
    .B2(_05566_),
    .C1(_07332_),
    .X(_07333_));
 sky130_fd_sc_hd__or4_1 _21960_ (.A(_07327_),
    .B(_07329_),
    .C(_07331_),
    .D(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__a22o_1 _21961_ (.A1(_05376_),
    .A2(\line_cache[140][6] ),
    .B1(_05375_),
    .B2(\line_cache[141][6] ),
    .X(_07335_));
 sky130_fd_sc_hd__a221o_1 _21962_ (.A1(\line_cache[143][6] ),
    .A2(_05382_),
    .B1(\line_cache[142][6] ),
    .B2(_05374_),
    .C1(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__a22o_1 _21963_ (.A1(_05604_),
    .A2(\line_cache[136][6] ),
    .B1(_05603_),
    .B2(\line_cache[137][6] ),
    .X(_07337_));
 sky130_fd_sc_hd__a221o_1 _21964_ (.A1(\line_cache[139][6] ),
    .A2(_05377_),
    .B1(\line_cache[138][6] ),
    .B2(_05602_),
    .C1(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__and2_1 _21965_ (.A(_05597_),
    .B(\line_cache[129][6] ),
    .X(_07339_));
 sky130_fd_sc_hd__a21o_1 _21966_ (.A1(_05594_),
    .A2(\line_cache[128][6] ),
    .B1(_07339_),
    .X(_07340_));
 sky130_fd_sc_hd__a221o_1 _21967_ (.A1(\line_cache[131][6] ),
    .A2(_05612_),
    .B1(\line_cache[130][6] ),
    .B2(_05598_),
    .C1(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__and2_1 _21968_ (.A(_05609_),
    .B(\line_cache[133][6] ),
    .X(_07342_));
 sky130_fd_sc_hd__and3_1 _21969_ (.A(_05611_),
    .B(\line_cache[132][6] ),
    .C(_05381_),
    .X(_07343_));
 sky130_fd_sc_hd__or2_1 _21970_ (.A(_07342_),
    .B(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__a221o_1 _21971_ (.A1(\line_cache[135][6] ),
    .A2(_05605_),
    .B1(\line_cache[134][6] ),
    .B2(_05608_),
    .C1(_07344_),
    .X(_07345_));
 sky130_fd_sc_hd__or4_1 _21972_ (.A(_07336_),
    .B(_07338_),
    .C(_07341_),
    .D(_07345_),
    .X(_07346_));
 sky130_fd_sc_hd__nor2_1 _21973_ (.A(_07334_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__a22o_1 _21974_ (.A1(_05464_),
    .A2(\line_cache[171][6] ),
    .B1(\line_cache[170][6] ),
    .B2(_05424_),
    .X(_07348_));
 sky130_fd_sc_hd__a221o_1 _21975_ (.A1(\line_cache[169][6] ),
    .A2(_05423_),
    .B1(\line_cache[168][6] ),
    .B2(_05427_),
    .C1(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__a32o_1 _21976_ (.A1(_05409_),
    .A2(\line_cache[162][6] ),
    .A3(_05410_),
    .B1(\line_cache[163][6] ),
    .B2(_05433_),
    .X(_07350_));
 sky130_fd_sc_hd__a221oi_1 _21977_ (.A1(\line_cache[161][6] ),
    .A2(_05406_),
    .B1(\line_cache[160][6] ),
    .B2(_05414_),
    .C1(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__a22o_1 _21978_ (.A1(_05434_),
    .A2(\line_cache[164][6] ),
    .B1(\line_cache[165][6] ),
    .B2(_05432_),
    .X(_07352_));
 sky130_fd_sc_hd__a221oi_2 _21979_ (.A1(\line_cache[167][6] ),
    .A2(_05425_),
    .B1(\line_cache[166][6] ),
    .B2(_05431_),
    .C1(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__a22o_1 _21980_ (.A1(_05463_),
    .A2(\line_cache[172][6] ),
    .B1(_05462_),
    .B2(\line_cache[173][6] ),
    .X(_07354_));
 sky130_fd_sc_hd__a221oi_1 _21981_ (.A1(\line_cache[175][6] ),
    .A2(_05456_),
    .B1(\line_cache[174][6] ),
    .B2(_05461_),
    .C1(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__and4b_1 _21982_ (.A_N(_07349_),
    .B(_07351_),
    .C(_07353_),
    .D(_07355_),
    .X(_07356_));
 sky130_fd_sc_hd__a22o_1 _21983_ (.A1(_05438_),
    .A2(\line_cache[184][6] ),
    .B1(_05440_),
    .B2(\line_cache[185][6] ),
    .X(_07357_));
 sky130_fd_sc_hd__a221o_1 _21984_ (.A1(\line_cache[187][6] ),
    .A2(_05481_),
    .B1(\line_cache[186][6] ),
    .B2(_06131_),
    .C1(_07357_),
    .X(_07358_));
 sky130_fd_sc_hd__a22o_1 _21985_ (.A1(_05449_),
    .A2(\line_cache[180][6] ),
    .B1(_05446_),
    .B2(\line_cache[181][6] ),
    .X(_07359_));
 sky130_fd_sc_hd__a221oi_2 _21986_ (.A1(\line_cache[183][6] ),
    .A2(_05439_),
    .B1(\line_cache[182][6] ),
    .B2(_05445_),
    .C1(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__a22o_1 _21987_ (.A1(_05447_),
    .A2(\line_cache[179][6] ),
    .B1(\line_cache[178][6] ),
    .B2(_05458_),
    .X(_07361_));
 sky130_fd_sc_hd__a221oi_1 _21988_ (.A1(\line_cache[177][6] ),
    .A2(_05457_),
    .B1(\line_cache[176][6] ),
    .B2(_05453_),
    .C1(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__a22o_1 _21989_ (.A1(_05480_),
    .A2(\line_cache[188][6] ),
    .B1(_05479_),
    .B2(\line_cache[189][6] ),
    .X(_07363_));
 sky130_fd_sc_hd__a221oi_2 _21990_ (.A1(\line_cache[191][6] ),
    .A2(_05468_),
    .B1(\line_cache[190][6] ),
    .B2(_05478_),
    .C1(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__and4b_1 _21991_ (.A_N(_07358_),
    .B(_07360_),
    .C(_07362_),
    .D(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__a22o_1 _21992_ (.A1(_05393_),
    .A2(\line_cache[148][6] ),
    .B1(\line_cache[149][6] ),
    .B2(_05391_),
    .X(_07366_));
 sky130_fd_sc_hd__a221oi_1 _21993_ (.A1(\line_cache[151][6] ),
    .A2(_05398_),
    .B1(\line_cache[150][6] ),
    .B2(_05390_),
    .C1(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__nand2_1 _21994_ (.A(_05386_),
    .B(\line_cache[146][6] ),
    .Y(_07368_));
 sky130_fd_sc_hd__nand2_1 _21995_ (.A(_05392_),
    .B(\line_cache[147][6] ),
    .Y(_07369_));
 sky130_fd_sc_hd__nand2_1 _21996_ (.A(_07368_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__a221oi_2 _21997_ (.A1(\line_cache[145][6] ),
    .A2(_05384_),
    .B1(_05380_),
    .B2(\line_cache[144][6] ),
    .C1(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__nand2_1 _21998_ (.A(_07367_),
    .B(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__a22o_1 _21999_ (.A1(_05418_),
    .A2(\line_cache[156][6] ),
    .B1(_05417_),
    .B2(\line_cache[157][6] ),
    .X(_07373_));
 sky130_fd_sc_hd__a221o_1 _22000_ (.A1(\line_cache[159][6] ),
    .A2(_05413_),
    .B1(\line_cache[158][6] ),
    .B2(_05416_),
    .C1(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__a22o_1 _22001_ (.A1(_05419_),
    .A2(\line_cache[155][6] ),
    .B1(\line_cache[154][6] ),
    .B2(_06107_),
    .X(_07375_));
 sky130_fd_sc_hd__a221o_1 _22002_ (.A1(\line_cache[153][6] ),
    .A2(_05399_),
    .B1(\line_cache[152][6] ),
    .B2(_05397_),
    .C1(_07375_),
    .X(_07376_));
 sky130_fd_sc_hd__nor3_1 _22003_ (.A(_07372_),
    .B(_07374_),
    .C(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__and3_1 _22004_ (.A(_07356_),
    .B(_07365_),
    .C(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__and3_1 _22005_ (.A(_07324_),
    .B(_07347_),
    .C(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__nand3_1 _22006_ (.A(_07202_),
    .B(_07304_),
    .C(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__o21a_4 _22007_ (.A1(_07134_),
    .A2(_07380_),
    .B1(_05884_),
    .X(net132));
 sky130_fd_sc_hd__nor3b_1 _22008_ (.A(_05258_),
    .B(_05372_),
    .C_N(\line_cache[0][7] ),
    .Y(_07381_));
 sky130_fd_sc_hd__a22o_1 _22009_ (.A1(_05531_),
    .A2(\line_cache[83][7] ),
    .B1(_05539_),
    .B2(\line_cache[82][7] ),
    .X(_07382_));
 sky130_fd_sc_hd__a221o_1 _22010_ (.A1(\line_cache[81][7] ),
    .A2(_05538_),
    .B1(\line_cache[80][7] ),
    .B2(_05535_),
    .C1(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__a22o_1 _22011_ (.A1(_05524_),
    .A2(\line_cache[92][7] ),
    .B1(_05523_),
    .B2(\line_cache[93][7] ),
    .X(_07384_));
 sky130_fd_sc_hd__a221o_1 _22012_ (.A1(\line_cache[95][7] ),
    .A2(_05519_),
    .B1(\line_cache[94][7] ),
    .B2(_05522_),
    .C1(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__a22o_1 _22013_ (.A1(_05532_),
    .A2(\line_cache[84][7] ),
    .B1(\line_cache[85][7] ),
    .B2(_05530_),
    .X(_07386_));
 sky130_fd_sc_hd__a221o_1 _22014_ (.A1(\line_cache[87][7] ),
    .A2(_05551_),
    .B1(\line_cache[86][7] ),
    .B2(_05529_),
    .C1(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__a22o_1 _22015_ (.A1(_05553_),
    .A2(\line_cache[88][7] ),
    .B1(_05549_),
    .B2(\line_cache[89][7] ),
    .X(_07388_));
 sky130_fd_sc_hd__a221o_1 _22016_ (.A1(\line_cache[91][7] ),
    .A2(_05525_),
    .B1(\line_cache[90][7] ),
    .B2(_05550_),
    .C1(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__or4_2 _22017_ (.A(_07383_),
    .B(_07385_),
    .C(_07387_),
    .D(_07389_),
    .X(_07390_));
 sky130_fd_sc_hd__a22o_1 _22018_ (.A1(_05510_),
    .A2(\line_cache[99][7] ),
    .B1(_05516_),
    .B2(\line_cache[98][7] ),
    .X(_07391_));
 sky130_fd_sc_hd__a221o_1 _22019_ (.A1(\line_cache[97][7] ),
    .A2(_05515_),
    .B1(\line_cache[96][7] ),
    .B2(_05520_),
    .C1(_07391_),
    .X(_07392_));
 sky130_fd_sc_hd__a22o_1 _22020_ (.A1(_05575_),
    .A2(\line_cache[108][7] ),
    .B1(_05574_),
    .B2(\line_cache[109][7] ),
    .X(_07393_));
 sky130_fd_sc_hd__a221o_1 _22021_ (.A1(\line_cache[111][7] ),
    .A2(_05580_),
    .B1(\line_cache[110][7] ),
    .B2(_05573_),
    .C1(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__a22o_1 _22022_ (.A1(_05511_),
    .A2(\line_cache[100][7] ),
    .B1(\line_cache[101][7] ),
    .B2(_05509_),
    .X(_07395_));
 sky130_fd_sc_hd__a221o_1 _22023_ (.A1(\line_cache[103][7] ),
    .A2(_05504_),
    .B1(\line_cache[102][7] ),
    .B2(_05502_),
    .C1(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__a22o_1 _22024_ (.A1(_05503_),
    .A2(\line_cache[104][7] ),
    .B1(_05508_),
    .B2(\line_cache[105][7] ),
    .X(_07397_));
 sky130_fd_sc_hd__a221o_1 _22025_ (.A1(\line_cache[107][7] ),
    .A2(_05576_),
    .B1(\line_cache[106][7] ),
    .B2(_05506_),
    .C1(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__or4_1 _22026_ (.A(_07392_),
    .B(_07394_),
    .C(_07396_),
    .D(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__and2_1 _22027_ (.A(_05589_),
    .B(\line_cache[125][7] ),
    .X(_07400_));
 sky130_fd_sc_hd__and3_1 _22028_ (.A(_05586_),
    .B(\line_cache[126][7] ),
    .C(_05562_),
    .X(_07401_));
 sky130_fd_sc_hd__a21o_1 _22029_ (.A1(\line_cache[127][7] ),
    .A2(_05596_),
    .B1(_07401_),
    .X(_07402_));
 sky130_fd_sc_hd__a211o_1 _22030_ (.A1(\line_cache[124][7] ),
    .A2(_05590_),
    .B1(_07400_),
    .C1(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__and3_1 _22031_ (.A(_05207_),
    .B(\line_cache[121][7] ),
    .C(_05562_),
    .X(_07404_));
 sky130_fd_sc_hd__a21o_1 _22032_ (.A1(\line_cache[120][7] ),
    .A2(_05561_),
    .B1(_07404_),
    .X(_07405_));
 sky130_fd_sc_hd__a221o_1 _22033_ (.A1(\line_cache[123][7] ),
    .A2(_05591_),
    .B1(\line_cache[122][7] ),
    .B2(_05559_),
    .C1(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__a22o_1 _22034_ (.A1(_05569_),
    .A2(\line_cache[115][7] ),
    .B1(_05582_),
    .B2(\line_cache[114][7] ),
    .X(_07407_));
 sky130_fd_sc_hd__a221o_1 _22035_ (.A1(\line_cache[113][7] ),
    .A2(_05581_),
    .B1(\line_cache[112][7] ),
    .B2(_05579_),
    .C1(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__a22o_1 _22036_ (.A1(_05568_),
    .A2(\line_cache[116][7] ),
    .B1(_05567_),
    .B2(\line_cache[117][7] ),
    .X(_07409_));
 sky130_fd_sc_hd__a221o_1 _22037_ (.A1(\line_cache[119][7] ),
    .A2(_06088_),
    .B1(\line_cache[118][7] ),
    .B2(_05566_),
    .C1(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__or4_1 _22038_ (.A(_07403_),
    .B(_07406_),
    .C(_07408_),
    .D(_07410_),
    .X(_07411_));
 sky130_fd_sc_hd__and3_1 _22039_ (.A(_05207_),
    .B(\line_cache[137][7] ),
    .C(_05381_),
    .X(_07412_));
 sky130_fd_sc_hd__a21o_1 _22040_ (.A1(\line_cache[136][7] ),
    .A2(_05604_),
    .B1(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__a221o_1 _22041_ (.A1(\line_cache[139][7] ),
    .A2(_05377_),
    .B1(\line_cache[138][7] ),
    .B2(_05602_),
    .C1(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__a22o_1 _22042_ (.A1(_05376_),
    .A2(\line_cache[140][7] ),
    .B1(_05375_),
    .B2(\line_cache[141][7] ),
    .X(_07415_));
 sky130_fd_sc_hd__a221o_1 _22043_ (.A1(\line_cache[143][7] ),
    .A2(_05382_),
    .B1(\line_cache[142][7] ),
    .B2(_05374_),
    .C1(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__and2_1 _22044_ (.A(_05597_),
    .B(\line_cache[129][7] ),
    .X(_07417_));
 sky130_fd_sc_hd__a21o_1 _22045_ (.A1(_05594_),
    .A2(\line_cache[128][7] ),
    .B1(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__a221o_1 _22046_ (.A1(\line_cache[131][7] ),
    .A2(_05612_),
    .B1(\line_cache[130][7] ),
    .B2(_05598_),
    .C1(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__and2_1 _22047_ (.A(_05609_),
    .B(\line_cache[133][7] ),
    .X(_07420_));
 sky130_fd_sc_hd__and3_1 _22048_ (.A(_05610_),
    .B(\line_cache[132][7] ),
    .C(_05381_),
    .X(_07421_));
 sky130_fd_sc_hd__or2_1 _22049_ (.A(_07420_),
    .B(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__a221o_1 _22050_ (.A1(\line_cache[135][7] ),
    .A2(_05605_),
    .B1(\line_cache[134][7] ),
    .B2(_05608_),
    .C1(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__or4_1 _22051_ (.A(_07414_),
    .B(_07416_),
    .C(_07419_),
    .D(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__or2_1 _22052_ (.A(_07411_),
    .B(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__nor3_2 _22053_ (.A(_07390_),
    .B(_07399_),
    .C(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__a22o_1 _22054_ (.A1(_05449_),
    .A2(\line_cache[180][7] ),
    .B1(_05446_),
    .B2(\line_cache[181][7] ),
    .X(_07427_));
 sky130_fd_sc_hd__a221o_1 _22055_ (.A1(\line_cache[183][7] ),
    .A2(_05439_),
    .B1(\line_cache[182][7] ),
    .B2(_05445_),
    .C1(_07427_),
    .X(_07428_));
 sky130_fd_sc_hd__a22o_1 _22056_ (.A1(\line_cache[177][7] ),
    .A2(_05457_),
    .B1(_05453_),
    .B2(\line_cache[176][7] ),
    .X(_07429_));
 sky130_fd_sc_hd__a221o_1 _22057_ (.A1(\line_cache[179][7] ),
    .A2(_05447_),
    .B1(\line_cache[178][7] ),
    .B2(_05458_),
    .C1(_07429_),
    .X(_07430_));
 sky130_fd_sc_hd__and2_1 _22058_ (.A(_05479_),
    .B(\line_cache[189][7] ),
    .X(_07431_));
 sky130_fd_sc_hd__a22o_1 _22059_ (.A1(_05478_),
    .A2(\line_cache[190][7] ),
    .B1(_05468_),
    .B2(\line_cache[191][7] ),
    .X(_07432_));
 sky130_fd_sc_hd__a22o_1 _22060_ (.A1(_05438_),
    .A2(\line_cache[184][7] ),
    .B1(_05440_),
    .B2(\line_cache[185][7] ),
    .X(_07433_));
 sky130_fd_sc_hd__a221o_1 _22061_ (.A1(\line_cache[187][7] ),
    .A2(_05481_),
    .B1(\line_cache[186][7] ),
    .B2(_06131_),
    .C1(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__a2111o_1 _22062_ (.A1(\line_cache[188][7] ),
    .A2(_05480_),
    .B1(_07431_),
    .C1(_07432_),
    .D1(_07434_),
    .X(_07435_));
 sky130_fd_sc_hd__nor3_1 _22063_ (.A(_07428_),
    .B(_07430_),
    .C(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__a22o_1 _22064_ (.A1(_05419_),
    .A2(\line_cache[155][7] ),
    .B1(\line_cache[154][7] ),
    .B2(_06107_),
    .X(_07437_));
 sky130_fd_sc_hd__a221o_1 _22065_ (.A1(\line_cache[153][7] ),
    .A2(_05399_),
    .B1(\line_cache[152][7] ),
    .B2(_05397_),
    .C1(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__a22o_1 _22066_ (.A1(_05392_),
    .A2(\line_cache[147][7] ),
    .B1(_05386_),
    .B2(\line_cache[146][7] ),
    .X(_07439_));
 sky130_fd_sc_hd__a221oi_2 _22067_ (.A1(\line_cache[145][7] ),
    .A2(_05384_),
    .B1(\line_cache[144][7] ),
    .B2(_05380_),
    .C1(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__a22o_1 _22068_ (.A1(_05393_),
    .A2(\line_cache[148][7] ),
    .B1(\line_cache[149][7] ),
    .B2(_05391_),
    .X(_07441_));
 sky130_fd_sc_hd__a221oi_2 _22069_ (.A1(\line_cache[151][7] ),
    .A2(_05398_),
    .B1(\line_cache[150][7] ),
    .B2(_05390_),
    .C1(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__a22o_1 _22070_ (.A1(_05418_),
    .A2(\line_cache[156][7] ),
    .B1(_05417_),
    .B2(\line_cache[157][7] ),
    .X(_07443_));
 sky130_fd_sc_hd__a221oi_1 _22071_ (.A1(\line_cache[159][7] ),
    .A2(_05413_),
    .B1(\line_cache[158][7] ),
    .B2(_05416_),
    .C1(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__and4b_1 _22072_ (.A_N(_07438_),
    .B(_07440_),
    .C(_07442_),
    .D(_07444_),
    .X(_07445_));
 sky130_fd_sc_hd__a22o_1 _22073_ (.A1(_05464_),
    .A2(\line_cache[171][7] ),
    .B1(\line_cache[170][7] ),
    .B2(_05424_),
    .X(_07446_));
 sky130_fd_sc_hd__a221o_1 _22074_ (.A1(\line_cache[169][7] ),
    .A2(_05423_),
    .B1(\line_cache[168][7] ),
    .B2(_05427_),
    .C1(_07446_),
    .X(_07447_));
 sky130_fd_sc_hd__a32o_1 _22075_ (.A1(_05409_),
    .A2(\line_cache[162][7] ),
    .A3(_05410_),
    .B1(\line_cache[163][7] ),
    .B2(_05433_),
    .X(_07448_));
 sky130_fd_sc_hd__a221oi_2 _22076_ (.A1(\line_cache[161][7] ),
    .A2(_05406_),
    .B1(\line_cache[160][7] ),
    .B2(_05414_),
    .C1(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__a22o_1 _22077_ (.A1(_05434_),
    .A2(\line_cache[164][7] ),
    .B1(\line_cache[165][7] ),
    .B2(_05432_),
    .X(_07450_));
 sky130_fd_sc_hd__nand2_1 _22078_ (.A(_05431_),
    .B(\line_cache[166][7] ),
    .Y(_07451_));
 sky130_fd_sc_hd__nand2_1 _22079_ (.A(_05425_),
    .B(\line_cache[167][7] ),
    .Y(_07452_));
 sky130_fd_sc_hd__and3b_1 _22080_ (.A_N(_07450_),
    .B(_07451_),
    .C(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__nand2_1 _22081_ (.A(_05462_),
    .B(\line_cache[173][7] ),
    .Y(_07454_));
 sky130_fd_sc_hd__nand2_1 _22082_ (.A(_05463_),
    .B(\line_cache[172][7] ),
    .Y(_07455_));
 sky130_fd_sc_hd__nand2_1 _22083_ (.A(_07454_),
    .B(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__a221oi_1 _22084_ (.A1(_05461_),
    .A2(\line_cache[174][7] ),
    .B1(_05456_),
    .B2(\line_cache[175][7] ),
    .C1(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__and4b_1 _22085_ (.A_N(_07447_),
    .B(_07449_),
    .C(_07453_),
    .D(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__and4_2 _22086_ (.A(_07426_),
    .B(_07436_),
    .C(_07445_),
    .D(_07458_),
    .X(_07459_));
 sky130_fd_sc_hd__and2_1 _22087_ (.A(_05797_),
    .B(\line_cache[1][7] ),
    .X(_07460_));
 sky130_fd_sc_hd__and3_1 _22088_ (.A(_05779_),
    .B(_05991_),
    .C(\line_cache[2][7] ),
    .X(_07461_));
 sky130_fd_sc_hd__a211o_1 _22089_ (.A1(\line_cache[15][7] ),
    .A2(_05798_),
    .B1(_07460_),
    .C1(_07461_),
    .X(_07462_));
 sky130_fd_sc_hd__and3_1 _22090_ (.A(_05778_),
    .B(_05792_),
    .C(\line_cache[3][7] ),
    .X(_07463_));
 sky130_fd_sc_hd__a31o_1 _22091_ (.A1(_05840_),
    .A2(\line_cache[4][7] ),
    .A3(_05771_),
    .B1(_07463_),
    .X(_07464_));
 sky130_fd_sc_hd__a221o_1 _22092_ (.A1(_05343_),
    .A2(\line_cache[5][7] ),
    .B1(\line_cache[6][7] ),
    .B2(_05348_),
    .C1(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__and3_1 _22093_ (.A(_05112_),
    .B(_05151_),
    .C(\line_cache[319][7] ),
    .X(_07466_));
 sky130_fd_sc_hd__a32o_1 _22094_ (.A1(_05991_),
    .A2(_05180_),
    .A3(\line_cache[31][7] ),
    .B1(_05998_),
    .B2(\line_cache[47][7] ),
    .X(_07467_));
 sky130_fd_sc_hd__a311o_1 _22095_ (.A1(_05188_),
    .A2(\line_cache[63][7] ),
    .A3(_05112_),
    .B1(_07466_),
    .C1(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__nand2_1 _22096_ (.A(_05787_),
    .B(\line_cache[303][7] ),
    .Y(_07469_));
 sky130_fd_sc_hd__nand2_1 _22097_ (.A(_05791_),
    .B(\line_cache[271][7] ),
    .Y(_07470_));
 sky130_fd_sc_hd__nand2_1 _22098_ (.A(_07469_),
    .B(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__a221oi_4 _22099_ (.A1(\line_cache[255][7] ),
    .A2(_05220_),
    .B1(\line_cache[287][7] ),
    .B2(_05788_),
    .C1(_07471_),
    .Y(_07472_));
 sky130_fd_sc_hd__or4b_1 _22100_ (.A(_07462_),
    .B(_07465_),
    .C(_07468_),
    .D_N(_07472_),
    .X(_07473_));
 sky130_fd_sc_hd__a22o_1 _22101_ (.A1(_05283_),
    .A2(\line_cache[45][7] ),
    .B1(\line_cache[46][7] ),
    .B2(_05285_),
    .X(_07474_));
 sky130_fd_sc_hd__a22o_1 _22102_ (.A1(_05298_),
    .A2(\line_cache[48][7] ),
    .B1(\line_cache[49][7] ),
    .B2(_05300_),
    .X(_07475_));
 sky130_fd_sc_hd__nand2_1 _22103_ (.A(_05279_),
    .B(\line_cache[41][7] ),
    .Y(_07476_));
 sky130_fd_sc_hd__nand2_1 _22104_ (.A(_05281_),
    .B(\line_cache[42][7] ),
    .Y(_07477_));
 sky130_fd_sc_hd__nand2_1 _22105_ (.A(_07476_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__a221oi_2 _22106_ (.A1(_05277_),
    .A2(\line_cache[43][7] ),
    .B1(\line_cache[44][7] ),
    .B2(_05287_),
    .C1(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__or3b_1 _22107_ (.A(_07474_),
    .B(_07475_),
    .C_N(_07479_),
    .X(_07480_));
 sky130_fd_sc_hd__a22o_1 _22108_ (.A1(_05106_),
    .A2(\line_cache[317][7] ),
    .B1(\line_cache[316][7] ),
    .B2(_05108_),
    .X(_07481_));
 sky130_fd_sc_hd__a22o_1 _22109_ (.A1(_05292_),
    .A2(\line_cache[61][7] ),
    .B1(\line_cache[60][7] ),
    .B2(_05294_),
    .X(_07482_));
 sky130_fd_sc_hd__a22o_1 _22110_ (.A1(_05312_),
    .A2(\line_cache[58][7] ),
    .B1(_05317_),
    .B2(\line_cache[59][7] ),
    .X(_07483_));
 sky130_fd_sc_hd__and3_1 _22111_ (.A(_05109_),
    .B(_05021_),
    .C(\line_cache[318][7] ),
    .X(_07484_));
 sky130_fd_sc_hd__a21o_1 _22112_ (.A1(\line_cache[62][7] ),
    .A2(_05296_),
    .B1(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__or4_1 _22113_ (.A(_07481_),
    .B(_07482_),
    .C(_07483_),
    .D(_07485_),
    .X(_07486_));
 sky130_fd_sc_hd__a22o_1 _22114_ (.A1(_05129_),
    .A2(\line_cache[304][7] ),
    .B1(\line_cache[305][7] ),
    .B2(_05127_),
    .X(_07487_));
 sky130_fd_sc_hd__a22o_1 _22115_ (.A1(_05119_),
    .A2(\line_cache[312][7] ),
    .B1(\line_cache[313][7] ),
    .B2(_05121_),
    .X(_07488_));
 sky130_fd_sc_hd__a22o_1 _22116_ (.A1(_05123_),
    .A2(\line_cache[314][7] ),
    .B1(_05644_),
    .B2(\line_cache[315][7] ),
    .X(_07489_));
 sky130_fd_sc_hd__a22o_1 _22117_ (.A1(_05132_),
    .A2(\line_cache[306][7] ),
    .B1(\line_cache[307][7] ),
    .B2(_05136_),
    .X(_07490_));
 sky130_fd_sc_hd__or4_2 _22118_ (.A(_07487_),
    .B(_07488_),
    .C(_07489_),
    .D(_07490_),
    .X(_07491_));
 sky130_fd_sc_hd__a22o_1 _22119_ (.A1(_05314_),
    .A2(\line_cache[56][7] ),
    .B1(\line_cache[57][7] ),
    .B2(_05315_),
    .X(_07492_));
 sky130_fd_sc_hd__a22o_1 _22120_ (.A1(_05304_),
    .A2(\line_cache[52][7] ),
    .B1(\line_cache[53][7] ),
    .B2(_05306_),
    .X(_07493_));
 sky130_fd_sc_hd__a22o_1 _22121_ (.A1(_05301_),
    .A2(\line_cache[50][7] ),
    .B1(\line_cache[51][7] ),
    .B2(_05302_),
    .X(_07494_));
 sky130_fd_sc_hd__a22o_1 _22122_ (.A1(_05307_),
    .A2(\line_cache[54][7] ),
    .B1(_05309_),
    .B2(\line_cache[55][7] ),
    .X(_07495_));
 sky130_fd_sc_hd__or4_1 _22123_ (.A(_07492_),
    .B(_07493_),
    .C(_07494_),
    .D(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__or4_1 _22124_ (.A(_07480_),
    .B(_07486_),
    .C(_07491_),
    .D(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__or2b_1 _22125_ (.A(_05365_),
    .B_N(\line_cache[12][7] ),
    .X(_07498_));
 sky130_fd_sc_hd__nand2_1 _22126_ (.A(_05358_),
    .B(\line_cache[11][7] ),
    .Y(_07499_));
 sky130_fd_sc_hd__nand2_1 _22127_ (.A(_07498_),
    .B(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__a221oi_1 _22128_ (.A1(\line_cache[14][7] ),
    .A2(_05838_),
    .B1(\line_cache[13][7] ),
    .B2(_05839_),
    .C1(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__nand2_1 _22129_ (.A(_05353_),
    .B(\line_cache[10][7] ),
    .Y(_07502_));
 sky130_fd_sc_hd__nand2_1 _22130_ (.A(_05351_),
    .B(\line_cache[9][7] ),
    .Y(_07503_));
 sky130_fd_sc_hd__nand2_1 _22131_ (.A(_07502_),
    .B(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__a221oi_1 _22132_ (.A1(_05355_),
    .A2(\line_cache[8][7] ),
    .B1(_05346_),
    .B2(\line_cache[7][7] ),
    .C1(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__nand2_1 _22133_ (.A(_07501_),
    .B(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__and3_1 _22134_ (.A(_05163_),
    .B(_05187_),
    .C(\line_cache[21][7] ),
    .X(_07507_));
 sky130_fd_sc_hd__and3_1 _22135_ (.A(_05167_),
    .B(_05187_),
    .C(\line_cache[20][7] ),
    .X(_07508_));
 sky130_fd_sc_hd__a22o_1 _22136_ (.A1(_05825_),
    .A2(\line_cache[23][7] ),
    .B1(\line_cache[22][7] ),
    .B2(_05826_),
    .X(_07509_));
 sky130_fd_sc_hd__a22o_1 _22137_ (.A1(_05329_),
    .A2(\line_cache[16][7] ),
    .B1(\line_cache[17][7] ),
    .B2(_05330_),
    .X(_07510_));
 sky130_fd_sc_hd__a221o_1 _22138_ (.A1(\line_cache[19][7] ),
    .A2(_05831_),
    .B1(\line_cache[18][7] ),
    .B2(_05832_),
    .C1(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__or4_1 _22139_ (.A(_07507_),
    .B(_07508_),
    .C(_07509_),
    .D(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__a22o_1 _22140_ (.A1(_05262_),
    .A2(\line_cache[33][7] ),
    .B1(\line_cache[34][7] ),
    .B2(_05263_),
    .X(_07513_));
 sky130_fd_sc_hd__a221o_1 _22141_ (.A1(\line_cache[36][7] ),
    .A2(_05266_),
    .B1(\line_cache[35][7] ),
    .B2(_05261_),
    .C1(_07513_),
    .X(_07514_));
 sky130_fd_sc_hd__and3_1 _22142_ (.A(_05146_),
    .B(_05186_),
    .C(\line_cache[25][7] ),
    .X(_07515_));
 sky130_fd_sc_hd__a31o_1 _22143_ (.A1(_05991_),
    .A2(\line_cache[24][7] ),
    .A3(_05320_),
    .B1(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__a221oi_2 _22144_ (.A1(\line_cache[27][7] ),
    .A2(_05817_),
    .B1(\line_cache[26][7] ),
    .B2(_05819_),
    .C1(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__a32o_1 _22145_ (.A1(_05175_),
    .A2(_05812_),
    .A3(\line_cache[30][7] ),
    .B1(_05260_),
    .B2(\line_cache[32][7] ),
    .X(_07518_));
 sky130_fd_sc_hd__a32o_1 _22146_ (.A1(_05991_),
    .A2(_05173_),
    .A3(\line_cache[29][7] ),
    .B1(_06051_),
    .B2(\line_cache[28][7] ),
    .X(_07519_));
 sky130_fd_sc_hd__nor2_1 _22147_ (.A(_07518_),
    .B(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__nand2_1 _22148_ (.A(_05270_),
    .B(\line_cache[38][7] ),
    .Y(_07521_));
 sky130_fd_sc_hd__nand2_1 _22149_ (.A(_05272_),
    .B(\line_cache[37][7] ),
    .Y(_07522_));
 sky130_fd_sc_hd__nand2_1 _22150_ (.A(_07521_),
    .B(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__a221oi_2 _22151_ (.A1(_05268_),
    .A2(\line_cache[39][7] ),
    .B1(\line_cache[40][7] ),
    .B2(_05275_),
    .C1(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__and4b_1 _22152_ (.A_N(_07514_),
    .B(_07517_),
    .C(_07520_),
    .D(_07524_),
    .X(_07525_));
 sky130_fd_sc_hd__or3b_2 _22153_ (.A(_07506_),
    .B(_07512_),
    .C_N(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__nor3_2 _22154_ (.A(_07473_),
    .B(_07497_),
    .C(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__and3_1 _22155_ (.A(_05058_),
    .B(_05034_),
    .C(\line_cache[302][7] ),
    .X(_07528_));
 sky130_fd_sc_hd__a22o_1 _22156_ (.A1(_05056_),
    .A2(\line_cache[301][7] ),
    .B1(\line_cache[300][7] ),
    .B2(_05053_),
    .X(_07529_));
 sky130_fd_sc_hd__a211o_1 _22157_ (.A1(\line_cache[256][7] ),
    .A2(_05777_),
    .B1(_07528_),
    .C1(_07529_),
    .X(_07530_));
 sky130_fd_sc_hd__and3_1 _22158_ (.A(_05779_),
    .B(_05021_),
    .C(\line_cache[258][7] ),
    .X(_07531_));
 sky130_fd_sc_hd__and3_1 _22159_ (.A(_05771_),
    .B(_05034_),
    .C(\line_cache[260][7] ),
    .X(_07532_));
 sky130_fd_sc_hd__and3_1 _22160_ (.A(_05778_),
    .B(_05176_),
    .C(\line_cache[259][7] ),
    .X(_07533_));
 sky130_fd_sc_hd__a2111o_1 _22161_ (.A1(\line_cache[257][7] ),
    .A2(_05776_),
    .B1(_07531_),
    .C1(_07532_),
    .D1(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__and3_1 _22162_ (.A(_05356_),
    .B(_05176_),
    .C(\line_cache[267][7] ),
    .X(_07535_));
 sky130_fd_sc_hd__a22o_1 _22163_ (.A1(_05760_),
    .A2(\line_cache[266][7] ),
    .B1(\line_cache[265][7] ),
    .B2(_05764_),
    .X(_07536_));
 sky130_fd_sc_hd__a311o_1 _22164_ (.A1(_05113_),
    .A2(\line_cache[268][7] ),
    .A3(_05364_),
    .B1(_07535_),
    .C1(_07536_),
    .X(_07537_));
 sky130_fd_sc_hd__nand2_1 _22165_ (.A(_05768_),
    .B(\line_cache[262][7] ),
    .Y(_07538_));
 sky130_fd_sc_hd__nand2_1 _22166_ (.A(_05773_),
    .B(\line_cache[261][7] ),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_1 _22167_ (.A(_07538_),
    .B(_07539_),
    .Y(_07540_));
 sky130_fd_sc_hd__a221oi_2 _22168_ (.A1(_05763_),
    .A2(\line_cache[264][7] ),
    .B1(_05770_),
    .B2(\line_cache[263][7] ),
    .C1(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__or4b_1 _22169_ (.A(_07530_),
    .B(_07534_),
    .C(_07537_),
    .D_N(_07541_),
    .X(_07542_));
 sky130_fd_sc_hd__a22o_1 _22170_ (.A1(_05098_),
    .A2(\line_cache[308][7] ),
    .B1(\line_cache[309][7] ),
    .B2(_05093_),
    .X(_07543_));
 sky130_fd_sc_hd__a221o_1 _22171_ (.A1(\line_cache[311][7] ),
    .A2(_05097_),
    .B1(\line_cache[310][7] ),
    .B2(_05103_),
    .C1(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__a22o_1 _22172_ (.A1(_05046_),
    .A2(\line_cache[295][7] ),
    .B1(\line_cache[294][7] ),
    .B2(_05043_),
    .X(_07545_));
 sky130_fd_sc_hd__a221o_1 _22173_ (.A1(\line_cache[293][7] ),
    .A2(_05628_),
    .B1(\line_cache[292][7] ),
    .B2(_05627_),
    .C1(_07545_),
    .X(_07546_));
 sky130_fd_sc_hd__a22o_1 _22174_ (.A1(_05069_),
    .A2(\line_cache[296][7] ),
    .B1(\line_cache[297][7] ),
    .B2(_05076_),
    .X(_07547_));
 sky130_fd_sc_hd__a221o_1 _22175_ (.A1(\line_cache[299][7] ),
    .A2(_05073_),
    .B1(\line_cache[298][7] ),
    .B2(_05079_),
    .C1(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__a22o_1 _22176_ (.A1(_05632_),
    .A2(\line_cache[288][7] ),
    .B1(\line_cache[289][7] ),
    .B2(_05633_),
    .X(_07549_));
 sky130_fd_sc_hd__a221o_1 _22177_ (.A1(\line_cache[291][7] ),
    .A2(_05623_),
    .B1(\line_cache[290][7] ),
    .B2(_05624_),
    .C1(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__or4_1 _22178_ (.A(_07544_),
    .B(_07546_),
    .C(_07548_),
    .D(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__nor2_1 _22179_ (.A(_07542_),
    .B(_07551_),
    .Y(_07552_));
 sky130_fd_sc_hd__and3_1 _22180_ (.A(_05203_),
    .B(\line_cache[203][7] ),
    .C(_05471_),
    .X(_07553_));
 sky130_fd_sc_hd__and3_1 _22181_ (.A(_05586_),
    .B(\line_cache[206][7] ),
    .C(_05471_),
    .X(_07554_));
 sky130_fd_sc_hd__and2b_1 _22182_ (.A_N(_05687_),
    .B(\line_cache[204][7] ),
    .X(_07555_));
 sky130_fd_sc_hd__a2111o_1 _22183_ (.A1(\line_cache[205][7] ),
    .A2(_05683_),
    .B1(_07553_),
    .C1(_07554_),
    .D1(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__a22o_1 _22184_ (.A1(_05484_),
    .A2(\line_cache[195][7] ),
    .B1(_05485_),
    .B2(\line_cache[196][7] ),
    .X(_07557_));
 sky130_fd_sc_hd__a221o_1 _22185_ (.A1(\line_cache[198][7] ),
    .A2(_05487_),
    .B1(\line_cache[197][7] ),
    .B2(_05489_),
    .C1(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__a22o_1 _22186_ (.A1(_05495_),
    .A2(\line_cache[200][7] ),
    .B1(_05493_),
    .B2(\line_cache[199][7] ),
    .X(_07559_));
 sky130_fd_sc_hd__a221o_1 _22187_ (.A1(\line_cache[202][7] ),
    .A2(_05492_),
    .B1(\line_cache[201][7] ),
    .B2(_05491_),
    .C1(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__and3_1 _22188_ (.A(_05470_),
    .B(\line_cache[193][7] ),
    .C(_05685_),
    .X(_07561_));
 sky130_fd_sc_hd__and3_1 _22189_ (.A(_05475_),
    .B(\line_cache[192][7] ),
    .C(_05685_),
    .X(_07562_));
 sky130_fd_sc_hd__and3_1 _22190_ (.A(_05408_),
    .B(\line_cache[194][7] ),
    .C(_05472_),
    .X(_07563_));
 sky130_fd_sc_hd__a2111o_1 _22191_ (.A1(_05630_),
    .A2(\line_cache[286][7] ),
    .B1(_07561_),
    .C1(_07562_),
    .D1(_07563_),
    .X(_07564_));
 sky130_fd_sc_hd__or4_1 _22192_ (.A(_07556_),
    .B(_07558_),
    .C(_07560_),
    .D(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__a22o_1 _22193_ (.A1(_05659_),
    .A2(\line_cache[275][7] ),
    .B1(\line_cache[274][7] ),
    .B2(_05662_),
    .X(_07566_));
 sky130_fd_sc_hd__a22o_1 _22194_ (.A1(_05658_),
    .A2(\line_cache[276][7] ),
    .B1(\line_cache[277][7] ),
    .B2(_05655_),
    .X(_07567_));
 sky130_fd_sc_hd__a22o_1 _22195_ (.A1(_05668_),
    .A2(\line_cache[270][7] ),
    .B1(\line_cache[269][7] ),
    .B2(_05670_),
    .X(_07568_));
 sky130_fd_sc_hd__a221o_1 _22196_ (.A1(\line_cache[273][7] ),
    .A2(_05660_),
    .B1(\line_cache[272][7] ),
    .B2(_05666_),
    .C1(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__a22oi_1 _22197_ (.A1(_05676_),
    .A2(\line_cache[283][7] ),
    .B1(_05678_),
    .B2(\line_cache[282][7] ),
    .Y(_07570_));
 sky130_fd_sc_hd__a22oi_1 _22198_ (.A1(_05674_),
    .A2(\line_cache[284][7] ),
    .B1(_05631_),
    .B2(\line_cache[285][7] ),
    .Y(_07571_));
 sky130_fd_sc_hd__nand2_1 _22199_ (.A(_07570_),
    .B(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__a22o_1 _22200_ (.A1(_05144_),
    .A2(\line_cache[280][7] ),
    .B1(_05677_),
    .B2(\line_cache[281][7] ),
    .X(_07573_));
 sky130_fd_sc_hd__a32o_1 _22201_ (.A1(_05165_),
    .A2(_05151_),
    .A3(\line_cache[278][7] ),
    .B1(_05654_),
    .B2(\line_cache[279][7] ),
    .X(_07574_));
 sky130_fd_sc_hd__nor3_1 _22202_ (.A(_07572_),
    .B(_07573_),
    .C(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__or4b_2 _22203_ (.A(_07566_),
    .B(_07567_),
    .C(_07569_),
    .D_N(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__nor2_1 _22204_ (.A(_07565_),
    .B(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__a22o_1 _22205_ (.A1(_05746_),
    .A2(\line_cache[236][7] ),
    .B1(_05747_),
    .B2(\line_cache[235][7] ),
    .X(_07578_));
 sky130_fd_sc_hd__a221o_1 _22206_ (.A1(\line_cache[238][7] ),
    .A2(_05744_),
    .B1(\line_cache[237][7] ),
    .B2(_05745_),
    .C1(_07578_),
    .X(_07579_));
 sky130_fd_sc_hd__and3_1 _22207_ (.A(_05469_),
    .B(\line_cache[225][7] ),
    .C(_05732_),
    .X(_07580_));
 sky130_fd_sc_hd__and3_1 _22208_ (.A(_05408_),
    .B(\line_cache[226][7] ),
    .C(_05721_),
    .X(_07581_));
 sky130_fd_sc_hd__and3_1 _22209_ (.A(_05475_),
    .B(\line_cache[224][7] ),
    .C(_05721_),
    .X(_07582_));
 sky130_fd_sc_hd__a2111o_1 _22210_ (.A1(\line_cache[223][7] ),
    .A2(_05720_),
    .B1(_07580_),
    .C1(_07581_),
    .D1(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__and3_1 _22211_ (.A(_05704_),
    .B(\line_cache[227][7] ),
    .C(_05193_),
    .X(_07584_));
 sky130_fd_sc_hd__and3_1 _22212_ (.A(_05610_),
    .B(\line_cache[228][7] ),
    .C(_05193_),
    .X(_07585_));
 sky130_fd_sc_hd__and3_1 _22213_ (.A(_05710_),
    .B(\line_cache[229][7] ),
    .C(_05193_),
    .X(_07586_));
 sky130_fd_sc_hd__and3_1 _22214_ (.A(_05708_),
    .B(\line_cache[230][7] ),
    .C(_05732_),
    .X(_07587_));
 sky130_fd_sc_hd__or4_1 _22215_ (.A(_07584_),
    .B(_07585_),
    .C(_07586_),
    .D(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__a22o_1 _22216_ (.A1(_05728_),
    .A2(\line_cache[232][7] ),
    .B1(_05729_),
    .B2(\line_cache[231][7] ),
    .X(_07589_));
 sky130_fd_sc_hd__a221o_1 _22217_ (.A1(\line_cache[234][7] ),
    .A2(_05726_),
    .B1(\line_cache[233][7] ),
    .B2(_05727_),
    .C1(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__or4_1 _22218_ (.A(_07579_),
    .B(_07583_),
    .C(_07588_),
    .D(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__a22o_1 _22219_ (.A1(_05716_),
    .A2(\line_cache[220][7] ),
    .B1(_05717_),
    .B2(\line_cache[219][7] ),
    .X(_07592_));
 sky130_fd_sc_hd__a221o_1 _22220_ (.A1(\line_cache[222][7] ),
    .A2(_05714_),
    .B1(\line_cache[221][7] ),
    .B2(_05715_),
    .C1(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__a22o_1 _22221_ (.A1(_05700_),
    .A2(\line_cache[209][7] ),
    .B1(\line_cache[210][7] ),
    .B2(_05701_),
    .X(_07594_));
 sky130_fd_sc_hd__a221o_1 _22222_ (.A1(\line_cache[208][7] ),
    .A2(_05698_),
    .B1(\line_cache[207][7] ),
    .B2(_05699_),
    .C1(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__and3_1 _22223_ (.A(_05704_),
    .B(\line_cache[211][7] ),
    .C(_05693_),
    .X(_07596_));
 sky130_fd_sc_hd__and3_1 _22224_ (.A(_05610_),
    .B(\line_cache[212][7] ),
    .C(_05694_),
    .X(_07597_));
 sky130_fd_sc_hd__and3_1 _22225_ (.A(_05710_),
    .B(\line_cache[213][7] ),
    .C(_05694_),
    .X(_07598_));
 sky130_fd_sc_hd__and3_1 _22226_ (.A(_05708_),
    .B(\line_cache[214][7] ),
    .C(_05706_),
    .X(_07599_));
 sky130_fd_sc_hd__or4_1 _22227_ (.A(_07596_),
    .B(_07597_),
    .C(_07598_),
    .D(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__a22o_1 _22228_ (.A1(_05692_),
    .A2(\line_cache[216][7] ),
    .B1(_05983_),
    .B2(\line_cache[215][7] ),
    .X(_07601_));
 sky130_fd_sc_hd__a221o_1 _22229_ (.A1(\line_cache[218][7] ),
    .A2(_05690_),
    .B1(\line_cache[217][7] ),
    .B2(_05691_),
    .C1(_07601_),
    .X(_07602_));
 sky130_fd_sc_hd__or4_2 _22230_ (.A(_07593_),
    .B(_07595_),
    .C(_07600_),
    .D(_07602_),
    .X(_07603_));
 sky130_fd_sc_hd__nor2_1 _22231_ (.A(_07591_),
    .B(_07603_),
    .Y(_07604_));
 sky130_fd_sc_hd__and3_1 _22232_ (.A(_05454_),
    .B(\line_cache[239][7] ),
    .C(_05732_),
    .X(_07605_));
 sky130_fd_sc_hd__and3_1 _22233_ (.A(_05469_),
    .B(\line_cache[241][7] ),
    .C(_05206_),
    .X(_07606_));
 sky130_fd_sc_hd__and3_1 _22234_ (.A(_05408_),
    .B(\line_cache[242][7] ),
    .C(_05206_),
    .X(_07607_));
 sky130_fd_sc_hd__a2111o_1 _22235_ (.A1(_05233_),
    .A2(\line_cache[240][7] ),
    .B1(_07605_),
    .C1(_07606_),
    .D1(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__and2_1 _22236_ (.A(_05235_),
    .B(\line_cache[243][7] ),
    .X(_07609_));
 sky130_fd_sc_hd__a21o_1 _22237_ (.A1(\line_cache[244][7] ),
    .A2(_05224_),
    .B1(_07609_),
    .X(_07610_));
 sky130_fd_sc_hd__a221o_1 _22238_ (.A1(\line_cache[246][7] ),
    .A2(_05753_),
    .B1(\line_cache[245][7] ),
    .B2(_05226_),
    .C1(_07610_),
    .X(_07611_));
 sky130_fd_sc_hd__a22o_1 _22239_ (.A1(_05212_),
    .A2(\line_cache[252][7] ),
    .B1(_05205_),
    .B2(\line_cache[251][7] ),
    .X(_07612_));
 sky130_fd_sc_hd__a221o_1 _22240_ (.A1(\line_cache[254][7] ),
    .A2(_05217_),
    .B1(\line_cache[253][7] ),
    .B2(_05214_),
    .C1(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__a22o_1 _22241_ (.A1(_05750_),
    .A2(\line_cache[248][7] ),
    .B1(_05229_),
    .B2(\line_cache[247][7] ),
    .X(_07614_));
 sky130_fd_sc_hd__a221o_1 _22242_ (.A1(\line_cache[250][7] ),
    .A2(_05202_),
    .B1(\line_cache[249][7] ),
    .B2(_05209_),
    .C1(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__or4_1 _22243_ (.A(_07608_),
    .B(_07611_),
    .C(_07613_),
    .D(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__a22o_1 _22244_ (.A1(_05875_),
    .A2(\line_cache[67][7] ),
    .B1(_05861_),
    .B2(\line_cache[66][7] ),
    .X(_07617_));
 sky130_fd_sc_hd__a221o_1 _22245_ (.A1(\line_cache[65][7] ),
    .A2(_05860_),
    .B1(\line_cache[64][7] ),
    .B2(_05858_),
    .C1(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__a22o_1 _22246_ (.A1(_05867_),
    .A2(\line_cache[72][7] ),
    .B1(_05866_),
    .B2(\line_cache[73][7] ),
    .X(_07619_));
 sky130_fd_sc_hd__a221o_1 _22247_ (.A1(\line_cache[75][7] ),
    .A2(_05543_),
    .B1(\line_cache[74][7] ),
    .B2(_05865_),
    .C1(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__a22o_1 _22248_ (.A1(_05873_),
    .A2(\line_cache[68][7] ),
    .B1(_05872_),
    .B2(\line_cache[69][7] ),
    .X(_07621_));
 sky130_fd_sc_hd__a221o_1 _22249_ (.A1(\line_cache[71][7] ),
    .A2(_05868_),
    .B1(\line_cache[70][7] ),
    .B2(_05871_),
    .C1(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__and2_1 _22250_ (.A(_05542_),
    .B(\line_cache[76][7] ),
    .X(_07623_));
 sky130_fd_sc_hd__and3_1 _22251_ (.A(_05544_),
    .B(\line_cache[77][7] ),
    .C(_05536_),
    .X(_07624_));
 sky130_fd_sc_hd__or2_1 _22252_ (.A(_07623_),
    .B(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__a221o_1 _22253_ (.A1(\line_cache[79][7] ),
    .A2(_05537_),
    .B1(\line_cache[78][7] ),
    .B2(_05545_),
    .C1(_07625_),
    .X(_07626_));
 sky130_fd_sc_hd__or4_2 _22254_ (.A(_07618_),
    .B(_07620_),
    .C(_07622_),
    .D(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__nor2_1 _22255_ (.A(_07616_),
    .B(_07627_),
    .Y(_07628_));
 sky130_fd_sc_hd__and4_1 _22256_ (.A(_07552_),
    .B(_07577_),
    .C(_07604_),
    .D(_07628_),
    .X(_07629_));
 sky130_fd_sc_hd__nand3_1 _22257_ (.A(_07459_),
    .B(_07527_),
    .C(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__o21a_4 _22258_ (.A1(_07381_),
    .A2(_07630_),
    .B1(_05884_),
    .X(net133));
 sky130_fd_sc_hd__or2_1 _22259_ (.A(net4215),
    .B(net125),
    .X(_07631_));
 sky130_fd_sc_hd__clkbuf_1 _22260_ (.A(net4216),
    .X(_02572_));
 sky130_fd_sc_hd__inv_2 _22261_ (.A(net4215),
    .Y(_07632_));
 sky130_fd_sc_hd__nor2_2 _22262_ (.A(_08726_),
    .B(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__o21a_1 _22263_ (.A1(net4221),
    .A2(_07633_),
    .B1(_08771_),
    .X(_02573_));
 sky130_fd_sc_hd__nand2_1 _22264_ (.A(net2713),
    .B(_09359_),
    .Y(_07634_));
 sky130_fd_sc_hd__inv_2 _22265_ (.A(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__mux2_1 _22266_ (.A0(_07635_),
    .A1(_08728_),
    .S(net4297),
    .X(_07636_));
 sky130_fd_sc_hd__clkbuf_1 _22267_ (.A(_07636_),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_1 _22268_ (.A(_10040_),
    .B(_10095_),
    .Y(_07637_));
 sky130_fd_sc_hd__a22o_1 _22269_ (.A1(net2781),
    .A2(_08728_),
    .B1(_07635_),
    .B2(_07637_),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_1 _22270_ (.A(_09173_),
    .B(net3791),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_1 _22271_ (.A(_09172_),
    .B(_08756_),
    .Y(_07639_));
 sky130_fd_sc_hd__a32o_1 _22272_ (.A1(_07635_),
    .A2(_07638_),
    .A3(_07639_),
    .B1(net3791),
    .B2(_08728_),
    .X(_02576_));
 sky130_fd_sc_hd__nor2_1 _22273_ (.A(_09167_),
    .B(_09172_),
    .Y(_07640_));
 sky130_fd_sc_hd__inv_2 _22274_ (.A(_07640_),
    .Y(_07641_));
 sky130_fd_sc_hd__nand2_1 _22275_ (.A(_07638_),
    .B(_08758_),
    .Y(_07642_));
 sky130_fd_sc_hd__a32o_1 _22276_ (.A1(_07635_),
    .A2(_07641_),
    .A3(_07642_),
    .B1(net2787),
    .B2(_08728_),
    .X(_02577_));
 sky130_fd_sc_hd__nand2_1 _22277_ (.A(_07640_),
    .B(net3899),
    .Y(_07643_));
 sky130_fd_sc_hd__nand2_1 _22278_ (.A(_07641_),
    .B(_03162_),
    .Y(_07644_));
 sky130_fd_sc_hd__a32o_1 _22279_ (.A1(_07635_),
    .A2(_07643_),
    .A3(_07644_),
    .B1(net3899),
    .B2(_08728_),
    .X(_02578_));
 sky130_fd_sc_hd__inv_2 _22280_ (.A(_10234_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand2_1 _22281_ (.A(_07643_),
    .B(_08738_),
    .Y(_07646_));
 sky130_fd_sc_hd__a32o_1 _22282_ (.A1(_07635_),
    .A2(_07645_),
    .A3(_07646_),
    .B1(net2927),
    .B2(_08728_),
    .X(_02579_));
 sky130_fd_sc_hd__a31o_1 _22283_ (.A1(_07640_),
    .A2(_04828_),
    .A3(_10466_),
    .B1(_09444_),
    .X(_07647_));
 sky130_fd_sc_hd__o2bb2a_1 _22284_ (.A1_N(_10238_),
    .A2_N(_07647_),
    .B1(_08728_),
    .B2(net2713),
    .X(_02580_));
 sky130_fd_sc_hd__and3_1 _22285_ (.A(_10234_),
    .B(_08736_),
    .C(_09225_),
    .X(_07648_));
 sky130_fd_sc_hd__nand2_1 _22286_ (.A(_07648_),
    .B(net4281),
    .Y(_07649_));
 sky130_fd_sc_hd__or2_1 _22287_ (.A(net4281),
    .B(_07648_),
    .X(_07650_));
 sky130_fd_sc_hd__and3_1 _22288_ (.A(_08771_),
    .B(_07649_),
    .C(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__clkbuf_1 _22289_ (.A(_07651_),
    .X(_02581_));
 sky130_fd_sc_hd__inv_2 _22290_ (.A(net3018),
    .Y(_07652_));
 sky130_fd_sc_hd__inv_2 _22291_ (.A(net3517),
    .Y(_07653_));
 sky130_fd_sc_hd__inv_2 _22292_ (.A(net2729),
    .Y(_07654_));
 sky130_fd_sc_hd__inv_2 _22293_ (.A(net2668),
    .Y(_07655_));
 sky130_fd_sc_hd__and4_1 _22294_ (.A(_07652_),
    .B(_07653_),
    .C(_07654_),
    .D(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__nor2_1 _22295_ (.A(net2687),
    .B(net2685),
    .Y(_07657_));
 sky130_fd_sc_hd__nor2_1 _22296_ (.A(net2778),
    .B(\res_v_counter[0] ),
    .Y(_07658_));
 sky130_fd_sc_hd__inv_2 _22297_ (.A(net2826),
    .Y(_07659_));
 sky130_fd_sc_hd__inv_2 _22298_ (.A(net2691),
    .Y(_07660_));
 sky130_fd_sc_hd__and3_1 _22299_ (.A(_07658_),
    .B(_07659_),
    .C(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__a31o_4 _22300_ (.A1(_07656_),
    .A2(_07657_),
    .A3(_07661_),
    .B1(_07632_),
    .X(_07662_));
 sky130_fd_sc_hd__or2_4 _22301_ (.A(_09225_),
    .B(_07633_),
    .X(_07663_));
 sky130_fd_sc_hd__nand2_8 _22302_ (.A(_07662_),
    .B(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__clkinv_4 _22303_ (.A(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__nand2_1 _22304_ (.A(_07665_),
    .B(_08726_),
    .Y(_07666_));
 sky130_fd_sc_hd__inv_2 _22305_ (.A(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__buf_4 _22306_ (.A(_07665_),
    .X(_07668_));
 sky130_fd_sc_hd__nand2_1 _22307_ (.A(_07668_),
    .B(net2716),
    .Y(_07669_));
 sky130_fd_sc_hd__o21a_1 _22308_ (.A1(net2716),
    .A2(_07667_),
    .B1(_07669_),
    .X(_02582_));
 sky130_fd_sc_hd__nand2_1 _22309_ (.A(net2716),
    .B(net4270),
    .Y(_07670_));
 sky130_fd_sc_hd__or2_1 _22310_ (.A(net2716),
    .B(net4270),
    .X(_07671_));
 sky130_fd_sc_hd__and2_1 _22311_ (.A(_07664_),
    .B(net4270),
    .X(_07672_));
 sky130_fd_sc_hd__a41o_1 _22312_ (.A1(_07668_),
    .A2(_08791_),
    .A3(_07670_),
    .A4(_07671_),
    .B1(_07672_),
    .X(_02583_));
 sky130_fd_sc_hd__or2_1 _22313_ (.A(_07670_),
    .B(_07664_),
    .X(_07673_));
 sky130_fd_sc_hd__inv_2 _22314_ (.A(net2741),
    .Y(_07674_));
 sky130_fd_sc_hd__nand2_4 _22315_ (.A(_07665_),
    .B(_09192_),
    .Y(_07675_));
 sky130_fd_sc_hd__inv_2 _22316_ (.A(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__or2_1 _22317_ (.A(_07674_),
    .B(_07670_),
    .X(_07677_));
 sky130_fd_sc_hd__or2_1 _22318_ (.A(_07677_),
    .B(_07664_),
    .X(_07678_));
 sky130_fd_sc_hd__inv_2 _22319_ (.A(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__a211oi_1 _22320_ (.A1(_07673_),
    .A2(_07674_),
    .B1(_07676_),
    .C1(_07679_),
    .Y(_02584_));
 sky130_fd_sc_hd__nor2b_1 _22321_ (.A(_07677_),
    .B_N(net3129),
    .Y(_07680_));
 sky130_fd_sc_hd__nand2_1 _22322_ (.A(_07668_),
    .B(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__o211a_1 _22323_ (.A1(net3129),
    .A2(_07679_),
    .B1(_07675_),
    .C1(_07681_),
    .X(_02585_));
 sky130_fd_sc_hd__nand2_1 _22324_ (.A(_07680_),
    .B(net3795),
    .Y(_07682_));
 sky130_fd_sc_hd__a31o_1 _22325_ (.A1(_07662_),
    .A2(_07663_),
    .A3(_07680_),
    .B1(net3795),
    .X(_07683_));
 sky130_fd_sc_hd__o211a_1 _22326_ (.A1(_07664_),
    .A2(_07682_),
    .B1(_07675_),
    .C1(net3796),
    .X(_02586_));
 sky130_fd_sc_hd__a31o_1 _22327_ (.A1(_07665_),
    .A2(net3795),
    .A3(_07680_),
    .B1(net4331),
    .X(_07684_));
 sky130_fd_sc_hd__nand2b_1 _22328_ (.A_N(_07682_),
    .B(net4331),
    .Y(_07685_));
 sky130_fd_sc_hd__or2_1 _22329_ (.A(_07685_),
    .B(_07664_),
    .X(_07686_));
 sky130_fd_sc_hd__and3_1 _22330_ (.A(_07684_),
    .B(_07675_),
    .C(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__clkbuf_1 _22331_ (.A(net4332),
    .X(_02587_));
 sky130_fd_sc_hd__inv_2 _22332_ (.A(net2748),
    .Y(_07688_));
 sky130_fd_sc_hd__or2_1 _22333_ (.A(_07688_),
    .B(_07685_),
    .X(_07689_));
 sky130_fd_sc_hd__inv_2 _22334_ (.A(_07689_),
    .Y(_07690_));
 sky130_fd_sc_hd__nand2_1 _22335_ (.A(_07665_),
    .B(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__inv_2 _22336_ (.A(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__a211oi_1 _22337_ (.A1(_07686_),
    .A2(_07688_),
    .B1(_07676_),
    .C1(_07692_),
    .Y(_02588_));
 sky130_fd_sc_hd__nand2_1 _22338_ (.A(_07690_),
    .B(net2793),
    .Y(_07693_));
 sky130_fd_sc_hd__inv_2 _22339_ (.A(_07693_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand2_1 _22340_ (.A(_07694_),
    .B(_07665_),
    .Y(_07695_));
 sky130_fd_sc_hd__o211a_1 _22341_ (.A1(net2793),
    .A2(_07692_),
    .B1(_07675_),
    .C1(_07695_),
    .X(_02589_));
 sky130_fd_sc_hd__inv_2 _22342_ (.A(net2743),
    .Y(_07696_));
 sky130_fd_sc_hd__nor2_1 _22343_ (.A(_07696_),
    .B(_07695_),
    .Y(_07697_));
 sky130_fd_sc_hd__or2_1 _22344_ (.A(_07676_),
    .B(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__a21oi_1 _22345_ (.A1(_07696_),
    .A2(_07695_),
    .B1(_07698_),
    .Y(_02590_));
 sky130_fd_sc_hd__nand2_1 _22346_ (.A(net2743),
    .B(net2809),
    .Y(_07699_));
 sky130_fd_sc_hd__nor2_1 _22347_ (.A(_07699_),
    .B(_07693_),
    .Y(_07700_));
 sky130_fd_sc_hd__nand2_1 _22348_ (.A(_07700_),
    .B(_07665_),
    .Y(_07701_));
 sky130_fd_sc_hd__o211a_1 _22349_ (.A1(net2809),
    .A2(_07697_),
    .B1(_07675_),
    .C1(_07701_),
    .X(_02591_));
 sky130_fd_sc_hd__inv_2 _22350_ (.A(net3188),
    .Y(_07702_));
 sky130_fd_sc_hd__nor2_1 _22351_ (.A(_07702_),
    .B(_07701_),
    .Y(_07703_));
 sky130_fd_sc_hd__or2_1 _22352_ (.A(_07676_),
    .B(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__a21oi_1 _22353_ (.A1(_07702_),
    .A2(_07701_),
    .B1(_07704_),
    .Y(_02592_));
 sky130_fd_sc_hd__inv_2 _22354_ (.A(net2726),
    .Y(_07705_));
 sky130_fd_sc_hd__inv_2 _22355_ (.A(_07700_),
    .Y(_07706_));
 sky130_fd_sc_hd__or4_1 _22356_ (.A(_07702_),
    .B(_07705_),
    .C(_07664_),
    .D(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__o211a_1 _22357_ (.A1(net2726),
    .A2(_07703_),
    .B1(_07675_),
    .C1(_07707_),
    .X(_02593_));
 sky130_fd_sc_hd__inv_2 _22358_ (.A(net2956),
    .Y(_07708_));
 sky130_fd_sc_hd__or4_1 _22359_ (.A(_07702_),
    .B(_07705_),
    .C(_07708_),
    .D(_07706_),
    .X(_07709_));
 sky130_fd_sc_hd__nor2_1 _22360_ (.A(_07664_),
    .B(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__a211oi_1 _22361_ (.A1(_07707_),
    .A2(_07708_),
    .B1(_07676_),
    .C1(_07710_),
    .Y(_02594_));
 sky130_fd_sc_hd__nor2b_1 _22362_ (.A(_07709_),
    .B_N(net2734),
    .Y(_07711_));
 sky130_fd_sc_hd__nand2_1 _22363_ (.A(_07711_),
    .B(_07665_),
    .Y(_07712_));
 sky130_fd_sc_hd__o211a_1 _22364_ (.A1(net2734),
    .A2(_07710_),
    .B1(_07675_),
    .C1(_07712_),
    .X(_02595_));
 sky130_fd_sc_hd__inv_2 _22365_ (.A(net2887),
    .Y(_07713_));
 sky130_fd_sc_hd__nor2_1 _22366_ (.A(_07713_),
    .B(_07712_),
    .Y(_07714_));
 sky130_fd_sc_hd__or2_1 _22367_ (.A(_07676_),
    .B(_07714_),
    .X(_07715_));
 sky130_fd_sc_hd__a21oi_1 _22368_ (.A1(_07713_),
    .A2(_07712_),
    .B1(_07715_),
    .Y(_02596_));
 sky130_fd_sc_hd__inv_2 _22369_ (.A(net2765),
    .Y(_07716_));
 sky130_fd_sc_hd__or3b_1 _22370_ (.A(_07713_),
    .B(_07716_),
    .C_N(_07711_),
    .X(_07717_));
 sky130_fd_sc_hd__o221a_1 _22371_ (.A1(net2765),
    .A2(_07714_),
    .B1(_07664_),
    .B2(_07717_),
    .C1(_07675_),
    .X(_02597_));
 sky130_fd_sc_hd__nand2_1 _22372_ (.A(net2956),
    .B(net2734),
    .Y(_07718_));
 sky130_fd_sc_hd__or3_1 _22373_ (.A(_07702_),
    .B(_07705_),
    .C(_07699_),
    .X(_07719_));
 sky130_fd_sc_hd__or4_1 _22374_ (.A(_07713_),
    .B(_07716_),
    .C(_07718_),
    .D(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__nor2_2 _22375_ (.A(_07693_),
    .B(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__or2_1 _22376_ (.A(net4242),
    .B(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__nand2_1 _22377_ (.A(_07721_),
    .B(net4242),
    .Y(_07723_));
 sky130_fd_sc_hd__and2_1 _22378_ (.A(_07664_),
    .B(net4242),
    .X(_07724_));
 sky130_fd_sc_hd__a41o_1 _22379_ (.A1(_07722_),
    .A2(_08791_),
    .A3(_07723_),
    .A4(_07668_),
    .B1(_07724_),
    .X(_02598_));
 sky130_fd_sc_hd__nand2_1 _22380_ (.A(net109),
    .B(net2671),
    .Y(_07725_));
 sky130_fd_sc_hd__or2_1 _22381_ (.A(_07725_),
    .B(_07717_),
    .X(_07726_));
 sky130_fd_sc_hd__a21o_1 _22382_ (.A1(_07721_),
    .A2(net109),
    .B1(net2671),
    .X(_07727_));
 sky130_fd_sc_hd__a32o_1 _22383_ (.A1(_07726_),
    .A2(_07667_),
    .A3(_07727_),
    .B1(net2671),
    .B2(_07664_),
    .X(_02599_));
 sky130_fd_sc_hd__nor2_1 _22384_ (.A(_07664_),
    .B(_07726_),
    .Y(_07728_));
 sky130_fd_sc_hd__a21oi_1 _22385_ (.A1(_07728_),
    .A2(net2719),
    .B1(_07676_),
    .Y(_07729_));
 sky130_fd_sc_hd__o21a_1 _22386_ (.A1(net2719),
    .A2(_07728_),
    .B1(_07729_),
    .X(_02600_));
 sky130_fd_sc_hd__inv_2 _22387_ (.A(net4193),
    .Y(_07730_));
 sky130_fd_sc_hd__inv_2 _22388_ (.A(_07725_),
    .Y(_07731_));
 sky130_fd_sc_hd__and2_1 _22389_ (.A(_07721_),
    .B(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__nand2_1 _22390_ (.A(_07732_),
    .B(net2719),
    .Y(_07733_));
 sky130_fd_sc_hd__or2_1 _22391_ (.A(_07730_),
    .B(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__nand2_1 _22392_ (.A(_07733_),
    .B(_07730_),
    .Y(_07735_));
 sky130_fd_sc_hd__nor2_1 _22393_ (.A(_07730_),
    .B(_07668_),
    .Y(_07736_));
 sky130_fd_sc_hd__a41o_1 _22394_ (.A1(_07734_),
    .A2(_07735_),
    .A3(_08791_),
    .A4(_07668_),
    .B1(_07736_),
    .X(_02601_));
 sky130_fd_sc_hd__inv_2 _22395_ (.A(net4211),
    .Y(_07737_));
 sky130_fd_sc_hd__and3_1 _22396_ (.A(_07731_),
    .B(net2719),
    .C(net4193),
    .X(_07738_));
 sky130_fd_sc_hd__nand2_1 _22397_ (.A(_07721_),
    .B(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__or2_1 _22398_ (.A(_07737_),
    .B(_07739_),
    .X(_07740_));
 sky130_fd_sc_hd__nand2_1 _22399_ (.A(_07739_),
    .B(_07737_),
    .Y(_07741_));
 sky130_fd_sc_hd__nor2_1 _22400_ (.A(_07737_),
    .B(_07668_),
    .Y(_07742_));
 sky130_fd_sc_hd__a41o_1 _22401_ (.A1(_07740_),
    .A2(_08791_),
    .A3(_07741_),
    .A4(_07668_),
    .B1(_07742_),
    .X(_02602_));
 sky130_fd_sc_hd__inv_2 _22402_ (.A(net4182),
    .Y(_07743_));
 sky130_fd_sc_hd__or2_1 _22403_ (.A(_07743_),
    .B(_07740_),
    .X(_07744_));
 sky130_fd_sc_hd__nand2_1 _22404_ (.A(_07740_),
    .B(_07743_),
    .Y(_07745_));
 sky130_fd_sc_hd__nor2_1 _22405_ (.A(_07743_),
    .B(_07668_),
    .Y(_07746_));
 sky130_fd_sc_hd__a41o_1 _22406_ (.A1(_07744_),
    .A2(_07745_),
    .A3(_08791_),
    .A4(_07668_),
    .B1(_07746_),
    .X(_02603_));
 sky130_fd_sc_hd__inv_2 _22407_ (.A(net4179),
    .Y(_07747_));
 sky130_fd_sc_hd__nand2_1 _22408_ (.A(net4211),
    .B(net4182),
    .Y(_07748_));
 sky130_fd_sc_hd__or2_1 _22409_ (.A(_07748_),
    .B(_07739_),
    .X(_07749_));
 sky130_fd_sc_hd__or2_1 _22410_ (.A(_07747_),
    .B(_07749_),
    .X(_07750_));
 sky130_fd_sc_hd__nand2_1 _22411_ (.A(_07749_),
    .B(_07747_),
    .Y(_07751_));
 sky130_fd_sc_hd__nor2_1 _22412_ (.A(_07747_),
    .B(_07668_),
    .Y(_07752_));
 sky130_fd_sc_hd__a41o_1 _22413_ (.A1(_07750_),
    .A2(_07751_),
    .A3(_08791_),
    .A4(_07668_),
    .B1(_07752_),
    .X(_02604_));
 sky130_fd_sc_hd__inv_2 _22414_ (.A(net4223),
    .Y(_07753_));
 sky130_fd_sc_hd__or2_1 _22415_ (.A(_07753_),
    .B(_07750_),
    .X(_07754_));
 sky130_fd_sc_hd__nand2_1 _22416_ (.A(_07750_),
    .B(_07753_),
    .Y(_07755_));
 sky130_fd_sc_hd__nor2_1 _22417_ (.A(_07753_),
    .B(_07668_),
    .Y(_07756_));
 sky130_fd_sc_hd__a41o_1 _22418_ (.A1(_07754_),
    .A2(_08791_),
    .A3(_07755_),
    .A4(_07665_),
    .B1(_07756_),
    .X(_02605_));
 sky130_fd_sc_hd__inv_2 _22419_ (.A(net4273),
    .Y(_07757_));
 sky130_fd_sc_hd__and4b_1 _22420_ (.A_N(_07748_),
    .B(_07738_),
    .C(net4179),
    .D(net4223),
    .X(_07758_));
 sky130_fd_sc_hd__nand2_1 _22421_ (.A(_07721_),
    .B(_07758_),
    .Y(_07759_));
 sky130_fd_sc_hd__or2_1 _22422_ (.A(_07757_),
    .B(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__nand2_1 _22423_ (.A(_07759_),
    .B(_07757_),
    .Y(_07761_));
 sky130_fd_sc_hd__nor2_1 _22424_ (.A(_07757_),
    .B(_07668_),
    .Y(_07762_));
 sky130_fd_sc_hd__a41o_1 _22425_ (.A1(_07760_),
    .A2(_08791_),
    .A3(_07761_),
    .A4(_07665_),
    .B1(_07762_),
    .X(_02606_));
 sky130_fd_sc_hd__inv_2 _22426_ (.A(net4257),
    .Y(_07763_));
 sky130_fd_sc_hd__or2_1 _22427_ (.A(_07763_),
    .B(_07760_),
    .X(_07764_));
 sky130_fd_sc_hd__nand2_1 _22428_ (.A(_07760_),
    .B(_07763_),
    .Y(_07765_));
 sky130_fd_sc_hd__nor2_1 _22429_ (.A(_07763_),
    .B(_07668_),
    .Y(_07766_));
 sky130_fd_sc_hd__a41o_1 _22430_ (.A1(_07764_),
    .A2(_07765_),
    .A3(_08791_),
    .A4(_07665_),
    .B1(_07766_),
    .X(_02607_));
 sky130_fd_sc_hd__inv_2 _22431_ (.A(net4285),
    .Y(_07767_));
 sky130_fd_sc_hd__or2_1 _22432_ (.A(_07767_),
    .B(_07764_),
    .X(_07768_));
 sky130_fd_sc_hd__nand2_1 _22433_ (.A(_07764_),
    .B(_07767_),
    .Y(_07769_));
 sky130_fd_sc_hd__nor2_1 _22434_ (.A(_07767_),
    .B(_07668_),
    .Y(_07770_));
 sky130_fd_sc_hd__a41o_1 _22435_ (.A1(_07768_),
    .A2(_07769_),
    .A3(_08791_),
    .A4(_07665_),
    .B1(_07770_),
    .X(_02608_));
 sky130_fd_sc_hd__inv_2 _22436_ (.A(net2673),
    .Y(_07771_));
 sky130_fd_sc_hd__or2_1 _22437_ (.A(_07771_),
    .B(_07768_),
    .X(_07772_));
 sky130_fd_sc_hd__nand2_1 _22438_ (.A(_07768_),
    .B(_07771_),
    .Y(_07773_));
 sky130_fd_sc_hd__a32o_1 _22439_ (.A1(_07772_),
    .A2(_07667_),
    .A3(_07773_),
    .B1(net2673),
    .B2(_07664_),
    .X(_02609_));
 sky130_fd_sc_hd__inv_2 _22440_ (.A(net4333),
    .Y(_07774_));
 sky130_fd_sc_hd__or3_1 _22441_ (.A(_07774_),
    .B(_07664_),
    .C(_07772_),
    .X(_07775_));
 sky130_fd_sc_hd__o21ai_1 _22442_ (.A1(_07664_),
    .A2(_07772_),
    .B1(_07774_),
    .Y(_07776_));
 sky130_fd_sc_hd__and3_1 _22443_ (.A(_07775_),
    .B(_07675_),
    .C(_07776_),
    .X(_07777_));
 sky130_fd_sc_hd__clkbuf_1 _22444_ (.A(net4334),
    .X(_02610_));
 sky130_fd_sc_hd__or2_1 _22445_ (.A(net2839),
    .B(_07775_),
    .X(_07778_));
 sky130_fd_sc_hd__nand2_1 _22446_ (.A(_07775_),
    .B(net2839),
    .Y(_07779_));
 sky130_fd_sc_hd__a21oi_1 _22447_ (.A1(_07778_),
    .A2(net2840),
    .B1(_07676_),
    .Y(_02611_));
 sky130_fd_sc_hd__nor2_1 _22448_ (.A(net88),
    .B(net89),
    .Y(_07780_));
 sky130_fd_sc_hd__inv_2 _22449_ (.A(net91),
    .Y(_07781_));
 sky130_fd_sc_hd__and3_1 _22450_ (.A(_07780_),
    .B(net90),
    .C(_07781_),
    .X(_07782_));
 sky130_fd_sc_hd__buf_6 _22451_ (.A(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__or3b_2 _22452_ (.A(net90),
    .B(_07781_),
    .C_N(_07780_),
    .X(_07784_));
 sky130_fd_sc_hd__inv_6 _22453_ (.A(_07784_),
    .Y(_07785_));
 sky130_fd_sc_hd__nor2_8 _22454_ (.A(_07783_),
    .B(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__a22o_1 _22455_ (.A1(net32),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net33),
    .X(_07787_));
 sky130_fd_sc_hd__a21o_1 _22456_ (.A1(net31),
    .A2(_07786_),
    .B1(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__inv_2 _22457_ (.A(net88),
    .Y(_07789_));
 sky130_fd_sc_hd__nor2_1 _22458_ (.A(net90),
    .B(net91),
    .Y(_07790_));
 sky130_fd_sc_hd__inv_2 _22459_ (.A(_07786_),
    .Y(_07791_));
 sky130_fd_sc_hd__a31o_1 _22460_ (.A1(_07789_),
    .A2(net89),
    .A3(_07790_),
    .B1(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__nand2_1 _22461_ (.A(_07792_),
    .B(_08723_),
    .Y(_07793_));
 sky130_fd_sc_hd__buf_6 _22462_ (.A(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__mux2_1 _22463_ (.A0(_07788_),
    .A1(net3502),
    .S(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__clkbuf_1 _22464_ (.A(_07795_),
    .X(_02612_));
 sky130_fd_sc_hd__a22o_1 _22465_ (.A1(net33),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net34),
    .X(_07796_));
 sky130_fd_sc_hd__a21o_1 _22466_ (.A1(net32),
    .A2(_07786_),
    .B1(_07796_),
    .X(_07797_));
 sky130_fd_sc_hd__mux2_1 _22467_ (.A0(_07797_),
    .A1(net3527),
    .S(_07794_),
    .X(_07798_));
 sky130_fd_sc_hd__clkbuf_1 _22468_ (.A(_07798_),
    .X(_02613_));
 sky130_fd_sc_hd__inv_2 _22469_ (.A(net33),
    .Y(_07799_));
 sky130_fd_sc_hd__nor2_1 _22470_ (.A(_07799_),
    .B(_07791_),
    .Y(_07800_));
 sky130_fd_sc_hd__a221o_1 _22471_ (.A1(net34),
    .A2(_07783_),
    .B1(net35),
    .B2(_07785_),
    .C1(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__mux2_1 _22472_ (.A0(_07801_),
    .A1(net2745),
    .S(_07794_),
    .X(_07802_));
 sky130_fd_sc_hd__clkbuf_1 _22473_ (.A(_07802_),
    .X(_02614_));
 sky130_fd_sc_hd__a22o_1 _22474_ (.A1(net35),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net36),
    .X(_07803_));
 sky130_fd_sc_hd__a21o_1 _22475_ (.A1(net34),
    .A2(_07786_),
    .B1(_07803_),
    .X(_07804_));
 sky130_fd_sc_hd__mux2_1 _22476_ (.A0(_07804_),
    .A1(net2738),
    .S(_07794_),
    .X(_07805_));
 sky130_fd_sc_hd__clkbuf_1 _22477_ (.A(_07805_),
    .X(_02615_));
 sky130_fd_sc_hd__inv_2 _22478_ (.A(net35),
    .Y(_07806_));
 sky130_fd_sc_hd__nor2_1 _22479_ (.A(_07806_),
    .B(_07791_),
    .Y(_07807_));
 sky130_fd_sc_hd__a221o_1 _22480_ (.A1(net36),
    .A2(_07783_),
    .B1(net37),
    .B2(_07785_),
    .C1(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__mux2_1 _22481_ (.A0(_07808_),
    .A1(net2772),
    .S(_07794_),
    .X(_07809_));
 sky130_fd_sc_hd__clkbuf_1 _22482_ (.A(_07809_),
    .X(_02616_));
 sky130_fd_sc_hd__a22o_1 _22483_ (.A1(net37),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net38),
    .X(_07810_));
 sky130_fd_sc_hd__a21o_1 _22484_ (.A1(net36),
    .A2(_07786_),
    .B1(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__mux2_1 _22485_ (.A0(_07811_),
    .A1(net2731),
    .S(_07794_),
    .X(_07812_));
 sky130_fd_sc_hd__clkbuf_1 _22486_ (.A(_07812_),
    .X(_02617_));
 sky130_fd_sc_hd__a22o_1 _22487_ (.A1(net38),
    .A2(_07783_),
    .B1(_07786_),
    .B2(net37),
    .X(_07813_));
 sky130_fd_sc_hd__mux2_1 _22488_ (.A0(_07813_),
    .A1(net2757),
    .S(_07794_),
    .X(_07814_));
 sky130_fd_sc_hd__clkbuf_1 _22489_ (.A(_07814_),
    .X(_02618_));
 sky130_fd_sc_hd__inv_2 _22490_ (.A(net38),
    .Y(_07815_));
 sky130_fd_sc_hd__nor2_1 _22491_ (.A(_07815_),
    .B(_07791_),
    .Y(_07816_));
 sky130_fd_sc_hd__mux2_1 _22492_ (.A0(_07816_),
    .A1(net3881),
    .S(_07794_),
    .X(_07817_));
 sky130_fd_sc_hd__clkbuf_1 _22493_ (.A(_07817_),
    .X(_02619_));
 sky130_fd_sc_hd__mux2_1 _22494_ (.A0(net1),
    .A1(net3871),
    .S(_03834_),
    .X(_07818_));
 sky130_fd_sc_hd__clkbuf_1 _22495_ (.A(_07818_),
    .X(_02620_));
 sky130_fd_sc_hd__mux2_1 _22496_ (.A0(net2),
    .A1(net4247),
    .S(_03834_),
    .X(_07819_));
 sky130_fd_sc_hd__clkbuf_1 _22497_ (.A(_07819_),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _22498_ (.A0(net3),
    .A1(net4209),
    .S(_03834_),
    .X(_07820_));
 sky130_fd_sc_hd__clkbuf_1 _22499_ (.A(_07820_),
    .X(_02622_));
 sky130_fd_sc_hd__mux2_1 _22500_ (.A0(net4),
    .A1(net4203),
    .S(_03834_),
    .X(_07821_));
 sky130_fd_sc_hd__clkbuf_1 _22501_ (.A(_07821_),
    .X(_02623_));
 sky130_fd_sc_hd__mux2_1 _22502_ (.A0(net5),
    .A1(net4037),
    .S(_03834_),
    .X(_07822_));
 sky130_fd_sc_hd__clkbuf_1 _22503_ (.A(_07822_),
    .X(_02624_));
 sky130_fd_sc_hd__clkbuf_8 _22504_ (.A(_09222_),
    .X(_07823_));
 sky130_fd_sc_hd__mux2_1 _22505_ (.A0(net6),
    .A1(net4236),
    .S(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__clkbuf_1 _22506_ (.A(_07824_),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _22507_ (.A0(net7),
    .A1(net4205),
    .S(_07823_),
    .X(_07825_));
 sky130_fd_sc_hd__clkbuf_1 _22508_ (.A(_07825_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _22509_ (.A0(net8),
    .A1(net3917),
    .S(_07823_),
    .X(_07826_));
 sky130_fd_sc_hd__clkbuf_1 _22510_ (.A(_07826_),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _22511_ (.A0(net9),
    .A1(net4234),
    .S(_07823_),
    .X(_07827_));
 sky130_fd_sc_hd__clkbuf_1 _22512_ (.A(_07827_),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _22513_ (.A0(net10),
    .A1(net4185),
    .S(_07823_),
    .X(_07828_));
 sky130_fd_sc_hd__clkbuf_1 _22514_ (.A(_07828_),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _22515_ (.A0(net18),
    .A1(net3282),
    .S(_07823_),
    .X(_07829_));
 sky130_fd_sc_hd__clkbuf_1 _22516_ (.A(_07829_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _22517_ (.A0(net19),
    .A1(net4007),
    .S(_07823_),
    .X(_07830_));
 sky130_fd_sc_hd__clkbuf_1 _22518_ (.A(_07830_),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _22519_ (.A0(net20),
    .A1(net3508),
    .S(_07823_),
    .X(_07831_));
 sky130_fd_sc_hd__clkbuf_1 _22520_ (.A(_07831_),
    .X(_02632_));
 sky130_fd_sc_hd__mux2_1 _22521_ (.A0(net21),
    .A1(net4210),
    .S(_07823_),
    .X(_07832_));
 sky130_fd_sc_hd__clkbuf_1 _22522_ (.A(_07832_),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _22523_ (.A0(net22),
    .A1(net2812),
    .S(_07823_),
    .X(_07833_));
 sky130_fd_sc_hd__clkbuf_1 _22524_ (.A(_07833_),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _22525_ (.A0(net23),
    .A1(net3754),
    .S(_07823_),
    .X(_07834_));
 sky130_fd_sc_hd__clkbuf_1 _22526_ (.A(_07834_),
    .X(_02635_));
 sky130_fd_sc_hd__mux2_1 _22527_ (.A0(net24),
    .A1(net4062),
    .S(_07823_),
    .X(_07835_));
 sky130_fd_sc_hd__clkbuf_1 _22528_ (.A(_07835_),
    .X(_02636_));
 sky130_fd_sc_hd__mux2_1 _22529_ (.A0(net25),
    .A1(net4137),
    .S(_07823_),
    .X(_07836_));
 sky130_fd_sc_hd__clkbuf_1 _22530_ (.A(_07836_),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _22531_ (.A0(net26),
    .A1(net4219),
    .S(_07823_),
    .X(_07837_));
 sky130_fd_sc_hd__clkbuf_1 _22532_ (.A(_07837_),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_1 _22533_ (.A0(net27),
    .A1(net4048),
    .S(_07823_),
    .X(_07838_));
 sky130_fd_sc_hd__clkbuf_1 _22534_ (.A(_07838_),
    .X(_02639_));
 sky130_fd_sc_hd__mux2_1 _22535_ (.A0(net28),
    .A1(net3735),
    .S(_07823_),
    .X(_07839_));
 sky130_fd_sc_hd__clkbuf_1 _22536_ (.A(_07839_),
    .X(_02640_));
 sky130_fd_sc_hd__buf_6 _22537_ (.A(_09222_),
    .X(_07840_));
 sky130_fd_sc_hd__mux2_1 _22538_ (.A0(net29),
    .A1(net3838),
    .S(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__clkbuf_1 _22539_ (.A(_07841_),
    .X(_02641_));
 sky130_fd_sc_hd__mux2_1 _22540_ (.A0(net11),
    .A1(net2733),
    .S(_07840_),
    .X(_07842_));
 sky130_fd_sc_hd__clkbuf_1 _22541_ (.A(_07842_),
    .X(_02642_));
 sky130_fd_sc_hd__mux2_1 _22542_ (.A0(net12),
    .A1(net3281),
    .S(_07840_),
    .X(_07843_));
 sky130_fd_sc_hd__clkbuf_1 _22543_ (.A(_07843_),
    .X(_02643_));
 sky130_fd_sc_hd__mux2_1 _22544_ (.A0(net13),
    .A1(net3227),
    .S(_07840_),
    .X(_07844_));
 sky130_fd_sc_hd__clkbuf_1 _22545_ (.A(_07844_),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _22546_ (.A0(net14),
    .A1(net3783),
    .S(_07840_),
    .X(_07845_));
 sky130_fd_sc_hd__clkbuf_1 _22547_ (.A(_07845_),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _22548_ (.A0(net15),
    .A1(net4198),
    .S(_07840_),
    .X(_07846_));
 sky130_fd_sc_hd__clkbuf_1 _22549_ (.A(_07846_),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _22550_ (.A0(net16),
    .A1(net3966),
    .S(_07840_),
    .X(_07847_));
 sky130_fd_sc_hd__clkbuf_1 _22551_ (.A(_07847_),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _22552_ (.A0(net17),
    .A1(net3922),
    .S(_07840_),
    .X(_07848_));
 sky130_fd_sc_hd__clkbuf_1 _22553_ (.A(_07848_),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_1 _22554_ (.A0(net30),
    .A1(net3940),
    .S(_07840_),
    .X(_07849_));
 sky130_fd_sc_hd__clkbuf_1 _22555_ (.A(_07849_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _22556_ (.A0(net31),
    .A1(net3372),
    .S(_07840_),
    .X(_07850_));
 sky130_fd_sc_hd__clkbuf_1 _22557_ (.A(_07850_),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _22558_ (.A0(net32),
    .A1(net3911),
    .S(_07840_),
    .X(_07851_));
 sky130_fd_sc_hd__clkbuf_1 _22559_ (.A(_07851_),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _22560_ (.A0(net33),
    .A1(net4161),
    .S(_07840_),
    .X(_07852_));
 sky130_fd_sc_hd__clkbuf_1 _22561_ (.A(_07852_),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _22562_ (.A0(net34),
    .A1(net3937),
    .S(_07840_),
    .X(_07853_));
 sky130_fd_sc_hd__clkbuf_1 _22563_ (.A(_07853_),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _22564_ (.A0(net35),
    .A1(net4157),
    .S(_07840_),
    .X(_07854_));
 sky130_fd_sc_hd__clkbuf_1 _22565_ (.A(_07854_),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _22566_ (.A0(net36),
    .A1(net3822),
    .S(_07840_),
    .X(_07855_));
 sky130_fd_sc_hd__clkbuf_1 _22567_ (.A(_07855_),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _22568_ (.A0(net37),
    .A1(net4237),
    .S(_07840_),
    .X(_07856_));
 sky130_fd_sc_hd__clkbuf_1 _22569_ (.A(_07856_),
    .X(_02656_));
 sky130_fd_sc_hd__buf_8 _22570_ (.A(_09222_),
    .X(_07857_));
 sky130_fd_sc_hd__mux2_1 _22571_ (.A0(net38),
    .A1(net3942),
    .S(_07857_),
    .X(_07858_));
 sky130_fd_sc_hd__clkbuf_1 _22572_ (.A(_07858_),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _22573_ (.A0(net43),
    .A1(net2728),
    .S(_07857_),
    .X(_07859_));
 sky130_fd_sc_hd__clkbuf_1 _22574_ (.A(_07859_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _22575_ (.A0(net44),
    .A1(net3136),
    .S(_07857_),
    .X(_07860_));
 sky130_fd_sc_hd__clkbuf_1 _22576_ (.A(_07860_),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _22577_ (.A0(net45),
    .A1(net2737),
    .S(_07857_),
    .X(_07861_));
 sky130_fd_sc_hd__clkbuf_1 _22578_ (.A(_07861_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _22579_ (.A0(net46),
    .A1(net2739),
    .S(_07857_),
    .X(_07862_));
 sky130_fd_sc_hd__clkbuf_1 _22580_ (.A(_07862_),
    .X(_02661_));
 sky130_fd_sc_hd__mux2_1 _22581_ (.A0(net47),
    .A1(net3206),
    .S(_07857_),
    .X(_07863_));
 sky130_fd_sc_hd__clkbuf_1 _22582_ (.A(_07863_),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _22583_ (.A0(net48),
    .A1(net4067),
    .S(_07857_),
    .X(_07864_));
 sky130_fd_sc_hd__clkbuf_1 _22584_ (.A(_07864_),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _22585_ (.A0(net39),
    .A1(net2732),
    .S(_07857_),
    .X(_07865_));
 sky130_fd_sc_hd__clkbuf_1 _22586_ (.A(_07865_),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _22587_ (.A0(net40),
    .A1(net3326),
    .S(_07857_),
    .X(_07866_));
 sky130_fd_sc_hd__clkbuf_1 _22588_ (.A(_07866_),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_1 _22589_ (.A0(net41),
    .A1(net4188),
    .S(_07857_),
    .X(_07867_));
 sky130_fd_sc_hd__clkbuf_1 _22590_ (.A(_07867_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _22591_ (.A0(net42),
    .A1(net3743),
    .S(_07857_),
    .X(_07868_));
 sky130_fd_sc_hd__clkbuf_1 _22592_ (.A(_07868_),
    .X(_02667_));
 sky130_fd_sc_hd__a22o_1 _22593_ (.A1(net3),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net4),
    .X(_07869_));
 sky130_fd_sc_hd__a21o_1 _22594_ (.A1(net2),
    .A2(_07786_),
    .B1(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__mux2_1 _22595_ (.A0(_07870_),
    .A1(net4026),
    .S(_07794_),
    .X(_07871_));
 sky130_fd_sc_hd__clkbuf_1 _22596_ (.A(_07871_),
    .X(_02668_));
 sky130_fd_sc_hd__a22o_1 _22597_ (.A1(net4),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net5),
    .X(_07872_));
 sky130_fd_sc_hd__a21o_1 _22598_ (.A1(net3),
    .A2(_07786_),
    .B1(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__mux2_1 _22599_ (.A0(_07873_),
    .A1(net3923),
    .S(_07794_),
    .X(_07874_));
 sky130_fd_sc_hd__clkbuf_1 _22600_ (.A(_07874_),
    .X(_02669_));
 sky130_fd_sc_hd__a22o_1 _22601_ (.A1(net5),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net6),
    .X(_07875_));
 sky130_fd_sc_hd__a21o_1 _22602_ (.A1(net4),
    .A2(_07786_),
    .B1(_07875_),
    .X(_07876_));
 sky130_fd_sc_hd__mux2_1 _22603_ (.A0(_07876_),
    .A1(net4086),
    .S(_07794_),
    .X(_07877_));
 sky130_fd_sc_hd__clkbuf_1 _22604_ (.A(_07877_),
    .X(_02670_));
 sky130_fd_sc_hd__a22o_1 _22605_ (.A1(net6),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net7),
    .X(_07878_));
 sky130_fd_sc_hd__a21o_1 _22606_ (.A1(net5),
    .A2(_07786_),
    .B1(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__mux2_1 _22607_ (.A0(_07879_),
    .A1(net3898),
    .S(_07794_),
    .X(_07880_));
 sky130_fd_sc_hd__clkbuf_1 _22608_ (.A(_07880_),
    .X(_02671_));
 sky130_fd_sc_hd__a22o_1 _22609_ (.A1(net7),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net8),
    .X(_07881_));
 sky130_fd_sc_hd__a21o_1 _22610_ (.A1(net6),
    .A2(_07786_),
    .B1(_07881_),
    .X(_07882_));
 sky130_fd_sc_hd__mux2_1 _22611_ (.A0(_07882_),
    .A1(net4287),
    .S(_07794_),
    .X(_07883_));
 sky130_fd_sc_hd__clkbuf_1 _22612_ (.A(_07883_),
    .X(_02672_));
 sky130_fd_sc_hd__a22o_1 _22613_ (.A1(net8),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net9),
    .X(_07884_));
 sky130_fd_sc_hd__a21o_1 _22614_ (.A1(net7),
    .A2(_07786_),
    .B1(_07884_),
    .X(_07885_));
 sky130_fd_sc_hd__mux2_1 _22615_ (.A0(_07885_),
    .A1(net4124),
    .S(_07794_),
    .X(_07886_));
 sky130_fd_sc_hd__clkbuf_1 _22616_ (.A(_07886_),
    .X(_02673_));
 sky130_fd_sc_hd__a22o_1 _22617_ (.A1(net9),
    .A2(_07783_),
    .B1(_07785_),
    .B2(net10),
    .X(_07887_));
 sky130_fd_sc_hd__a21o_1 _22618_ (.A1(net8),
    .A2(_07786_),
    .B1(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__mux2_1 _22619_ (.A0(_07888_),
    .A1(net4145),
    .S(_07794_),
    .X(_07889_));
 sky130_fd_sc_hd__clkbuf_1 _22620_ (.A(_07889_),
    .X(_02674_));
 sky130_fd_sc_hd__a22o_1 _22621_ (.A1(net10),
    .A2(_07783_),
    .B1(_07786_),
    .B2(net9),
    .X(_07890_));
 sky130_fd_sc_hd__mux2_1 _22622_ (.A0(_07890_),
    .A1(net4063),
    .S(_07794_),
    .X(_07891_));
 sky130_fd_sc_hd__clkbuf_1 _22623_ (.A(_07891_),
    .X(_02675_));
 sky130_fd_sc_hd__and2_1 _22624_ (.A(_07786_),
    .B(net10),
    .X(_07892_));
 sky130_fd_sc_hd__mux2_1 _22625_ (.A0(_07892_),
    .A1(net2712),
    .S(_07793_),
    .X(_07893_));
 sky130_fd_sc_hd__clkbuf_1 _22626_ (.A(_07893_),
    .X(_02676_));
 sky130_fd_sc_hd__inv_2 _22627_ (.A(\base_h_bporch[6] ),
    .Y(_07894_));
 sky130_fd_sc_hd__nand2_1 _22628_ (.A(_08966_),
    .B(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand3_2 _22629_ (.A(_08926_),
    .B(\base_h_bporch[6] ),
    .C(_08965_),
    .Y(_07896_));
 sky130_fd_sc_hd__nand2_1 _22630_ (.A(_07895_),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__nor2_1 _22631_ (.A(_08928_),
    .B(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__inv_2 _22632_ (.A(\base_h_bporch[1] ),
    .Y(_07899_));
 sky130_fd_sc_hd__nand2_1 _22633_ (.A(_08951_),
    .B(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__nand3_1 _22634_ (.A(_08880_),
    .B(_08950_),
    .C(\base_h_bporch[1] ),
    .Y(_07901_));
 sky130_fd_sc_hd__nand2_1 _22635_ (.A(_08955_),
    .B(\base_h_bporch[0] ),
    .Y(_07902_));
 sky130_fd_sc_hd__inv_2 _22636_ (.A(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand3_1 _22637_ (.A(_07900_),
    .B(_07901_),
    .C(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__nand2_1 _22638_ (.A(_07904_),
    .B(_07901_),
    .Y(_07905_));
 sky130_fd_sc_hd__nand3_2 _22639_ (.A(_08890_),
    .B(_08942_),
    .C(\base_h_bporch[2] ),
    .Y(_07906_));
 sky130_fd_sc_hd__inv_2 _22640_ (.A(\base_h_bporch[2] ),
    .Y(_07907_));
 sky130_fd_sc_hd__nand2_1 _22641_ (.A(_08943_),
    .B(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__nand3_1 _22642_ (.A(_07905_),
    .B(_07906_),
    .C(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__nand2_1 _22643_ (.A(_07909_),
    .B(_07906_),
    .Y(_07910_));
 sky130_fd_sc_hd__inv_2 _22644_ (.A(\base_h_bporch[3] ),
    .Y(_07911_));
 sky130_fd_sc_hd__nand2_1 _22645_ (.A(_08947_),
    .B(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__nand2_1 _22646_ (.A(_07910_),
    .B(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__or2_1 _22647_ (.A(_07911_),
    .B(_08947_),
    .X(_07914_));
 sky130_fd_sc_hd__nand2_1 _22648_ (.A(_07913_),
    .B(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__inv_2 _22649_ (.A(\base_h_bporch[5] ),
    .Y(_07916_));
 sky130_fd_sc_hd__nand2_1 _22650_ (.A(_08936_),
    .B(_07916_),
    .Y(_07917_));
 sky130_fd_sc_hd__nand3_2 _22651_ (.A(_08933_),
    .B(_08935_),
    .C(\base_h_bporch[5] ),
    .Y(_07918_));
 sky130_fd_sc_hd__inv_2 _22652_ (.A(\base_h_bporch[4] ),
    .Y(_07919_));
 sky130_fd_sc_hd__nand2_1 _22653_ (.A(_08938_),
    .B(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__nand3_2 _22654_ (.A(_08931_),
    .B(_08937_),
    .C(\base_h_bporch[4] ),
    .Y(_07921_));
 sky130_fd_sc_hd__nand2_1 _22655_ (.A(_07920_),
    .B(_07921_),
    .Y(_07922_));
 sky130_fd_sc_hd__inv_2 _22656_ (.A(_07922_),
    .Y(_07923_));
 sky130_fd_sc_hd__nand3_1 _22657_ (.A(_07917_),
    .B(_07918_),
    .C(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__inv_2 _22658_ (.A(_07924_),
    .Y(_07925_));
 sky130_fd_sc_hd__nand3_1 _22659_ (.A(_07898_),
    .B(_07915_),
    .C(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__nor2_1 _22660_ (.A(_07896_),
    .B(_08928_),
    .Y(_07927_));
 sky130_fd_sc_hd__inv_2 _22661_ (.A(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__clkinvlp_2 _22662_ (.A(_07921_),
    .Y(_07929_));
 sky130_fd_sc_hd__nand3_1 _22663_ (.A(_07917_),
    .B(_07918_),
    .C(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__nand2_1 _22664_ (.A(_07930_),
    .B(_07918_),
    .Y(_07931_));
 sky130_fd_sc_hd__nand2_1 _22665_ (.A(_07898_),
    .B(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__nand3_1 _22666_ (.A(_07926_),
    .B(_07928_),
    .C(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__nand2_1 _22667_ (.A(_07933_),
    .B(_08916_),
    .Y(_07934_));
 sky130_fd_sc_hd__nand2_1 _22668_ (.A(_07934_),
    .B(_08919_),
    .Y(_07935_));
 sky130_fd_sc_hd__nand3_1 _22669_ (.A(_07933_),
    .B(_08920_),
    .C(_08916_),
    .Y(_07936_));
 sky130_fd_sc_hd__nand2_1 _22670_ (.A(_07935_),
    .B(_07936_),
    .Y(_07937_));
 sky130_fd_sc_hd__nand2_1 _22671_ (.A(_07923_),
    .B(_07915_),
    .Y(_07938_));
 sky130_fd_sc_hd__nand2_1 _22672_ (.A(_07938_),
    .B(_07921_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_1 _22673_ (.A(_08936_),
    .B(\base_h_bporch[5] ),
    .Y(_07940_));
 sky130_fd_sc_hd__nand3_1 _22674_ (.A(_08933_),
    .B(_08935_),
    .C(_07916_),
    .Y(_07941_));
 sky130_fd_sc_hd__nand2_1 _22675_ (.A(_07940_),
    .B(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__nand2_1 _22676_ (.A(_07939_),
    .B(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_1 _22677_ (.A(_07943_),
    .B(_07918_),
    .Y(_07944_));
 sky130_fd_sc_hd__clkinvlp_2 _22678_ (.A(_07897_),
    .Y(_07945_));
 sky130_fd_sc_hd__nand2_1 _22679_ (.A(_07944_),
    .B(_07945_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand3_1 _22680_ (.A(_07943_),
    .B(_07918_),
    .C(_07897_),
    .Y(_07947_));
 sky130_fd_sc_hd__nand2_1 _22681_ (.A(_07946_),
    .B(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__nand2_1 _22682_ (.A(_07917_),
    .B(_07918_),
    .Y(_07949_));
 sky130_fd_sc_hd__nand3_1 _22683_ (.A(_07949_),
    .B(_07921_),
    .C(_07938_),
    .Y(_07950_));
 sky130_fd_sc_hd__nand2_1 _22684_ (.A(_07950_),
    .B(_07943_),
    .Y(_07951_));
 sky130_fd_sc_hd__nand3_1 _22685_ (.A(_07922_),
    .B(_07914_),
    .C(_07913_),
    .Y(_07952_));
 sky130_fd_sc_hd__nand2_1 _22686_ (.A(_07952_),
    .B(_07938_),
    .Y(_07953_));
 sky130_fd_sc_hd__a21boi_1 _22687_ (.A1(_07905_),
    .A2(_07908_),
    .B1_N(_07906_),
    .Y(_07954_));
 sky130_fd_sc_hd__nand3_1 _22688_ (.A(_08944_),
    .B(_08946_),
    .C(_07911_),
    .Y(_07955_));
 sky130_fd_sc_hd__nand2_1 _22689_ (.A(_08947_),
    .B(\base_h_bporch[3] ),
    .Y(_07956_));
 sky130_fd_sc_hd__nand3_1 _22690_ (.A(_07954_),
    .B(_07955_),
    .C(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__nand2_1 _22691_ (.A(_07956_),
    .B(_07955_),
    .Y(_07958_));
 sky130_fd_sc_hd__nand2_1 _22692_ (.A(_07958_),
    .B(_07910_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_1 _22693_ (.A(_07957_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__inv_2 _22694_ (.A(_07905_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand2_1 _22695_ (.A(_07908_),
    .B(_07906_),
    .Y(_07962_));
 sky130_fd_sc_hd__nand2_1 _22696_ (.A(_07961_),
    .B(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__nand2_1 _22697_ (.A(_07909_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__nand2_1 _22698_ (.A(_07900_),
    .B(_07901_),
    .Y(_07965_));
 sky130_fd_sc_hd__nand2_1 _22699_ (.A(_07965_),
    .B(_07902_),
    .Y(_07966_));
 sky130_fd_sc_hd__nand2_1 _22700_ (.A(_07966_),
    .B(_07904_),
    .Y(_07967_));
 sky130_fd_sc_hd__or2_1 _22701_ (.A(\base_h_bporch[0] ),
    .B(_08955_),
    .X(_07968_));
 sky130_fd_sc_hd__nand2_1 _22702_ (.A(_07968_),
    .B(_07902_),
    .Y(_07969_));
 sky130_fd_sc_hd__nand2_1 _22703_ (.A(_07967_),
    .B(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__inv_2 _22704_ (.A(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__nand2_1 _22705_ (.A(_07964_),
    .B(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__inv_2 _22706_ (.A(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__nand2_1 _22707_ (.A(_07960_),
    .B(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__inv_2 _22708_ (.A(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__nand2_1 _22709_ (.A(_07953_),
    .B(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__inv_2 _22710_ (.A(_07976_),
    .Y(_07977_));
 sky130_fd_sc_hd__nand2_2 _22711_ (.A(_07951_),
    .B(_07977_),
    .Y(_07978_));
 sky130_fd_sc_hd__inv_2 _22712_ (.A(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__nand2_1 _22713_ (.A(_07948_),
    .B(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__nand2_1 _22714_ (.A(_07946_),
    .B(_07896_),
    .Y(_07981_));
 sky130_fd_sc_hd__nand2_1 _22715_ (.A(_07981_),
    .B(_08928_),
    .Y(_07982_));
 sky130_fd_sc_hd__nand3_1 _22716_ (.A(_07946_),
    .B(_08929_),
    .C(_07896_),
    .Y(_07983_));
 sky130_fd_sc_hd__nand2_1 _22717_ (.A(_07982_),
    .B(_07983_),
    .Y(_07984_));
 sky130_fd_sc_hd__nor2_1 _22718_ (.A(_07980_),
    .B(_07984_),
    .Y(_07985_));
 sky130_fd_sc_hd__a21oi_1 _22719_ (.A1(_07898_),
    .A2(_07931_),
    .B1(_07927_),
    .Y(_07986_));
 sky130_fd_sc_hd__nand3_1 _22720_ (.A(_07986_),
    .B(_08915_),
    .C(_07926_),
    .Y(_07987_));
 sky130_fd_sc_hd__nand2_1 _22721_ (.A(_07934_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__nand3_1 _22722_ (.A(_07937_),
    .B(_07985_),
    .C(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__inv_2 _22723_ (.A(_07980_),
    .Y(_07990_));
 sky130_fd_sc_hd__nand2_1 _22724_ (.A(_07984_),
    .B(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__nand2_1 _22725_ (.A(_07981_),
    .B(_08929_),
    .Y(_07992_));
 sky130_fd_sc_hd__nand3_1 _22726_ (.A(_07946_),
    .B(_08928_),
    .C(_07896_),
    .Y(_07993_));
 sky130_fd_sc_hd__nand2_1 _22727_ (.A(_07992_),
    .B(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__nand2_1 _22728_ (.A(_07994_),
    .B(_07980_),
    .Y(_07995_));
 sky130_fd_sc_hd__nand2_1 _22729_ (.A(_07991_),
    .B(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_1 _22730_ (.A(_07996_),
    .B(net3443),
    .Y(_07997_));
 sky130_fd_sc_hd__nand2_1 _22731_ (.A(_07989_),
    .B(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__nand3_1 _22732_ (.A(_07991_),
    .B(_07995_),
    .C(_08512_),
    .Y(_07999_));
 sky130_fd_sc_hd__nand3_1 _22733_ (.A(_07974_),
    .B(_07952_),
    .C(_07938_),
    .Y(_08000_));
 sky130_fd_sc_hd__a21oi_1 _22734_ (.A1(_07976_),
    .A2(_08000_),
    .B1(\base_h_counter[4] ),
    .Y(_08001_));
 sky130_fd_sc_hd__nand3_1 _22735_ (.A(_07957_),
    .B(_07959_),
    .C(_07972_),
    .Y(_08002_));
 sky130_fd_sc_hd__a21oi_1 _22736_ (.A1(_07974_),
    .A2(_08002_),
    .B1(\base_h_counter[3] ),
    .Y(_08003_));
 sky130_fd_sc_hd__nand3_1 _22737_ (.A(_07909_),
    .B(_07963_),
    .C(_07970_),
    .Y(_08004_));
 sky130_fd_sc_hd__a21oi_1 _22738_ (.A1(_07972_),
    .A2(_08004_),
    .B1(\base_h_counter[2] ),
    .Y(_08005_));
 sky130_fd_sc_hd__nand3_1 _22739_ (.A(_07972_),
    .B(_08004_),
    .C(\base_h_counter[2] ),
    .Y(_08006_));
 sky130_fd_sc_hd__nand3_1 _22740_ (.A(_07966_),
    .B(_07904_),
    .C(_07969_),
    .Y(_08007_));
 sky130_fd_sc_hd__nand3_1 _22741_ (.A(_07965_),
    .B(_07902_),
    .C(_07968_),
    .Y(_08008_));
 sky130_fd_sc_hd__nand2_1 _22742_ (.A(_08007_),
    .B(_08008_),
    .Y(_08009_));
 sky130_fd_sc_hd__nand2_1 _22743_ (.A(_08009_),
    .B(_08526_),
    .Y(_08010_));
 sky130_fd_sc_hd__xor2_1 _22744_ (.A(_08525_),
    .B(_07969_),
    .X(_08011_));
 sky130_fd_sc_hd__nand3_1 _22745_ (.A(_08007_),
    .B(_08527_),
    .C(_08008_),
    .Y(_08012_));
 sky130_fd_sc_hd__nand3_1 _22746_ (.A(_08010_),
    .B(_08011_),
    .C(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__inv_2 _22747_ (.A(_08013_),
    .Y(_08014_));
 sky130_fd_sc_hd__nand2_1 _22748_ (.A(_08006_),
    .B(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__nor2_1 _22749_ (.A(_08005_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand3_1 _22750_ (.A(_07974_),
    .B(_08002_),
    .C(\base_h_counter[3] ),
    .Y(_08017_));
 sky130_fd_sc_hd__nand2_1 _22751_ (.A(_08016_),
    .B(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__nor2_1 _22752_ (.A(_08003_),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand3_1 _22753_ (.A(_07976_),
    .B(_08000_),
    .C(\base_h_counter[4] ),
    .Y(_08020_));
 sky130_fd_sc_hd__nand2_1 _22754_ (.A(_08019_),
    .B(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__nor2_1 _22755_ (.A(_08001_),
    .B(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__nand3_1 _22756_ (.A(_07976_),
    .B(_07950_),
    .C(_07943_),
    .Y(_08023_));
 sky130_fd_sc_hd__nand2_1 _22757_ (.A(_07978_),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__nand2_1 _22758_ (.A(_08024_),
    .B(_08519_),
    .Y(_08025_));
 sky130_fd_sc_hd__nand3_1 _22759_ (.A(_07978_),
    .B(_08023_),
    .C(\base_h_counter[5] ),
    .Y(_08026_));
 sky130_fd_sc_hd__nand3_1 _22760_ (.A(_08022_),
    .B(_08025_),
    .C(_08026_),
    .Y(_08027_));
 sky130_fd_sc_hd__nand3_1 _22761_ (.A(_07978_),
    .B(_07946_),
    .C(_07947_),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_1 _22762_ (.A(_07980_),
    .B(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__nor2_1 _22763_ (.A(_08509_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__nor2_1 _22764_ (.A(_08027_),
    .B(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__nand2_1 _22765_ (.A(_08029_),
    .B(_08509_),
    .Y(_08032_));
 sky130_fd_sc_hd__nand3_1 _22766_ (.A(_07999_),
    .B(_08031_),
    .C(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__nor2_1 _22767_ (.A(_07998_),
    .B(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand2_1 _22768_ (.A(_07985_),
    .B(_07988_),
    .Y(_08035_));
 sky130_fd_sc_hd__inv_2 _22769_ (.A(_07988_),
    .Y(_08036_));
 sky130_fd_sc_hd__nand2_1 _22770_ (.A(_07994_),
    .B(_07990_),
    .Y(_08037_));
 sky130_fd_sc_hd__nand2_1 _22771_ (.A(_08036_),
    .B(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__nand3_1 _22772_ (.A(_08035_),
    .B(_08038_),
    .C(net4150),
    .Y(_08039_));
 sky130_fd_sc_hd__nand2_1 _22773_ (.A(_07985_),
    .B(_08036_),
    .Y(_08040_));
 sky130_fd_sc_hd__nand2_1 _22774_ (.A(_08037_),
    .B(_07988_),
    .Y(_08041_));
 sky130_fd_sc_hd__nand3_1 _22775_ (.A(_08040_),
    .B(_08554_),
    .C(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__nand2_1 _22776_ (.A(_08039_),
    .B(_08042_),
    .Y(_08043_));
 sky130_fd_sc_hd__inv_2 _22777_ (.A(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__inv_2 _22778_ (.A(_07937_),
    .Y(_08045_));
 sky130_fd_sc_hd__nand2_1 _22779_ (.A(_08035_),
    .B(_08045_),
    .Y(_08046_));
 sky130_fd_sc_hd__nand2_1 _22780_ (.A(_08046_),
    .B(_08921_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand3_1 _22781_ (.A(_08035_),
    .B(_08045_),
    .C(net2896),
    .Y(_08048_));
 sky130_fd_sc_hd__nand2_1 _22782_ (.A(_08047_),
    .B(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__nand3_4 _22783_ (.A(_08034_),
    .B(_08044_),
    .C(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__nor2_4 _22784_ (.A(_08722_),
    .B(net4316),
    .Y(_08051_));
 sky130_fd_sc_hd__nand2_4 _22785_ (.A(_08050_),
    .B(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__inv_6 _22786_ (.A(_08052_),
    .Y(_08053_));
 sky130_fd_sc_hd__mux2_1 _22787_ (.A0(_08053_),
    .A1(_08793_),
    .S(net4319),
    .X(_08054_));
 sky130_fd_sc_hd__clkbuf_1 _22788_ (.A(_08054_),
    .X(_02677_));
 sky130_fd_sc_hd__nor2_1 _22789_ (.A(_08526_),
    .B(\base_h_counter[0] ),
    .Y(_08055_));
 sky130_fd_sc_hd__nand2_1 _22790_ (.A(_08526_),
    .B(net4319),
    .Y(_08056_));
 sky130_fd_sc_hd__inv_2 _22791_ (.A(_08056_),
    .Y(_08057_));
 sky130_fd_sc_hd__nor2_1 _22792_ (.A(_08055_),
    .B(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__a22o_1 _22793_ (.A1(_08526_),
    .A2(_08793_),
    .B1(_08053_),
    .B2(_08058_),
    .X(_02678_));
 sky130_fd_sc_hd__xor2_1 _22794_ (.A(net4320),
    .B(_08056_),
    .X(_08059_));
 sky130_fd_sc_hd__o22ai_1 _22795_ (.A1(_08535_),
    .A2(_04971_),
    .B1(_08059_),
    .B2(_08052_),
    .Y(_02679_));
 sky130_fd_sc_hd__and3_1 _22796_ (.A(_08057_),
    .B(net4323),
    .C(net4320),
    .X(_08060_));
 sky130_fd_sc_hd__inv_2 _22797_ (.A(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__o21ai_1 _22798_ (.A1(_08535_),
    .A2(_08056_),
    .B1(_08524_),
    .Y(_08062_));
 sky130_fd_sc_hd__nand2_1 _22799_ (.A(_08061_),
    .B(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__o22ai_1 _22800_ (.A1(_08524_),
    .A2(_04971_),
    .B1(_08063_),
    .B2(_08052_),
    .Y(_02680_));
 sky130_fd_sc_hd__nor2_1 _22801_ (.A(net3660),
    .B(_08060_),
    .Y(_08064_));
 sky130_fd_sc_hd__nor2_1 _22802_ (.A(_08522_),
    .B(_08061_),
    .Y(_08065_));
 sky130_fd_sc_hd__nor2_1 _22803_ (.A(_08064_),
    .B(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__a22o_1 _22804_ (.A1(net3660),
    .A2(_08793_),
    .B1(_08053_),
    .B2(_08066_),
    .X(_02681_));
 sky130_fd_sc_hd__or2_1 _22805_ (.A(net4327),
    .B(_08065_),
    .X(_08067_));
 sky130_fd_sc_hd__nand2_1 _22806_ (.A(_08065_),
    .B(net4327),
    .Y(_08068_));
 sky130_fd_sc_hd__nand2_1 _22807_ (.A(_08067_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__o22ai_1 _22808_ (.A1(_08519_),
    .A2(_04971_),
    .B1(_08069_),
    .B2(_08052_),
    .Y(_02682_));
 sky130_fd_sc_hd__or2_1 _22809_ (.A(_08509_),
    .B(_08068_),
    .X(_08070_));
 sky130_fd_sc_hd__nand2_1 _22810_ (.A(_08068_),
    .B(_08509_),
    .Y(_08071_));
 sky130_fd_sc_hd__nand2_1 _22811_ (.A(_08070_),
    .B(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__o22ai_1 _22812_ (.A1(_08509_),
    .A2(_04971_),
    .B1(_08072_),
    .B2(_08052_),
    .Y(_02683_));
 sky130_fd_sc_hd__nor2_1 _22813_ (.A(_08512_),
    .B(_08070_),
    .Y(_08073_));
 sky130_fd_sc_hd__nand2_1 _22814_ (.A(_08070_),
    .B(_08512_),
    .Y(_08074_));
 sky130_fd_sc_hd__and2b_1 _22815_ (.A_N(_08073_),
    .B(_08074_),
    .X(_08075_));
 sky130_fd_sc_hd__a22o_1 _22816_ (.A1(net3443),
    .A2(_08793_),
    .B1(_08053_),
    .B2(_08075_),
    .X(_02684_));
 sky130_fd_sc_hd__or2_1 _22817_ (.A(net4150),
    .B(_08073_),
    .X(_08076_));
 sky130_fd_sc_hd__nand2_1 _22818_ (.A(_08073_),
    .B(net4150),
    .Y(_08077_));
 sky130_fd_sc_hd__nand2_1 _22819_ (.A(_08076_),
    .B(net4151),
    .Y(_08078_));
 sky130_fd_sc_hd__o22ai_1 _22820_ (.A1(_08554_),
    .A2(_04971_),
    .B1(_08078_),
    .B2(_08052_),
    .Y(_02685_));
 sky130_fd_sc_hd__xor2_1 _22821_ (.A(_08921_),
    .B(_08077_),
    .X(_08079_));
 sky130_fd_sc_hd__a22o_1 _22822_ (.A1(net2896),
    .A2(_08793_),
    .B1(_08053_),
    .B2(_08079_),
    .X(_02686_));
 sky130_fd_sc_hd__nor2_2 _22823_ (.A(_08793_),
    .B(_08053_),
    .Y(_08080_));
 sky130_fd_sc_hd__buf_6 _22824_ (.A(_08080_),
    .X(_08081_));
 sky130_fd_sc_hd__inv_2 _22825_ (.A(\base_v_bporch[2] ),
    .Y(_08082_));
 sky130_fd_sc_hd__nand2_1 _22826_ (.A(_09143_),
    .B(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__nand3_2 _22827_ (.A(_09142_),
    .B(\base_v_bporch[2] ),
    .C(_09091_),
    .Y(_08084_));
 sky130_fd_sc_hd__nand2_1 _22828_ (.A(_09132_),
    .B(\base_v_bporch[0] ),
    .Y(_08085_));
 sky130_fd_sc_hd__inv_2 _22829_ (.A(\base_v_bporch[1] ),
    .Y(_08086_));
 sky130_fd_sc_hd__nand2_1 _22830_ (.A(_09135_),
    .B(_08086_),
    .Y(_08087_));
 sky130_fd_sc_hd__nand3_2 _22831_ (.A(_09134_),
    .B(\base_v_bporch[1] ),
    .C(_09086_),
    .Y(_08088_));
 sky130_fd_sc_hd__nand3b_1 _22832_ (.A_N(_08085_),
    .B(_08087_),
    .C(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__nand2_1 _22833_ (.A(_08089_),
    .B(_08088_),
    .Y(_08090_));
 sky130_fd_sc_hd__nand3_2 _22834_ (.A(_08083_),
    .B(_08084_),
    .C(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand2_1 _22835_ (.A(_08091_),
    .B(_08084_),
    .Y(_08092_));
 sky130_fd_sc_hd__nand3_2 _22836_ (.A(_09093_),
    .B(_09139_),
    .C(\base_v_bporch[3] ),
    .Y(_08093_));
 sky130_fd_sc_hd__a21o_1 _22837_ (.A1(_09093_),
    .A2(_09139_),
    .B1(\base_v_bporch[3] ),
    .X(_08094_));
 sky130_fd_sc_hd__nand3_2 _22838_ (.A(_08092_),
    .B(_08093_),
    .C(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__nand2_1 _22839_ (.A(_08095_),
    .B(_08093_),
    .Y(_08096_));
 sky130_fd_sc_hd__nand3_1 _22840_ (.A(_09094_),
    .B(_09013_),
    .C(_09095_),
    .Y(_08097_));
 sky130_fd_sc_hd__inv_2 _22841_ (.A(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__nand3b_1 _22842_ (.A_N(_09115_),
    .B(_08096_),
    .C(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand2_1 _22843_ (.A(_08099_),
    .B(_09112_),
    .Y(_08100_));
 sky130_fd_sc_hd__nand3_1 _22844_ (.A(_09109_),
    .B(_09069_),
    .C(_09114_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand3b_1 _22845_ (.A_N(_08101_),
    .B(_08096_),
    .C(_08098_),
    .Y(_08102_));
 sky130_fd_sc_hd__nand2_1 _22846_ (.A(_08100_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__inv_2 _22847_ (.A(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__nand2_1 _22848_ (.A(_08096_),
    .B(_09097_),
    .Y(_08105_));
 sky130_fd_sc_hd__nand3_1 _22849_ (.A(_08095_),
    .B(_09096_),
    .C(_08093_),
    .Y(_08106_));
 sky130_fd_sc_hd__nand2_1 _22850_ (.A(_08094_),
    .B(_08093_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand3_1 _22851_ (.A(_08107_),
    .B(_08091_),
    .C(_08084_),
    .Y(_08108_));
 sky130_fd_sc_hd__nand2_1 _22852_ (.A(_08108_),
    .B(_08095_),
    .Y(_08109_));
 sky130_fd_sc_hd__nand2_1 _22853_ (.A(_08083_),
    .B(_08084_),
    .Y(_08110_));
 sky130_fd_sc_hd__nand3_1 _22854_ (.A(_08110_),
    .B(_08088_),
    .C(_08089_),
    .Y(_08111_));
 sky130_fd_sc_hd__nand2_1 _22855_ (.A(_08111_),
    .B(_08091_),
    .Y(_08112_));
 sky130_fd_sc_hd__nand2_1 _22856_ (.A(_08087_),
    .B(_08088_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand2_1 _22857_ (.A(_08113_),
    .B(_08085_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_1 _22858_ (.A(_08114_),
    .B(_08089_),
    .Y(_08115_));
 sky130_fd_sc_hd__or2_1 _22859_ (.A(\base_v_bporch[0] ),
    .B(_09132_),
    .X(_08116_));
 sky130_fd_sc_hd__nand2_1 _22860_ (.A(_08116_),
    .B(_08085_),
    .Y(_08117_));
 sky130_fd_sc_hd__nand2_1 _22861_ (.A(_08115_),
    .B(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__inv_2 _22862_ (.A(_08118_),
    .Y(_08119_));
 sky130_fd_sc_hd__nand2_1 _22863_ (.A(_08112_),
    .B(_08119_),
    .Y(_08120_));
 sky130_fd_sc_hd__inv_2 _22864_ (.A(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__nand2_1 _22865_ (.A(_08109_),
    .B(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__a21oi_2 _22866_ (.A1(_08105_),
    .A2(_08106_),
    .B1(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__nand2_1 _22867_ (.A(_08105_),
    .B(_09103_),
    .Y(_08124_));
 sky130_fd_sc_hd__nand2_1 _22868_ (.A(_08096_),
    .B(_08098_),
    .Y(_08125_));
 sky130_fd_sc_hd__nand2_2 _22869_ (.A(_08124_),
    .B(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__nand2_1 _22870_ (.A(_08125_),
    .B(_09115_),
    .Y(_08127_));
 sky130_fd_sc_hd__nand2_1 _22871_ (.A(_08127_),
    .B(_08099_),
    .Y(_08128_));
 sky130_fd_sc_hd__nand3_1 _22872_ (.A(_08123_),
    .B(_08126_),
    .C(_08128_),
    .Y(_08129_));
 sky130_fd_sc_hd__nor2_1 _22873_ (.A(_08104_),
    .B(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__inv_2 _22874_ (.A(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__nand2_1 _22875_ (.A(_08129_),
    .B(_08104_),
    .Y(_08132_));
 sky130_fd_sc_hd__nand2_1 _22876_ (.A(_08131_),
    .B(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__nand2_1 _22877_ (.A(_08133_),
    .B(_08565_),
    .Y(_08134_));
 sky130_fd_sc_hd__nand3_1 _22878_ (.A(_08131_),
    .B(\base_v_counter[7] ),
    .C(_08132_),
    .Y(_08135_));
 sky130_fd_sc_hd__or2_1 _22879_ (.A(_09125_),
    .B(_08102_),
    .X(_08136_));
 sky130_fd_sc_hd__nand2_1 _22880_ (.A(_08136_),
    .B(_09159_),
    .Y(_08137_));
 sky130_fd_sc_hd__or2_1 _22881_ (.A(_08606_),
    .B(_08137_),
    .X(_08138_));
 sky130_fd_sc_hd__nand3_1 _22882_ (.A(_08134_),
    .B(_08135_),
    .C(_08138_),
    .Y(_08139_));
 sky130_fd_sc_hd__nand2_1 _22883_ (.A(_08123_),
    .B(_08126_),
    .Y(_08140_));
 sky130_fd_sc_hd__nand2_1 _22884_ (.A(_08140_),
    .B(_08128_),
    .Y(_08141_));
 sky130_fd_sc_hd__inv_2 _22885_ (.A(_08128_),
    .Y(_08142_));
 sky130_fd_sc_hd__nand3_1 _22886_ (.A(_08142_),
    .B(_08123_),
    .C(_08126_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand3_1 _22887_ (.A(_08141_),
    .B(_08143_),
    .C(_08562_),
    .Y(_08144_));
 sky130_fd_sc_hd__nand2_1 _22888_ (.A(_08140_),
    .B(_08142_),
    .Y(_08145_));
 sky130_fd_sc_hd__nand3_1 _22889_ (.A(_08145_),
    .B(\base_v_counter[6] ),
    .C(_08129_),
    .Y(_08146_));
 sky130_fd_sc_hd__nand2_1 _22890_ (.A(_08144_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__nand2_1 _22891_ (.A(_08105_),
    .B(_08106_),
    .Y(_08148_));
 sky130_fd_sc_hd__nand2b_1 _22892_ (.A_N(_08148_),
    .B(_08122_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand3_1 _22893_ (.A(_08148_),
    .B(_08121_),
    .C(_08109_),
    .Y(_08150_));
 sky130_fd_sc_hd__nand2_1 _22894_ (.A(_08149_),
    .B(_08150_),
    .Y(_08151_));
 sky130_fd_sc_hd__nand2_1 _22895_ (.A(_08151_),
    .B(_08577_),
    .Y(_08152_));
 sky130_fd_sc_hd__nand3_1 _22896_ (.A(_08120_),
    .B(_08108_),
    .C(_08095_),
    .Y(_08153_));
 sky130_fd_sc_hd__a21oi_1 _22897_ (.A1(_08122_),
    .A2(_08153_),
    .B1(\base_v_counter[3] ),
    .Y(_08154_));
 sky130_fd_sc_hd__nand3_1 _22898_ (.A(_08111_),
    .B(_08091_),
    .C(_08118_),
    .Y(_08155_));
 sky130_fd_sc_hd__a21oi_1 _22899_ (.A1(_08120_),
    .A2(_08155_),
    .B1(\base_v_counter[2] ),
    .Y(_08156_));
 sky130_fd_sc_hd__nand3_1 _22900_ (.A(_08120_),
    .B(\base_v_counter[2] ),
    .C(_08155_),
    .Y(_08157_));
 sky130_fd_sc_hd__or2b_1 _22901_ (.A(_08115_),
    .B_N(_08117_),
    .X(_08158_));
 sky130_fd_sc_hd__or2b_1 _22902_ (.A(_08117_),
    .B_N(_08115_),
    .X(_08159_));
 sky130_fd_sc_hd__nand2_1 _22903_ (.A(_08158_),
    .B(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand2_1 _22904_ (.A(_08160_),
    .B(\base_v_counter[1] ),
    .Y(_08161_));
 sky130_fd_sc_hd__nand3_1 _22905_ (.A(_08158_),
    .B(_08159_),
    .C(_09041_),
    .Y(_08162_));
 sky130_fd_sc_hd__xor2_1 _22906_ (.A(_08581_),
    .B(_08117_),
    .X(_08163_));
 sky130_fd_sc_hd__nand3_1 _22907_ (.A(_08161_),
    .B(_08162_),
    .C(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__inv_2 _22908_ (.A(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__nand2_1 _22909_ (.A(_08157_),
    .B(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__nor2_1 _22910_ (.A(_08156_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand3_1 _22911_ (.A(_08122_),
    .B(_08153_),
    .C(\base_v_counter[3] ),
    .Y(_08168_));
 sky130_fd_sc_hd__nand2_1 _22912_ (.A(_08167_),
    .B(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__nor2_1 _22913_ (.A(_08154_),
    .B(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__nand3_1 _22914_ (.A(_08149_),
    .B(\base_v_counter[4] ),
    .C(_08150_),
    .Y(_08171_));
 sky130_fd_sc_hd__nand3_1 _22915_ (.A(_08152_),
    .B(_08170_),
    .C(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_1 _22916_ (.A(_08150_),
    .B(_08126_),
    .Y(_08173_));
 sky130_fd_sc_hd__inv_2 _22917_ (.A(_08126_),
    .Y(_08174_));
 sky130_fd_sc_hd__nand2_1 _22918_ (.A(_08174_),
    .B(_08123_),
    .Y(_08175_));
 sky130_fd_sc_hd__nand2_1 _22919_ (.A(_08173_),
    .B(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__nand2_1 _22920_ (.A(_08176_),
    .B(\base_v_counter[5] ),
    .Y(_08177_));
 sky130_fd_sc_hd__nand3_1 _22921_ (.A(_08173_),
    .B(_08175_),
    .C(_08572_),
    .Y(_08178_));
 sky130_fd_sc_hd__nand2_1 _22922_ (.A(_08177_),
    .B(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__nor2_1 _22923_ (.A(_08172_),
    .B(_08179_),
    .Y(_08180_));
 sky130_fd_sc_hd__nand2_1 _22924_ (.A(_08137_),
    .B(_08606_),
    .Y(_08181_));
 sky130_fd_sc_hd__nand2_1 _22925_ (.A(_08102_),
    .B(_09125_),
    .Y(_08182_));
 sky130_fd_sc_hd__nand2_1 _22926_ (.A(_08136_),
    .B(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__nand3_1 _22927_ (.A(_08181_),
    .B(_08130_),
    .C(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__nand3b_1 _22928_ (.A_N(_08147_),
    .B(_08180_),
    .C(_08184_),
    .Y(_08185_));
 sky130_fd_sc_hd__nor2_1 _22929_ (.A(_08139_),
    .B(_08185_),
    .Y(_08186_));
 sky130_fd_sc_hd__inv_2 _22930_ (.A(_08183_),
    .Y(_08187_));
 sky130_fd_sc_hd__nand2_1 _22931_ (.A(_08131_),
    .B(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__nand2_1 _22932_ (.A(_08130_),
    .B(_08183_),
    .Y(_08189_));
 sky130_fd_sc_hd__a21oi_1 _22933_ (.A1(_08188_),
    .A2(_08189_),
    .B1(net4318),
    .Y(_08190_));
 sky130_fd_sc_hd__nand3_1 _22934_ (.A(_08188_),
    .B(_08189_),
    .C(net4318),
    .Y(_08191_));
 sky130_fd_sc_hd__nand2b_1 _22935_ (.A_N(_08181_),
    .B(_08189_),
    .Y(_08192_));
 sky130_fd_sc_hd__nand2_1 _22936_ (.A(_08191_),
    .B(_08192_),
    .Y(_08193_));
 sky130_fd_sc_hd__nor2_1 _22937_ (.A(_08190_),
    .B(_08193_),
    .Y(_08194_));
 sky130_fd_sc_hd__nand2_4 _22938_ (.A(_08186_),
    .B(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__nor2_1 _22939_ (.A(net4303),
    .B(_08723_),
    .Y(_08196_));
 sky130_fd_sc_hd__nand2_1 _22940_ (.A(_08195_),
    .B(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__or2_1 _22941_ (.A(net43),
    .B(net30),
    .X(_08198_));
 sky130_fd_sc_hd__nand2_1 _22942_ (.A(net43),
    .B(net30),
    .Y(_08199_));
 sky130_fd_sc_hd__nand2_1 _22943_ (.A(_08198_),
    .B(_08199_),
    .Y(_08200_));
 sky130_fd_sc_hd__inv_2 _22944_ (.A(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__nor2_1 _22945_ (.A(net46),
    .B(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_1 _22946_ (.A(_08201_),
    .B(net46),
    .Y(_08203_));
 sky130_fd_sc_hd__or3b_1 _22947_ (.A(_09222_),
    .B(_08202_),
    .C_N(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__nand2_1 _22948_ (.A(_08197_),
    .B(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__nand2_1 _22949_ (.A(_08205_),
    .B(_08081_),
    .Y(_08206_));
 sky130_fd_sc_hd__o21ai_1 _22950_ (.A1(_08581_),
    .A2(_08081_),
    .B1(_08206_),
    .Y(_02687_));
 sky130_fd_sc_hd__nor2_1 _22951_ (.A(net4312),
    .B(net4303),
    .Y(_08207_));
 sky130_fd_sc_hd__nand2_1 _22952_ (.A(net4312),
    .B(net4303),
    .Y(_08208_));
 sky130_fd_sc_hd__or3b_1 _22953_ (.A(_08722_),
    .B(_08207_),
    .C_N(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__inv_2 _22954_ (.A(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__nand2_1 _22955_ (.A(_08195_),
    .B(_08210_),
    .Y(_08211_));
 sky130_fd_sc_hd__and2_1 _22956_ (.A(_08203_),
    .B(_08199_),
    .X(_08212_));
 sky130_fd_sc_hd__or2_1 _22957_ (.A(net44),
    .B(net31),
    .X(_08213_));
 sky130_fd_sc_hd__nand2_1 _22958_ (.A(net44),
    .B(net31),
    .Y(_08214_));
 sky130_fd_sc_hd__nand2_1 _22959_ (.A(_08213_),
    .B(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__xor2_1 _22960_ (.A(net47),
    .B(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__nor2_1 _22961_ (.A(_08216_),
    .B(_08212_),
    .Y(_08217_));
 sky130_fd_sc_hd__inv_2 _22962_ (.A(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__nand2_1 _22963_ (.A(_08218_),
    .B(_08723_),
    .Y(_08219_));
 sky130_fd_sc_hd__a21o_1 _22964_ (.A1(_08212_),
    .A2(_08216_),
    .B1(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__nand2_1 _22965_ (.A(_08211_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__nand2_1 _22966_ (.A(_08221_),
    .B(_08081_),
    .Y(_08222_));
 sky130_fd_sc_hd__o21ai_1 _22967_ (.A1(_09041_),
    .A2(_08081_),
    .B1(_08222_),
    .Y(_02688_));
 sky130_fd_sc_hd__nor2_1 _22968_ (.A(_08593_),
    .B(_08208_),
    .Y(_08223_));
 sky130_fd_sc_hd__inv_2 _22969_ (.A(_08223_),
    .Y(_08224_));
 sky130_fd_sc_hd__nand2_1 _22970_ (.A(_08208_),
    .B(_08593_),
    .Y(_08225_));
 sky130_fd_sc_hd__and3_1 _22971_ (.A(_08224_),
    .B(_10310_),
    .C(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__nand2_1 _22972_ (.A(_08195_),
    .B(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__a21boi_1 _22973_ (.A1(_08213_),
    .A2(net47),
    .B1_N(_08214_),
    .Y(_08228_));
 sky130_fd_sc_hd__inv_2 _22974_ (.A(net48),
    .Y(_08229_));
 sky130_fd_sc_hd__or2_1 _22975_ (.A(net45),
    .B(net32),
    .X(_08230_));
 sky130_fd_sc_hd__nand2_1 _22976_ (.A(net45),
    .B(net32),
    .Y(_08231_));
 sky130_fd_sc_hd__nand2_1 _22977_ (.A(_08230_),
    .B(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__or2_1 _22978_ (.A(_08229_),
    .B(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__nand2_1 _22979_ (.A(_08232_),
    .B(_08229_),
    .Y(_08234_));
 sky130_fd_sc_hd__nand2_1 _22980_ (.A(_08233_),
    .B(_08234_),
    .Y(_08235_));
 sky130_fd_sc_hd__or2_1 _22981_ (.A(_08228_),
    .B(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__nand2_1 _22982_ (.A(_08235_),
    .B(_08228_),
    .Y(_08237_));
 sky130_fd_sc_hd__nand2_1 _22983_ (.A(_08236_),
    .B(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__or2_1 _22984_ (.A(_08218_),
    .B(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__nand2_1 _22985_ (.A(_08239_),
    .B(_08723_),
    .Y(_08240_));
 sky130_fd_sc_hd__a21o_1 _22986_ (.A1(_08218_),
    .A2(_08238_),
    .B1(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__nand2_1 _22987_ (.A(_08227_),
    .B(_08241_),
    .Y(_08242_));
 sky130_fd_sc_hd__nand2_1 _22988_ (.A(_08242_),
    .B(_08081_),
    .Y(_08243_));
 sky130_fd_sc_hd__o21ai_1 _22989_ (.A1(_08593_),
    .A2(_08081_),
    .B1(_08243_),
    .Y(_02689_));
 sky130_fd_sc_hd__nor2_1 _22990_ (.A(_08588_),
    .B(_08224_),
    .Y(_08244_));
 sky130_fd_sc_hd__inv_2 _22991_ (.A(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__nand2_1 _22992_ (.A(_08224_),
    .B(_08588_),
    .Y(_08246_));
 sky130_fd_sc_hd__and3_1 _22993_ (.A(_08245_),
    .B(_10310_),
    .C(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__nand2_1 _22994_ (.A(_08195_),
    .B(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__nand2_1 _22995_ (.A(_08233_),
    .B(_08231_),
    .Y(_08249_));
 sky130_fd_sc_hd__inv_2 _22996_ (.A(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__nor2_1 _22997_ (.A(_07799_),
    .B(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_1 _22998_ (.A(_08250_),
    .B(_07799_),
    .Y(_08252_));
 sky130_fd_sc_hd__or2b_1 _22999_ (.A(_08251_),
    .B_N(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__nand2_1 _23000_ (.A(_08239_),
    .B(_08236_),
    .Y(_08254_));
 sky130_fd_sc_hd__or2_1 _23001_ (.A(_08253_),
    .B(_08254_),
    .X(_08255_));
 sky130_fd_sc_hd__nand2_1 _23002_ (.A(_08254_),
    .B(_08253_),
    .Y(_08256_));
 sky130_fd_sc_hd__a21o_1 _23003_ (.A1(_08255_),
    .A2(_08256_),
    .B1(_03834_),
    .X(_08257_));
 sky130_fd_sc_hd__nand2_1 _23004_ (.A(_08248_),
    .B(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__nand2_1 _23005_ (.A(_08258_),
    .B(_08081_),
    .Y(_08259_));
 sky130_fd_sc_hd__o21ai_1 _23006_ (.A1(_08588_),
    .A2(_08081_),
    .B1(_08259_),
    .Y(_02690_));
 sky130_fd_sc_hd__nor2_1 _23007_ (.A(net4306),
    .B(_08244_),
    .Y(_08260_));
 sky130_fd_sc_hd__nor2_1 _23008_ (.A(_08577_),
    .B(_08245_),
    .Y(_08261_));
 sky130_fd_sc_hd__or3_1 _23009_ (.A(_08722_),
    .B(_08260_),
    .C(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__inv_2 _23010_ (.A(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__nand2_1 _23011_ (.A(_08195_),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__a21o_1 _23012_ (.A1(_08254_),
    .A2(_08252_),
    .B1(_08251_),
    .X(_08265_));
 sky130_fd_sc_hd__or2_1 _23013_ (.A(net34),
    .B(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__nand2_1 _23014_ (.A(_08265_),
    .B(net34),
    .Y(_08267_));
 sky130_fd_sc_hd__nand3_1 _23015_ (.A(_08266_),
    .B(_08723_),
    .C(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand2_1 _23016_ (.A(_08264_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__nand2_1 _23017_ (.A(_08269_),
    .B(_08081_),
    .Y(_08270_));
 sky130_fd_sc_hd__o21ai_1 _23018_ (.A1(_08577_),
    .A2(_08081_),
    .B1(_08270_),
    .Y(_02691_));
 sky130_fd_sc_hd__inv_2 _23019_ (.A(_08261_),
    .Y(_08271_));
 sky130_fd_sc_hd__nor2_1 _23020_ (.A(_08572_),
    .B(_08271_),
    .Y(_08272_));
 sky130_fd_sc_hd__nor2_1 _23021_ (.A(_08723_),
    .B(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__o21a_1 _23022_ (.A1(net4325),
    .A2(_08261_),
    .B1(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__nand2_1 _23023_ (.A(_08195_),
    .B(_08274_),
    .Y(_08275_));
 sky130_fd_sc_hd__nor2_1 _23024_ (.A(_07806_),
    .B(_08267_),
    .Y(_08276_));
 sky130_fd_sc_hd__or2_1 _23025_ (.A(_09222_),
    .B(_08276_),
    .X(_08277_));
 sky130_fd_sc_hd__a21o_1 _23026_ (.A1(_07806_),
    .A2(_08267_),
    .B1(_08277_),
    .X(_08278_));
 sky130_fd_sc_hd__nand2_1 _23027_ (.A(_08275_),
    .B(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__nand2_1 _23028_ (.A(_08279_),
    .B(_08081_),
    .Y(_08280_));
 sky130_fd_sc_hd__o21ai_1 _23029_ (.A1(_08572_),
    .A2(_08081_),
    .B1(_08280_),
    .Y(_02692_));
 sky130_fd_sc_hd__nor2_1 _23030_ (.A(net4298),
    .B(_08272_),
    .Y(_08281_));
 sky130_fd_sc_hd__nand2_1 _23031_ (.A(_08272_),
    .B(net4298),
    .Y(_08282_));
 sky130_fd_sc_hd__or3b_1 _23032_ (.A(_08722_),
    .B(_08281_),
    .C_N(_08282_),
    .X(_08283_));
 sky130_fd_sc_hd__inv_2 _23033_ (.A(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__nand2_1 _23034_ (.A(_08195_),
    .B(_08284_),
    .Y(_08285_));
 sky130_fd_sc_hd__nor2_1 _23035_ (.A(net36),
    .B(_08276_),
    .Y(_08286_));
 sky130_fd_sc_hd__nand2_1 _23036_ (.A(_08276_),
    .B(net36),
    .Y(_08287_));
 sky130_fd_sc_hd__inv_2 _23037_ (.A(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__or3_1 _23038_ (.A(_09222_),
    .B(_08286_),
    .C(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__nand2_1 _23039_ (.A(_08285_),
    .B(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__nand2_1 _23040_ (.A(_08290_),
    .B(_08081_),
    .Y(_08291_));
 sky130_fd_sc_hd__o21ai_1 _23041_ (.A1(_08562_),
    .A2(_08080_),
    .B1(_08291_),
    .Y(_02693_));
 sky130_fd_sc_hd__nor2_1 _23042_ (.A(_08565_),
    .B(_08282_),
    .Y(_08292_));
 sky130_fd_sc_hd__nand2_1 _23043_ (.A(_08282_),
    .B(_08565_),
    .Y(_08293_));
 sky130_fd_sc_hd__or3b_1 _23044_ (.A(_08722_),
    .B(_08292_),
    .C_N(_08293_),
    .X(_08294_));
 sky130_fd_sc_hd__inv_2 _23045_ (.A(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__nand2_1 _23046_ (.A(_08195_),
    .B(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__inv_2 _23047_ (.A(net37),
    .Y(_08297_));
 sky130_fd_sc_hd__nor2_1 _23048_ (.A(_08297_),
    .B(_08287_),
    .Y(_08298_));
 sky130_fd_sc_hd__nor2_1 _23049_ (.A(_09223_),
    .B(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__o21ai_1 _23050_ (.A1(net37),
    .A2(_08288_),
    .B1(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__nand2_1 _23051_ (.A(_08296_),
    .B(_08300_),
    .Y(_08301_));
 sky130_fd_sc_hd__nand2_1 _23052_ (.A(_08301_),
    .B(_08081_),
    .Y(_08302_));
 sky130_fd_sc_hd__o21ai_1 _23053_ (.A1(_08565_),
    .A2(_08080_),
    .B1(_08302_),
    .Y(_02694_));
 sky130_fd_sc_hd__or2_1 _23054_ (.A(net4318),
    .B(_08292_),
    .X(_08303_));
 sky130_fd_sc_hd__nand2_1 _23055_ (.A(_08292_),
    .B(net4318),
    .Y(_08304_));
 sky130_fd_sc_hd__and3_1 _23056_ (.A(_08303_),
    .B(_10310_),
    .C(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__nand2_1 _23057_ (.A(_08195_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__inv_2 _23058_ (.A(_08298_),
    .Y(_08307_));
 sky130_fd_sc_hd__a21o_1 _23059_ (.A1(_08298_),
    .A2(net38),
    .B1(_08776_),
    .X(_08308_));
 sky130_fd_sc_hd__a21o_1 _23060_ (.A1(_07815_),
    .A2(_08307_),
    .B1(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__nand2_1 _23061_ (.A(_08306_),
    .B(_08309_),
    .Y(_08310_));
 sky130_fd_sc_hd__nand2_1 _23062_ (.A(_08310_),
    .B(_08081_),
    .Y(_08311_));
 sky130_fd_sc_hd__o21ai_1 _23063_ (.A1(_08584_),
    .A2(_08080_),
    .B1(_08311_),
    .Y(_02695_));
 sky130_fd_sc_hd__a21oi_1 _23064_ (.A1(_08304_),
    .A2(_08606_),
    .B1(_08723_),
    .Y(_08312_));
 sky130_fd_sc_hd__o21a_1 _23065_ (.A1(_08606_),
    .A2(_08304_),
    .B1(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__nand2_1 _23066_ (.A(_08195_),
    .B(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__or3_1 _23067_ (.A(_09222_),
    .B(_07815_),
    .C(_08307_),
    .X(_08315_));
 sky130_fd_sc_hd__nand2_1 _23068_ (.A(_08314_),
    .B(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__nand2_1 _23069_ (.A(_08316_),
    .B(_08081_),
    .Y(_08317_));
 sky130_fd_sc_hd__o21ai_1 _23070_ (.A1(_08606_),
    .A2(_08080_),
    .B1(_08317_),
    .Y(_02696_));
 sky130_fd_sc_hd__buf_8 _23071_ (.A(_08050_),
    .X(_08318_));
 sky130_fd_sc_hd__nand2_1 _23072_ (.A(_08785_),
    .B(_09222_),
    .Y(_08319_));
 sky130_fd_sc_hd__inv_2 _23073_ (.A(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__nand3_1 _23074_ (.A(_08318_),
    .B(_08696_),
    .C(_08320_),
    .Y(_08321_));
 sky130_fd_sc_hd__nand3_2 _23075_ (.A(_08050_),
    .B(_08614_),
    .C(_08051_),
    .Y(_08322_));
 sky130_fd_sc_hd__nor2_1 _23076_ (.A(_08722_),
    .B(_08655_),
    .Y(_08323_));
 sky130_fd_sc_hd__and2_1 _23077_ (.A(_08802_),
    .B(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__nand2_1 _23078_ (.A(_08318_),
    .B(_08324_),
    .Y(_08325_));
 sky130_fd_sc_hd__nand3_4 _23079_ (.A(_08322_),
    .B(_08792_),
    .C(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__buf_6 _23080_ (.A(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__nand2_1 _23081_ (.A(_08327_),
    .B(net2770),
    .Y(_08328_));
 sky130_fd_sc_hd__o21ai_1 _23082_ (.A1(_08321_),
    .A2(_08327_),
    .B1(_08328_),
    .Y(_02697_));
 sky130_fd_sc_hd__o211ai_1 _23083_ (.A1(_05012_),
    .A2(_05017_),
    .B1(_08320_),
    .C1(_08318_),
    .Y(_08329_));
 sky130_fd_sc_hd__nand2_1 _23084_ (.A(_08327_),
    .B(net3038),
    .Y(_08330_));
 sky130_fd_sc_hd__o21ai_1 _23085_ (.A1(_08329_),
    .A2(_08327_),
    .B1(_08330_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_1 _23086_ (.A(_05024_),
    .B(net3919),
    .Y(_08331_));
 sky130_fd_sc_hd__nand2_1 _23087_ (.A(_05023_),
    .B(_05029_),
    .Y(_08332_));
 sky130_fd_sc_hd__and3_1 _23088_ (.A(_08331_),
    .B(_10310_),
    .C(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__nand3_1 _23089_ (.A(_08318_),
    .B(_08720_),
    .C(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__nand2_1 _23090_ (.A(_08327_),
    .B(net3919),
    .Y(_08335_));
 sky130_fd_sc_hd__o21ai_1 _23091_ (.A1(_08334_),
    .A2(_08327_),
    .B1(_08335_),
    .Y(_02699_));
 sky130_fd_sc_hd__nand2_1 _23092_ (.A(_08331_),
    .B(_08705_),
    .Y(_08336_));
 sky130_fd_sc_hd__and3_1 _23093_ (.A(_08336_),
    .B(_10310_),
    .C(_05062_),
    .X(_08337_));
 sky130_fd_sc_hd__nand3_1 _23094_ (.A(_08318_),
    .B(_08720_),
    .C(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__nand2_1 _23095_ (.A(_08327_),
    .B(net2785),
    .Y(_08339_));
 sky130_fd_sc_hd__o21ai_1 _23096_ (.A1(_08338_),
    .A2(_08327_),
    .B1(_08339_),
    .Y(_02700_));
 sky130_fd_sc_hd__nor2_1 _23097_ (.A(net4288),
    .B(_05061_),
    .Y(_08340_));
 sky130_fd_sc_hd__nor2_1 _23098_ (.A(_08684_),
    .B(_05062_),
    .Y(_08341_));
 sky130_fd_sc_hd__nor2_1 _23099_ (.A(_08340_),
    .B(_08341_),
    .Y(_08342_));
 sky130_fd_sc_hd__nand3_1 _23100_ (.A(_08318_),
    .B(_08320_),
    .C(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__nand2_1 _23101_ (.A(_08327_),
    .B(net4288),
    .Y(_08344_));
 sky130_fd_sc_hd__o21ai_1 _23102_ (.A1(_08343_),
    .A2(_08327_),
    .B1(_08344_),
    .Y(_02701_));
 sky130_fd_sc_hd__or2_1 _23103_ (.A(net4186),
    .B(_08341_),
    .X(_08345_));
 sky130_fd_sc_hd__nand2_1 _23104_ (.A(_05061_),
    .B(_05088_),
    .Y(_08346_));
 sky130_fd_sc_hd__and3_1 _23105_ (.A(_08345_),
    .B(_10310_),
    .C(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__nand3_1 _23106_ (.A(_08318_),
    .B(_08720_),
    .C(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nand2_1 _23107_ (.A(_08327_),
    .B(net4186),
    .Y(_08349_));
 sky130_fd_sc_hd__o21ai_1 _23108_ (.A1(_08348_),
    .A2(_08327_),
    .B1(_08349_),
    .Y(_02702_));
 sky130_fd_sc_hd__or2_1 _23109_ (.A(_08709_),
    .B(_08346_),
    .X(_08350_));
 sky130_fd_sc_hd__nand2_1 _23110_ (.A(_08346_),
    .B(_08709_),
    .Y(_08351_));
 sky130_fd_sc_hd__and3_1 _23111_ (.A(_08350_),
    .B(_10310_),
    .C(_08351_),
    .X(_08352_));
 sky130_fd_sc_hd__nand3_1 _23112_ (.A(_08318_),
    .B(_08720_),
    .C(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand2_1 _23113_ (.A(_08327_),
    .B(net2750),
    .Y(_08354_));
 sky130_fd_sc_hd__o21ai_1 _23114_ (.A1(_08353_),
    .A2(_08326_),
    .B1(_08354_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand2_1 _23115_ (.A(_08350_),
    .B(_08662_),
    .Y(_08355_));
 sky130_fd_sc_hd__and3_1 _23116_ (.A(_08355_),
    .B(_10310_),
    .C(_05219_),
    .X(_08356_));
 sky130_fd_sc_hd__nand3_1 _23117_ (.A(_08318_),
    .B(_08720_),
    .C(_08356_),
    .Y(_08357_));
 sky130_fd_sc_hd__nand2_1 _23118_ (.A(_08327_),
    .B(net3652),
    .Y(_08358_));
 sky130_fd_sc_hd__o21ai_1 _23119_ (.A1(_08357_),
    .A2(_08326_),
    .B1(_08358_),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2_1 _23120_ (.A(_05219_),
    .B(_05188_),
    .Y(_08359_));
 sky130_fd_sc_hd__nand2_1 _23121_ (.A(_05218_),
    .B(_05113_),
    .Y(_08360_));
 sky130_fd_sc_hd__and3_1 _23122_ (.A(_08359_),
    .B(_10310_),
    .C(_08360_),
    .X(_08361_));
 sky130_fd_sc_hd__nand3_1 _23123_ (.A(_08318_),
    .B(_08720_),
    .C(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__nand2_1 _23124_ (.A(_08327_),
    .B(_05113_),
    .Y(_08363_));
 sky130_fd_sc_hd__o21ai_1 _23125_ (.A1(_08362_),
    .A2(_08326_),
    .B1(_08363_),
    .Y(_02705_));
 sky130_fd_sc_hd__nand2_1 _23126_ (.A(_08360_),
    .B(_08700_),
    .Y(_08364_));
 sky130_fd_sc_hd__o21a_1 _23127_ (.A1(_08700_),
    .A2(_08360_),
    .B1(_08800_),
    .X(_08365_));
 sky130_fd_sc_hd__nand3_1 _23128_ (.A(_08318_),
    .B(_08364_),
    .C(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__nand2_1 _23129_ (.A(_08327_),
    .B(net1859),
    .Y(_08367_));
 sky130_fd_sc_hd__o21ai_1 _23130_ (.A1(_08366_),
    .A2(_08326_),
    .B1(_08367_),
    .Y(_02706_));
 sky130_fd_sc_hd__inv_2 _23131_ (.A(net2958),
    .Y(_08368_));
 sky130_fd_sc_hd__inv_2 _23132_ (.A(_08774_),
    .Y(_08369_));
 sky130_fd_sc_hd__nor2_1 _23133_ (.A(_08368_),
    .B(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__nor2_1 _23134_ (.A(\res_v_active[0] ),
    .B(\res_v_active[1] ),
    .Y(_08371_));
 sky130_fd_sc_hd__inv_2 _23135_ (.A(\res_v_active[2] ),
    .Y(_08372_));
 sky130_fd_sc_hd__nand2_1 _23136_ (.A(_08371_),
    .B(_08372_),
    .Y(_08373_));
 sky130_fd_sc_hd__or2_1 _23137_ (.A(\res_v_active[3] ),
    .B(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__nor2_1 _23138_ (.A(\res_v_active[4] ),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__inv_2 _23139_ (.A(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__or2_1 _23140_ (.A(\res_v_active[5] ),
    .B(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__nor2_1 _23141_ (.A(net2757),
    .B(_08377_),
    .Y(_08378_));
 sky130_fd_sc_hd__inv_2 _23142_ (.A(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand2_1 _23143_ (.A(_08374_),
    .B(net2772),
    .Y(_08380_));
 sky130_fd_sc_hd__nand2_1 _23144_ (.A(_08376_),
    .B(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__xor2_1 _23145_ (.A(\res_v_counter[4] ),
    .B(_08381_),
    .X(_08382_));
 sky130_fd_sc_hd__inv_2 _23146_ (.A(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__nand2_1 _23147_ (.A(_08377_),
    .B(\res_v_active[6] ),
    .Y(_08384_));
 sky130_fd_sc_hd__nand2_1 _23148_ (.A(_08379_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__or2_1 _23149_ (.A(_07655_),
    .B(_08385_),
    .X(_08386_));
 sky130_fd_sc_hd__nand2_1 _23150_ (.A(_08376_),
    .B(\res_v_active[5] ),
    .Y(_08387_));
 sky130_fd_sc_hd__nand2_1 _23151_ (.A(_08377_),
    .B(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__nand2_1 _23152_ (.A(_08388_),
    .B(_07652_),
    .Y(_08389_));
 sky130_fd_sc_hd__nand2_1 _23153_ (.A(_08385_),
    .B(_07655_),
    .Y(_08390_));
 sky130_fd_sc_hd__and3_1 _23154_ (.A(_08386_),
    .B(_08389_),
    .C(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__a21o_1 _23155_ (.A1(_08379_),
    .A2(\res_v_active[7] ),
    .B1(_07654_),
    .X(_08392_));
 sky130_fd_sc_hd__nand2_1 _23156_ (.A(_08373_),
    .B(\res_v_active[3] ),
    .Y(_08393_));
 sky130_fd_sc_hd__nand2_1 _23157_ (.A(_08374_),
    .B(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__or2_1 _23158_ (.A(_08372_),
    .B(_08371_),
    .X(_08395_));
 sky130_fd_sc_hd__nand2_1 _23159_ (.A(_08395_),
    .B(_08373_),
    .Y(_08396_));
 sky130_fd_sc_hd__nand2_1 _23160_ (.A(_08396_),
    .B(_07660_),
    .Y(_08397_));
 sky130_fd_sc_hd__or2_1 _23161_ (.A(_07660_),
    .B(_08396_),
    .X(_08398_));
 sky130_fd_sc_hd__xnor2_1 _23162_ (.A(\res_v_counter[1] ),
    .B(\res_v_active[1] ),
    .Y(_08399_));
 sky130_fd_sc_hd__nand2_1 _23163_ (.A(_08368_),
    .B(\res_v_active[0] ),
    .Y(_08400_));
 sky130_fd_sc_hd__o21ai_1 _23164_ (.A1(\res_v_active[0] ),
    .A2(_08399_),
    .B1(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__o211ai_1 _23165_ (.A1(\res_v_counter[0] ),
    .A2(_08399_),
    .B1(_07657_),
    .C1(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__a21oi_1 _23166_ (.A1(_07659_),
    .A2(_08394_),
    .B1(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__o2111a_1 _23167_ (.A1(_07659_),
    .A2(_08394_),
    .B1(_08397_),
    .C1(_08398_),
    .D1(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__or3b_1 _23168_ (.A(net2729),
    .B(_08378_),
    .C_N(\res_v_active[7] ),
    .X(_08405_));
 sky130_fd_sc_hd__o2111a_1 _23169_ (.A1(_07652_),
    .A2(_08388_),
    .B1(_08392_),
    .C1(_08404_),
    .D1(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__o2111ai_4 _23170_ (.A1(\res_v_active[7] ),
    .A2(_08379_),
    .B1(_08383_),
    .C1(_08391_),
    .D1(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__and3_1 _23171_ (.A(_08369_),
    .B(_08368_),
    .C(_08407_),
    .X(_08408_));
 sky130_fd_sc_hd__o21ai_1 _23172_ (.A1(_08370_),
    .A2(_08408_),
    .B1(_08051_),
    .Y(_08409_));
 sky130_fd_sc_hd__nor2_4 _23173_ (.A(_08318_),
    .B(_08195_),
    .Y(_08410_));
 sky130_fd_sc_hd__o22ai_1 _23174_ (.A1(_08368_),
    .A2(_04971_),
    .B1(_08409_),
    .B2(_08410_),
    .Y(_02707_));
 sky130_fd_sc_hd__inv_2 _23175_ (.A(net2778),
    .Y(_08411_));
 sky130_fd_sc_hd__nor2_1 _23176_ (.A(_08411_),
    .B(_08369_),
    .Y(_08412_));
 sky130_fd_sc_hd__nand2_1 _23177_ (.A(net2778),
    .B(\res_v_counter[0] ),
    .Y(_08413_));
 sky130_fd_sc_hd__inv_2 _23178_ (.A(_08413_),
    .Y(_08414_));
 sky130_fd_sc_hd__nor2_1 _23179_ (.A(_07658_),
    .B(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__and3_1 _23180_ (.A(_08369_),
    .B(_08407_),
    .C(_08415_),
    .X(_08416_));
 sky130_fd_sc_hd__o21ai_1 _23181_ (.A1(_08412_),
    .A2(_08416_),
    .B1(_08051_),
    .Y(_08417_));
 sky130_fd_sc_hd__o22ai_1 _23182_ (.A1(_08411_),
    .A2(_04971_),
    .B1(_08417_),
    .B2(_08410_),
    .Y(_02708_));
 sky130_fd_sc_hd__xor2_1 _23183_ (.A(net2691),
    .B(_08413_),
    .X(_08418_));
 sky130_fd_sc_hd__or3b_1 _23184_ (.A(_08418_),
    .B(_08774_),
    .C_N(_08407_),
    .X(_08419_));
 sky130_fd_sc_hd__nand2_1 _23185_ (.A(_08774_),
    .B(net2691),
    .Y(_08420_));
 sky130_fd_sc_hd__inv_2 _23186_ (.A(_08051_),
    .Y(_08421_));
 sky130_fd_sc_hd__a21o_1 _23187_ (.A1(_08419_),
    .A2(_08420_),
    .B1(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__nand2_1 _23188_ (.A(_08793_),
    .B(net2691),
    .Y(_08423_));
 sky130_fd_sc_hd__o21ai_1 _23189_ (.A1(_08410_),
    .A2(_08422_),
    .B1(net2692),
    .Y(_02709_));
 sky130_fd_sc_hd__and3_1 _23190_ (.A(_08414_),
    .B(net2826),
    .C(net2691),
    .X(_08424_));
 sky130_fd_sc_hd__inv_2 _23191_ (.A(_08424_),
    .Y(_08425_));
 sky130_fd_sc_hd__o21ai_1 _23192_ (.A1(_07660_),
    .A2(_08413_),
    .B1(_07659_),
    .Y(_08426_));
 sky130_fd_sc_hd__a31o_1 _23193_ (.A1(_08407_),
    .A2(_08425_),
    .A3(_08426_),
    .B1(_08774_),
    .X(_08427_));
 sky130_fd_sc_hd__o211ai_1 _23194_ (.A1(net2826),
    .A2(_08369_),
    .B1(_08051_),
    .C1(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__o22ai_1 _23195_ (.A1(_07659_),
    .A2(_04971_),
    .B1(_08428_),
    .B2(_08410_),
    .Y(_02710_));
 sky130_fd_sc_hd__nor2_1 _23196_ (.A(_07653_),
    .B(_08369_),
    .Y(_08429_));
 sky130_fd_sc_hd__nor2_1 _23197_ (.A(net3517),
    .B(_08424_),
    .Y(_08430_));
 sky130_fd_sc_hd__nor2_1 _23198_ (.A(_07653_),
    .B(_08425_),
    .Y(_08431_));
 sky130_fd_sc_hd__or3b_1 _23199_ (.A(_08430_),
    .B(_08431_),
    .C_N(_08407_),
    .X(_08432_));
 sky130_fd_sc_hd__nor2_1 _23200_ (.A(_08774_),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__o21ai_1 _23201_ (.A1(_08429_),
    .A2(_08433_),
    .B1(_08051_),
    .Y(_08434_));
 sky130_fd_sc_hd__o22ai_1 _23202_ (.A1(_07653_),
    .A2(_04971_),
    .B1(_08434_),
    .B2(_08410_),
    .Y(_02711_));
 sky130_fd_sc_hd__or2_1 _23203_ (.A(net3018),
    .B(_08431_),
    .X(_08435_));
 sky130_fd_sc_hd__nand2_1 _23204_ (.A(_08431_),
    .B(net3018),
    .Y(_08436_));
 sky130_fd_sc_hd__nand3_1 _23205_ (.A(_08407_),
    .B(_08435_),
    .C(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__nor2_1 _23206_ (.A(_08437_),
    .B(_08774_),
    .Y(_08438_));
 sky130_fd_sc_hd__nor2_1 _23207_ (.A(_07652_),
    .B(_08369_),
    .Y(_08439_));
 sky130_fd_sc_hd__o21ai_1 _23208_ (.A1(_08438_),
    .A2(_08439_),
    .B1(_08051_),
    .Y(_08440_));
 sky130_fd_sc_hd__o22ai_1 _23209_ (.A1(_07652_),
    .A2(_04971_),
    .B1(_08440_),
    .B2(_08410_),
    .Y(_02712_));
 sky130_fd_sc_hd__or2_1 _23210_ (.A(_07655_),
    .B(_08436_),
    .X(_08441_));
 sky130_fd_sc_hd__nand2_1 _23211_ (.A(_08436_),
    .B(_07655_),
    .Y(_08442_));
 sky130_fd_sc_hd__nand2_1 _23212_ (.A(_08441_),
    .B(_08442_),
    .Y(_08443_));
 sky130_fd_sc_hd__or3b_1 _23213_ (.A(_08443_),
    .B(_08774_),
    .C_N(_08407_),
    .X(_08444_));
 sky130_fd_sc_hd__nand2_1 _23214_ (.A(_08774_),
    .B(net2668),
    .Y(_08445_));
 sky130_fd_sc_hd__a21o_1 _23215_ (.A1(_08444_),
    .A2(_08445_),
    .B1(_08421_),
    .X(_08446_));
 sky130_fd_sc_hd__nand2_1 _23216_ (.A(_08793_),
    .B(net2668),
    .Y(_08447_));
 sky130_fd_sc_hd__o21ai_1 _23217_ (.A1(_08410_),
    .A2(_08446_),
    .B1(net2669),
    .Y(_02713_));
 sky130_fd_sc_hd__or2_1 _23218_ (.A(_07654_),
    .B(_08441_),
    .X(_08448_));
 sky130_fd_sc_hd__a21o_1 _23219_ (.A1(_08407_),
    .A2(_08448_),
    .B1(_08774_),
    .X(_08449_));
 sky130_fd_sc_hd__o21ai_1 _23220_ (.A1(_08441_),
    .A2(_08774_),
    .B1(_07654_),
    .Y(_08450_));
 sky130_fd_sc_hd__nand3_1 _23221_ (.A(_08449_),
    .B(_08450_),
    .C(_08051_),
    .Y(_08451_));
 sky130_fd_sc_hd__o22ai_1 _23222_ (.A1(_07654_),
    .A2(_04971_),
    .B1(_08451_),
    .B2(_08410_),
    .Y(_02714_));
 sky130_fd_sc_hd__or2_1 _23223_ (.A(net2685),
    .B(_08448_),
    .X(_08452_));
 sky130_fd_sc_hd__or3b_1 _23224_ (.A(_08452_),
    .B(_08774_),
    .C_N(_08407_),
    .X(_08453_));
 sky130_fd_sc_hd__nand2_1 _23225_ (.A(_08449_),
    .B(net2685),
    .Y(_08454_));
 sky130_fd_sc_hd__a21o_1 _23226_ (.A1(_08453_),
    .A2(_08454_),
    .B1(_08421_),
    .X(_08455_));
 sky130_fd_sc_hd__nand2_1 _23227_ (.A(_08793_),
    .B(net2685),
    .Y(_08456_));
 sky130_fd_sc_hd__o21ai_1 _23228_ (.A1(_08410_),
    .A2(_08455_),
    .B1(_08456_),
    .Y(_02715_));
 sky130_fd_sc_hd__or2b_1 _23229_ (.A(_08193_),
    .B_N(_08184_),
    .X(_08457_));
 sky130_fd_sc_hd__nor3_1 _23230_ (.A(_08172_),
    .B(_08179_),
    .C(_08147_),
    .Y(_08458_));
 sky130_fd_sc_hd__nor3b_1 _23231_ (.A(_08190_),
    .B(_08139_),
    .C_N(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__inv_2 _23232_ (.A(_08318_),
    .Y(_08460_));
 sky130_fd_sc_hd__nand3b_1 _23233_ (.A_N(_08457_),
    .B(_08459_),
    .C(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__nor3b_1 _23234_ (.A(_08448_),
    .B(_08661_),
    .C_N(net2685),
    .Y(_08462_));
 sky130_fd_sc_hd__xnor2_1 _23235_ (.A(net2687),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__or3_2 _23236_ (.A(_08772_),
    .B(_08720_),
    .C(_08614_),
    .X(_08464_));
 sky130_fd_sc_hd__or2_1 _23237_ (.A(_08463_),
    .B(_08464_),
    .X(_08465_));
 sky130_fd_sc_hd__nand2_1 _23238_ (.A(_08464_),
    .B(net2687),
    .Y(_08466_));
 sky130_fd_sc_hd__a21oi_1 _23239_ (.A1(_08465_),
    .A2(_08466_),
    .B1(_08421_),
    .Y(_08467_));
 sky130_fd_sc_hd__nand2_1 _23240_ (.A(_08461_),
    .B(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__nand2_1 _23241_ (.A(_08793_),
    .B(net2687),
    .Y(_08469_));
 sky130_fd_sc_hd__nand2_1 _23242_ (.A(_08468_),
    .B(net2688),
    .Y(_02716_));
 sky130_fd_sc_hd__mux2_1 _23243_ (.A0(net84),
    .A1(net3788),
    .S(_07857_),
    .X(_08470_));
 sky130_fd_sc_hd__clkbuf_1 _23244_ (.A(_08470_),
    .X(_02717_));
 sky130_fd_sc_hd__mux2_1 _23245_ (.A0(net85),
    .A1(net3910),
    .S(_07857_),
    .X(_08471_));
 sky130_fd_sc_hd__clkbuf_1 _23246_ (.A(_08471_),
    .X(_02718_));
 sky130_fd_sc_hd__mux2_1 _23247_ (.A0(net86),
    .A1(net3819),
    .S(_07857_),
    .X(_08472_));
 sky130_fd_sc_hd__clkbuf_1 _23248_ (.A(_08472_),
    .X(_02719_));
 sky130_fd_sc_hd__mux2_1 _23249_ (.A0(net87),
    .A1(net2761),
    .S(_07857_),
    .X(_08473_));
 sky130_fd_sc_hd__clkbuf_1 _23250_ (.A(_08473_),
    .X(_02720_));
 sky130_fd_sc_hd__mux2_1 _23251_ (.A0(net88),
    .A1(net4292),
    .S(_07857_),
    .X(_08474_));
 sky130_fd_sc_hd__clkbuf_1 _23252_ (.A(_08474_),
    .X(_02721_));
 sky130_fd_sc_hd__mux2_1 _23253_ (.A0(net89),
    .A1(net3633),
    .S(_09375_),
    .X(_08475_));
 sky130_fd_sc_hd__clkbuf_1 _23254_ (.A(_08475_),
    .X(_02722_));
 sky130_fd_sc_hd__mux2_1 _23255_ (.A0(net90),
    .A1(net2775),
    .S(_09375_),
    .X(_08476_));
 sky130_fd_sc_hd__clkbuf_1 _23256_ (.A(_08476_),
    .X(_02723_));
 sky130_fd_sc_hd__mux2_1 _23257_ (.A0(net91),
    .A1(net2999),
    .S(_09375_),
    .X(_08477_));
 sky130_fd_sc_hd__clkbuf_1 _23258_ (.A(_08477_),
    .X(_02724_));
 sky130_fd_sc_hd__nand2_2 _23259_ (.A(_08322_),
    .B(_04971_),
    .Y(_08478_));
 sky130_fd_sc_hd__nand2_1 _23260_ (.A(_08323_),
    .B(_08639_),
    .Y(_08479_));
 sky130_fd_sc_hd__or2_1 _23261_ (.A(_08479_),
    .B(_08460_),
    .X(_08480_));
 sky130_fd_sc_hd__nand2_1 _23262_ (.A(_08478_),
    .B(net2648),
    .Y(_08481_));
 sky130_fd_sc_hd__o21ai_1 _23263_ (.A1(_08478_),
    .A2(_08480_),
    .B1(_08481_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_1 _23264_ (.A(_08639_),
    .B(_08634_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand2_1 _23265_ (.A(net2648),
    .B(net2655),
    .Y(_08483_));
 sky130_fd_sc_hd__and3_1 _23266_ (.A(_08323_),
    .B(_08482_),
    .C(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__nand2_1 _23267_ (.A(_08318_),
    .B(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__nand2_1 _23268_ (.A(_08478_),
    .B(net2655),
    .Y(_08486_));
 sky130_fd_sc_hd__o21ai_1 _23269_ (.A1(_08485_),
    .A2(_08478_),
    .B1(_08486_),
    .Y(_02726_));
 sky130_fd_sc_hd__nand2_1 _23270_ (.A(_08483_),
    .B(_08651_),
    .Y(_08487_));
 sky130_fd_sc_hd__or2_1 _23271_ (.A(_08651_),
    .B(_08483_),
    .X(_08488_));
 sky130_fd_sc_hd__and3_1 _23272_ (.A(_08323_),
    .B(_08487_),
    .C(_08488_),
    .X(_08489_));
 sky130_fd_sc_hd__nand2_1 _23273_ (.A(_08318_),
    .B(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_1 _23274_ (.A(_08478_),
    .B(net1912),
    .Y(_08491_));
 sky130_fd_sc_hd__o21ai_1 _23275_ (.A1(_08490_),
    .A2(_08478_),
    .B1(net1913),
    .Y(_02727_));
 sky130_fd_sc_hd__a21oi_1 _23276_ (.A1(_08488_),
    .A2(_08647_),
    .B1(_08723_),
    .Y(_08492_));
 sky130_fd_sc_hd__o211a_1 _23277_ (.A1(_08647_),
    .A2(_08488_),
    .B1(_08492_),
    .C1(_08772_),
    .X(_08493_));
 sky130_fd_sc_hd__nand2_1 _23278_ (.A(_08318_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__nand2_1 _23279_ (.A(_08478_),
    .B(net1876),
    .Y(_08495_));
 sky130_fd_sc_hd__o21ai_1 _23280_ (.A1(_08494_),
    .A2(_08478_),
    .B1(net1877),
    .Y(_02728_));
 sky130_fd_sc_hd__nand2_1 _23281_ (.A(_08661_),
    .B(_08776_),
    .Y(_08496_));
 sky130_fd_sc_hd__nor2_1 _23282_ (.A(net4058),
    .B(_08496_),
    .Y(_08497_));
 sky130_fd_sc_hd__o211ai_2 _23283_ (.A1(_08772_),
    .A2(_08785_),
    .B1(_08633_),
    .C1(_05882_),
    .Y(_08498_));
 sky130_fd_sc_hd__o21ai_4 _23284_ (.A1(_08723_),
    .A2(_08802_),
    .B1(_08498_),
    .Y(_08499_));
 sky130_fd_sc_hd__mux2_1 _23285_ (.A0(_08497_),
    .A1(net4058),
    .S(_08499_),
    .X(_08500_));
 sky130_fd_sc_hd__clkbuf_1 _23286_ (.A(_08500_),
    .X(_02729_));
 sky130_fd_sc_hd__or2b_1 _23287_ (.A(net2660),
    .B_N(\line_double_counter[0] ),
    .X(_08501_));
 sky130_fd_sc_hd__o21ai_1 _23288_ (.A1(_08497_),
    .A2(_08499_),
    .B1(net2660),
    .Y(_08502_));
 sky130_fd_sc_hd__o31ai_1 _23289_ (.A1(_08496_),
    .A2(_08501_),
    .A3(_08499_),
    .B1(net2661),
    .Y(_02730_));
 sky130_fd_sc_hd__a21oi_1 _23290_ (.A1(\line_double_counter[0] ),
    .A2(net2660),
    .B1(net2677),
    .Y(_08503_));
 sky130_fd_sc_hd__and3_1 _23291_ (.A(\line_double_counter[0] ),
    .B(net2660),
    .C(net2677),
    .X(_08504_));
 sky130_fd_sc_hd__or2_1 _23292_ (.A(_08503_),
    .B(_08504_),
    .X(_08505_));
 sky130_fd_sc_hd__nand2_1 _23293_ (.A(_08499_),
    .B(net2677),
    .Y(_08506_));
 sky130_fd_sc_hd__o31ai_1 _23294_ (.A1(_08496_),
    .A2(_08505_),
    .A3(_08499_),
    .B1(net2678),
    .Y(_02731_));
 sky130_fd_sc_hd__xnor2_1 _23295_ (.A(net2680),
    .B(_08504_),
    .Y(_08507_));
 sky130_fd_sc_hd__nand2_1 _23296_ (.A(_08499_),
    .B(net2680),
    .Y(_08508_));
 sky130_fd_sc_hd__o31ai_1 _23297_ (.A1(_08496_),
    .A2(_08507_),
    .A3(_08499_),
    .B1(net2681),
    .Y(_02732_));
 sky130_fd_sc_hd__dfstp_1 _23298_ (.CLK(clknet_leaf_21_clk_i),
    .D(net2703),
    .SET_B(net168),
    .Q(\fb_read_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23299_ (.CLK(clknet_leaf_21_clk_i),
    .D(net4317),
    .RESET_B(net168),
    .Q(\fb_read_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _23300_ (.CLK(clknet_leaf_21_clk_i),
    .D(net2715),
    .RESET_B(net168),
    .Q(\fb_read_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _23301_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02572_),
    .RESET_B(net253),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_4 _23302_ (.CLK(clknet_leaf_283_clk_i),
    .D(net4222),
    .RESET_B(net270),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_2 _23303_ (.CLK(clknet_leaf_24_clk_i),
    .D(_02574_),
    .RESET_B(net172),
    .Q(\line_cache_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23304_ (.CLK(clknet_leaf_24_clk_i),
    .D(net2782),
    .RESET_B(net172),
    .Q(\line_cache_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23305_ (.CLK(clknet_leaf_33_clk_i),
    .D(net3792),
    .RESET_B(net194),
    .Q(\line_cache_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23306_ (.CLK(clknet_leaf_33_clk_i),
    .D(net2788),
    .RESET_B(net194),
    .Q(\line_cache_idx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _23307_ (.CLK(clknet_leaf_33_clk_i),
    .D(net3900),
    .RESET_B(net172),
    .Q(\line_cache_idx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _23308_ (.CLK(clknet_leaf_33_clk_i),
    .D(net2928),
    .RESET_B(net194),
    .Q(\line_cache_idx[7] ));
 sky130_fd_sc_hd__dfrtp_4 _23309_ (.CLK(clknet_leaf_24_clk_i),
    .D(_02580_),
    .RESET_B(net172),
    .Q(\line_cache_idx[8] ));
 sky130_fd_sc_hd__dfrtp_1 _23310_ (.CLK(clknet_leaf_24_clk_i),
    .D(_02581_),
    .RESET_B(net173),
    .Q(\line_cache_idx[9] ));
 sky130_fd_sc_hd__dfrtp_1 _23311_ (.CLK(clknet_leaf_257_clk_i),
    .D(net2717),
    .RESET_B(net262),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _23312_ (.CLK(clknet_leaf_257_clk_i),
    .D(net4271),
    .RESET_B(net262),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _23313_ (.CLK(clknet_leaf_256_clk_i),
    .D(net2742),
    .RESET_B(net262),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _23314_ (.CLK(clknet_leaf_256_clk_i),
    .D(net3130),
    .RESET_B(net262),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _23315_ (.CLK(clknet_leaf_256_clk_i),
    .D(net3797),
    .RESET_B(net264),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _23316_ (.CLK(clknet_leaf_256_clk_i),
    .D(_02587_),
    .RESET_B(net264),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _23317_ (.CLK(clknet_leaf_255_clk_i),
    .D(net2749),
    .RESET_B(net264),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _23318_ (.CLK(clknet_leaf_255_clk_i),
    .D(net2794),
    .RESET_B(net264),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _23319_ (.CLK(clknet_leaf_255_clk_i),
    .D(net2744),
    .RESET_B(net264),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _23320_ (.CLK(clknet_leaf_255_clk_i),
    .D(net2810),
    .RESET_B(net264),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _23321_ (.CLK(clknet_leaf_255_clk_i),
    .D(net3189),
    .RESET_B(net285),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _23322_ (.CLK(clknet_leaf_243_clk_i),
    .D(net2727),
    .RESET_B(net285),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _23323_ (.CLK(clknet_leaf_243_clk_i),
    .D(net2957),
    .RESET_B(net285),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _23324_ (.CLK(clknet_leaf_243_clk_i),
    .D(net2735),
    .RESET_B(net285),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _23325_ (.CLK(clknet_leaf_242_clk_i),
    .D(net2888),
    .RESET_B(net285),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_1 _23326_ (.CLK(clknet_leaf_242_clk_i),
    .D(net2766),
    .RESET_B(net285),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_2 _23327_ (.CLK(clknet_leaf_242_clk_i),
    .D(net4243),
    .RESET_B(net285),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _23328_ (.CLK(clknet_leaf_242_clk_i),
    .D(net2672),
    .RESET_B(net287),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _23329_ (.CLK(clknet_leaf_242_clk_i),
    .D(net2720),
    .RESET_B(net287),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_1 _23330_ (.CLK(clknet_leaf_242_clk_i),
    .D(net4194),
    .RESET_B(net287),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_1 _23331_ (.CLK(clknet_leaf_242_clk_i),
    .D(net4212),
    .RESET_B(net287),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_1 _23332_ (.CLK(clknet_leaf_242_clk_i),
    .D(net4183),
    .RESET_B(net287),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_1 _23333_ (.CLK(clknet_leaf_241_clk_i),
    .D(net4180),
    .RESET_B(net287),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_1 _23334_ (.CLK(clknet_leaf_241_clk_i),
    .D(net4224),
    .RESET_B(net293),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _23335_ (.CLK(clknet_leaf_242_clk_i),
    .D(net4274),
    .RESET_B(net293),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_1 _23336_ (.CLK(clknet_leaf_238_clk_i),
    .D(net4258),
    .RESET_B(net293),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_1 _23337_ (.CLK(clknet_leaf_238_clk_i),
    .D(net4286),
    .RESET_B(net293),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_1 _23338_ (.CLK(clknet_leaf_238_clk_i),
    .D(net2674),
    .RESET_B(net293),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 _23339_ (.CLK(clknet_leaf_238_clk_i),
    .D(_02610_),
    .RESET_B(net293),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_1 _23340_ (.CLK(clknet_leaf_238_clk_i),
    .D(net2841),
    .RESET_B(net294),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_1 _23341_ (.CLK(clknet_leaf_76_clk_i),
    .D(_02612_),
    .RESET_B(net215),
    .Q(\res_v_active[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23342_ (.CLK(clknet_leaf_76_clk_i),
    .D(_02613_),
    .RESET_B(net215),
    .Q(\res_v_active[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23343_ (.CLK(clknet_leaf_76_clk_i),
    .D(_02614_),
    .RESET_B(net215),
    .Q(\res_v_active[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23344_ (.CLK(clknet_leaf_76_clk_i),
    .D(_02615_),
    .RESET_B(net215),
    .Q(\res_v_active[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23345_ (.CLK(clknet_leaf_76_clk_i),
    .D(_02616_),
    .RESET_B(net215),
    .Q(\res_v_active[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23346_ (.CLK(clknet_leaf_75_clk_i),
    .D(_02617_),
    .RESET_B(net215),
    .Q(\res_v_active[5] ));
 sky130_fd_sc_hd__dfrtp_1 _23347_ (.CLK(clknet_leaf_75_clk_i),
    .D(_02618_),
    .RESET_B(net216),
    .Q(\res_v_active[6] ));
 sky130_fd_sc_hd__dfrtp_2 _23348_ (.CLK(clknet_leaf_74_clk_i),
    .D(_02619_),
    .RESET_B(net216),
    .Q(\res_v_active[7] ));
 sky130_fd_sc_hd__dfrtp_2 _23349_ (.CLK(clknet_leaf_60_clk_i),
    .D(_02620_),
    .RESET_B(net166),
    .Q(\base_h_active[0] ));
 sky130_fd_sc_hd__dfrtp_4 _23350_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02621_),
    .RESET_B(net166),
    .Q(\base_h_active[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23351_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02622_),
    .RESET_B(net166),
    .Q(\base_h_active[2] ));
 sky130_fd_sc_hd__dfrtp_4 _23352_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02623_),
    .RESET_B(net166),
    .Q(\base_h_active[3] ));
 sky130_fd_sc_hd__dfrtp_2 _23353_ (.CLK(clknet_leaf_60_clk_i),
    .D(_02624_),
    .RESET_B(net204),
    .Q(\base_h_active[4] ));
 sky130_fd_sc_hd__dfrtp_2 _23354_ (.CLK(clknet_leaf_20_clk_i),
    .D(_02625_),
    .RESET_B(net166),
    .Q(\base_h_active[5] ));
 sky130_fd_sc_hd__dfrtp_4 _23355_ (.CLK(clknet_leaf_59_clk_i),
    .D(_02626_),
    .RESET_B(net204),
    .Q(\base_h_active[6] ));
 sky130_fd_sc_hd__dfrtp_1 _23356_ (.CLK(clknet_leaf_59_clk_i),
    .D(_02627_),
    .RESET_B(net204),
    .Q(\base_h_active[7] ));
 sky130_fd_sc_hd__dfrtp_4 _23357_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02628_),
    .RESET_B(net166),
    .Q(\base_h_active[8] ));
 sky130_fd_sc_hd__dfrtp_2 _23358_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02629_),
    .RESET_B(net166),
    .Q(\base_h_active[9] ));
 sky130_fd_sc_hd__dfrtp_1 _23359_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02630_),
    .RESET_B(net166),
    .Q(\base_h_fporch[0] ));
 sky130_fd_sc_hd__dfrtp_2 _23360_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02631_),
    .RESET_B(net166),
    .Q(\base_h_fporch[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23361_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02632_),
    .RESET_B(net166),
    .Q(\base_h_fporch[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23362_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02633_),
    .RESET_B(net166),
    .Q(\base_h_fporch[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23363_ (.CLK(clknet_leaf_59_clk_i),
    .D(_02634_),
    .RESET_B(net204),
    .Q(\base_h_fporch[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23364_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02635_),
    .RESET_B(net166),
    .Q(\base_h_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23365_ (.CLK(clknet_leaf_61_clk_i),
    .D(_02636_),
    .RESET_B(net204),
    .Q(\base_h_sync[1] ));
 sky130_fd_sc_hd__dfrtp_2 _23366_ (.CLK(clknet_leaf_61_clk_i),
    .D(_02637_),
    .RESET_B(net204),
    .Q(\base_h_sync[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23367_ (.CLK(clknet_leaf_60_clk_i),
    .D(_02638_),
    .RESET_B(net204),
    .Q(\base_h_sync[3] ));
 sky130_fd_sc_hd__dfrtp_2 _23368_ (.CLK(clknet_leaf_60_clk_i),
    .D(_02639_),
    .RESET_B(net204),
    .Q(\base_h_sync[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23369_ (.CLK(clknet_leaf_61_clk_i),
    .D(_02640_),
    .RESET_B(net204),
    .Q(\base_h_sync[5] ));
 sky130_fd_sc_hd__dfrtp_1 _23370_ (.CLK(clknet_leaf_62_clk_i),
    .D(_02641_),
    .RESET_B(net204),
    .Q(\base_h_sync[6] ));
 sky130_fd_sc_hd__dfrtp_1 _23371_ (.CLK(clknet_leaf_63_clk_i),
    .D(_02642_),
    .RESET_B(net206),
    .Q(\base_h_bporch[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23372_ (.CLK(clknet_leaf_61_clk_i),
    .D(_02643_),
    .RESET_B(net204),
    .Q(\base_h_bporch[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23373_ (.CLK(clknet_leaf_63_clk_i),
    .D(_02644_),
    .RESET_B(net206),
    .Q(\base_h_bporch[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23374_ (.CLK(clknet_leaf_63_clk_i),
    .D(_02645_),
    .RESET_B(net206),
    .Q(\base_h_bporch[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23375_ (.CLK(clknet_leaf_63_clk_i),
    .D(_02646_),
    .RESET_B(net206),
    .Q(\base_h_bporch[4] ));
 sky130_fd_sc_hd__dfrtp_2 _23376_ (.CLK(clknet_leaf_64_clk_i),
    .D(_02647_),
    .RESET_B(net206),
    .Q(\base_h_bporch[5] ));
 sky130_fd_sc_hd__dfrtp_2 _23377_ (.CLK(clknet_leaf_64_clk_i),
    .D(_02648_),
    .RESET_B(net206),
    .Q(\base_h_bporch[6] ));
 sky130_fd_sc_hd__dfrtp_2 _23378_ (.CLK(clknet_leaf_78_clk_i),
    .D(_02649_),
    .RESET_B(net215),
    .Q(\base_v_active[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23379_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02650_),
    .RESET_B(net217),
    .Q(\base_v_active[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23380_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02651_),
    .RESET_B(net217),
    .Q(\base_v_active[2] ));
 sky130_fd_sc_hd__dfrtp_2 _23381_ (.CLK(clknet_leaf_76_clk_i),
    .D(_02652_),
    .RESET_B(net215),
    .Q(\base_v_active[3] ));
 sky130_fd_sc_hd__dfrtp_2 _23382_ (.CLK(clknet_leaf_77_clk_i),
    .D(_02653_),
    .RESET_B(net215),
    .Q(\base_v_active[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23383_ (.CLK(clknet_leaf_78_clk_i),
    .D(_02654_),
    .RESET_B(net216),
    .Q(\base_v_active[5] ));
 sky130_fd_sc_hd__dfrtp_2 _23384_ (.CLK(clknet_leaf_79_clk_i),
    .D(_02655_),
    .RESET_B(net216),
    .Q(\base_v_active[6] ));
 sky130_fd_sc_hd__dfrtp_2 _23385_ (.CLK(clknet_leaf_78_clk_i),
    .D(_02656_),
    .RESET_B(net215),
    .Q(\base_v_active[7] ));
 sky130_fd_sc_hd__dfrtp_1 _23386_ (.CLK(clknet_leaf_78_clk_i),
    .D(_02657_),
    .RESET_B(net215),
    .Q(\base_v_active[8] ));
 sky130_fd_sc_hd__dfrtp_1 _23387_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02658_),
    .RESET_B(net217),
    .Q(\base_v_fporch[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23388_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02659_),
    .RESET_B(net217),
    .Q(\base_v_fporch[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23389_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02660_),
    .RESET_B(net217),
    .Q(\base_v_fporch[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23390_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02661_),
    .RESET_B(net217),
    .Q(\base_v_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23391_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02662_),
    .RESET_B(net217),
    .Q(\base_v_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23392_ (.CLK(clknet_leaf_80_clk_i),
    .D(_02663_),
    .RESET_B(net217),
    .Q(\base_v_sync[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23393_ (.CLK(clknet_leaf_81_clk_i),
    .D(_02664_),
    .RESET_B(net217),
    .Q(\base_v_bporch[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23394_ (.CLK(clknet_leaf_81_clk_i),
    .D(_02665_),
    .RESET_B(net217),
    .Q(\base_v_bporch[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23395_ (.CLK(clknet_leaf_81_clk_i),
    .D(_02666_),
    .RESET_B(net217),
    .Q(\base_v_bporch[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23396_ (.CLK(clknet_leaf_81_clk_i),
    .D(_02667_),
    .RESET_B(net217),
    .Q(\base_v_bporch[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23397_ (.CLK(clknet_leaf_2_clk_i),
    .D(_02560_),
    .RESET_B(net150),
    .Q(\prescaler_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23398_ (.CLK(clknet_leaf_2_clk_i),
    .D(_02561_),
    .RESET_B(net151),
    .Q(\prescaler_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23399_ (.CLK(clknet_leaf_3_clk_i),
    .D(_02562_),
    .RESET_B(net151),
    .Q(\prescaler_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23400_ (.CLK(clknet_leaf_13_clk_i),
    .D(_02563_),
    .RESET_B(net162),
    .Q(\prescaler_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23401_ (.CLK(clknet_leaf_13_clk_i),
    .D(_02564_),
    .RESET_B(net162),
    .Q(\prescaler_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23402_ (.CLK(clknet_leaf_13_clk_i),
    .D(_02565_),
    .RESET_B(net162),
    .Q(\prescaler_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _23403_ (.CLK(clknet_leaf_14_clk_i),
    .D(_02566_),
    .RESET_B(net162),
    .Q(\prescaler_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _23404_ (.CLK(clknet_leaf_14_clk_i),
    .D(_02567_),
    .RESET_B(net162),
    .Q(\prescaler_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _23405_ (.CLK(clknet_leaf_14_clk_i),
    .D(net2697),
    .RESET_B(net162),
    .Q(\prescaler_counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _23406_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02668_),
    .RESET_B(net166),
    .Q(\res_h_active[0] ));
 sky130_fd_sc_hd__dfrtp_2 _23407_ (.CLK(clknet_leaf_18_clk_i),
    .D(_02669_),
    .RESET_B(net166),
    .Q(\res_h_active[1] ));
 sky130_fd_sc_hd__dfrtp_2 _23408_ (.CLK(clknet_leaf_18_clk_i),
    .D(_02670_),
    .RESET_B(net167),
    .Q(\res_h_active[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23409_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02671_),
    .RESET_B(net168),
    .Q(\res_h_active[3] ));
 sky130_fd_sc_hd__dfrtp_4 _23410_ (.CLK(clknet_leaf_18_clk_i),
    .D(_02672_),
    .RESET_B(net167),
    .Q(\res_h_active[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23411_ (.CLK(clknet_leaf_16_clk_i),
    .D(_02673_),
    .RESET_B(net168),
    .Q(\res_h_active[5] ));
 sky130_fd_sc_hd__dfrtp_4 _23412_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02674_),
    .RESET_B(net167),
    .Q(\res_h_active[6] ));
 sky130_fd_sc_hd__dfrtp_2 _23413_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02675_),
    .RESET_B(net167),
    .Q(\res_h_active[7] ));
 sky130_fd_sc_hd__dfrtp_2 _23414_ (.CLK(clknet_leaf_18_clk_i),
    .D(_02676_),
    .RESET_B(net167),
    .Q(\res_h_active[8] ));
 sky130_fd_sc_hd__dfrtp_4 _23415_ (.CLK(clknet_leaf_64_clk_i),
    .D(_02677_),
    .RESET_B(net206),
    .Q(\base_h_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23416_ (.CLK(clknet_leaf_62_clk_i),
    .D(net4311),
    .RESET_B(net204),
    .Q(\base_h_counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _23417_ (.CLK(clknet_leaf_60_clk_i),
    .D(_02679_),
    .RESET_B(net166),
    .Q(\base_h_counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _23418_ (.CLK(clknet_leaf_59_clk_i),
    .D(_02680_),
    .RESET_B(net204),
    .Q(\base_h_counter[3] ));
 sky130_fd_sc_hd__dfrtp_4 _23419_ (.CLK(clknet_leaf_62_clk_i),
    .D(net3661),
    .RESET_B(net204),
    .Q(\base_h_counter[4] ));
 sky130_fd_sc_hd__dfrtp_4 _23420_ (.CLK(clknet_leaf_59_clk_i),
    .D(_02682_),
    .RESET_B(net204),
    .Q(\base_h_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _23421_ (.CLK(clknet_leaf_62_clk_i),
    .D(net4267),
    .RESET_B(net204),
    .Q(\base_h_counter[6] ));
 sky130_fd_sc_hd__dfrtp_2 _23422_ (.CLK(clknet_leaf_58_clk_i),
    .D(net3444),
    .RESET_B(net205),
    .Q(\base_h_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _23423_ (.CLK(clknet_leaf_58_clk_i),
    .D(net4152),
    .RESET_B(net205),
    .Q(\base_h_counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _23424_ (.CLK(clknet_leaf_53_clk_i),
    .D(net2897),
    .RESET_B(net206),
    .Q(\base_h_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _23425_ (.CLK(clknet_leaf_77_clk_i),
    .D(net4304),
    .RESET_B(net215),
    .Q(\base_v_counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _23426_ (.CLK(clknet_leaf_77_clk_i),
    .D(net4313),
    .RESET_B(net215),
    .Q(\base_v_counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _23427_ (.CLK(clknet_leaf_78_clk_i),
    .D(net4290),
    .RESET_B(net215),
    .Q(\base_v_counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _23428_ (.CLK(clknet_leaf_79_clk_i),
    .D(net4301),
    .RESET_B(net216),
    .Q(\base_v_counter[3] ));
 sky130_fd_sc_hd__dfrtp_4 _23429_ (.CLK(clknet_leaf_79_clk_i),
    .D(net4307),
    .RESET_B(net216),
    .Q(\base_v_counter[4] ));
 sky130_fd_sc_hd__dfrtp_4 _23430_ (.CLK(clknet_leaf_73_clk_i),
    .D(_02692_),
    .RESET_B(net216),
    .Q(\base_v_counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _23431_ (.CLK(clknet_leaf_79_clk_i),
    .D(net4299),
    .RESET_B(net216),
    .Q(\base_v_counter[6] ));
 sky130_fd_sc_hd__dfrtp_4 _23432_ (.CLK(clknet_leaf_73_clk_i),
    .D(_02694_),
    .RESET_B(net218),
    .Q(\base_v_counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _23433_ (.CLK(clknet_leaf_73_clk_i),
    .D(_02695_),
    .RESET_B(net218),
    .Q(\base_v_counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _23434_ (.CLK(clknet_leaf_73_clk_i),
    .D(net4230),
    .RESET_B(net216),
    .Q(\base_v_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _23435_ (.CLK(clknet_leaf_22_clk_i),
    .D(net2771),
    .RESET_B(net172),
    .Q(\res_h_counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _23436_ (.CLK(clknet_leaf_22_clk_i),
    .D(net3039),
    .RESET_B(net172),
    .Q(\res_h_counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _23437_ (.CLK(clknet_leaf_22_clk_i),
    .D(net3920),
    .RESET_B(net172),
    .Q(\res_h_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23438_ (.CLK(clknet_leaf_23_clk_i),
    .D(net2786),
    .RESET_B(net173),
    .Q(\res_h_counter[3] ));
 sky130_fd_sc_hd__dfrtp_4 _23439_ (.CLK(clknet_leaf_24_clk_i),
    .D(_02701_),
    .RESET_B(net173),
    .Q(\res_h_counter[4] ));
 sky130_fd_sc_hd__dfrtp_4 _23440_ (.CLK(clknet_leaf_24_clk_i),
    .D(net4187),
    .RESET_B(net173),
    .Q(\res_h_counter[5] ));
 sky130_fd_sc_hd__dfrtp_4 _23441_ (.CLK(clknet_leaf_23_clk_i),
    .D(net2751),
    .RESET_B(net173),
    .Q(\res_h_counter[6] ));
 sky130_fd_sc_hd__dfrtp_4 _23442_ (.CLK(clknet_leaf_22_clk_i),
    .D(net3653),
    .RESET_B(net173),
    .Q(\res_h_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _23443_ (.CLK(clknet_leaf_23_clk_i),
    .D(_02705_),
    .RESET_B(net173),
    .Q(\res_h_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _23444_ (.CLK(clknet_leaf_22_clk_i),
    .D(net1860),
    .RESET_B(net172),
    .Q(\res_h_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _23445_ (.CLK(clknet_leaf_64_clk_i),
    .D(net2959),
    .RESET_B(net206),
    .Q(\res_v_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23446_ (.CLK(clknet_leaf_64_clk_i),
    .D(net2779),
    .RESET_B(net206),
    .Q(\res_v_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23447_ (.CLK(clknet_leaf_64_clk_i),
    .D(net2693),
    .RESET_B(net206),
    .Q(\res_v_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23448_ (.CLK(clknet_leaf_75_clk_i),
    .D(net2827),
    .RESET_B(net215),
    .Q(\res_v_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23449_ (.CLK(clknet_leaf_74_clk_i),
    .D(net3518),
    .RESET_B(net215),
    .Q(\res_v_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _23450_ (.CLK(clknet_leaf_64_clk_i),
    .D(net3019),
    .RESET_B(net206),
    .Q(\res_v_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _23451_ (.CLK(clknet_leaf_74_clk_i),
    .D(net2670),
    .RESET_B(net216),
    .Q(\res_v_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _23452_ (.CLK(clknet_leaf_74_clk_i),
    .D(net2730),
    .RESET_B(net216),
    .Q(\res_v_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _23453_ (.CLK(clknet_leaf_65_clk_i),
    .D(net2686),
    .RESET_B(net206),
    .Q(\res_v_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _23454_ (.CLK(clknet_leaf_65_clk_i),
    .D(net2689),
    .RESET_B(net206),
    .Q(\res_v_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _23455_ (.CLK(clknet_leaf_1_clk_i),
    .D(_02717_),
    .RESET_B(net150),
    .Q(\prescaler[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23456_ (.CLK(clknet_leaf_1_clk_i),
    .D(_02718_),
    .RESET_B(net150),
    .Q(\prescaler[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23457_ (.CLK(clknet_leaf_1_clk_i),
    .D(_02719_),
    .RESET_B(net150),
    .Q(\prescaler[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23458_ (.CLK(clknet_leaf_1_clk_i),
    .D(_02720_),
    .RESET_B(net150),
    .Q(\prescaler[3] ));
 sky130_fd_sc_hd__dfrtp_4 _23459_ (.CLK(clknet_leaf_18_clk_i),
    .D(_02721_),
    .RESET_B(net167),
    .Q(\resolution[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23460_ (.CLK(clknet_leaf_18_clk_i),
    .D(_02722_),
    .RESET_B(net167),
    .Q(\resolution[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23461_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02723_),
    .RESET_B(net168),
    .Q(\resolution[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23462_ (.CLK(clknet_leaf_18_clk_i),
    .D(_02724_),
    .RESET_B(net167),
    .Q(\resolution[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23463_ (.CLK(clknet_leaf_59_clk_i),
    .D(net2649),
    .RESET_B(net205),
    .Q(\pixel_double_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23464_ (.CLK(clknet_leaf_59_clk_i),
    .D(net2656),
    .RESET_B(net205),
    .Q(\pixel_double_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23465_ (.CLK(clknet_leaf_59_clk_i),
    .D(net1914),
    .RESET_B(net205),
    .Q(\pixel_double_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23466_ (.CLK(clknet_leaf_57_clk_i),
    .D(net1878),
    .RESET_B(net168),
    .Q(\pixel_double_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23467_ (.CLK(clknet_leaf_19_clk_i),
    .D(_02729_),
    .RESET_B(net166),
    .Q(\line_double_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _23468_ (.CLK(clknet_leaf_20_clk_i),
    .D(net2662),
    .RESET_B(net168),
    .Q(\line_double_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _23469_ (.CLK(clknet_leaf_19_clk_i),
    .D(net2679),
    .RESET_B(net167),
    .Q(\line_double_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _23470_ (.CLK(clknet_leaf_20_clk_i),
    .D(net2682),
    .RESET_B(net168),
    .Q(\line_double_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _23471_ (.CLK(clknet_leaf_290_clk_i),
    .D(net608),
    .RESET_B(net196),
    .Q(\line_cache[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23472_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00001_),
    .RESET_B(net191),
    .Q(\line_cache[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23473_ (.CLK(clknet_leaf_290_clk_i),
    .D(net1746),
    .RESET_B(net196),
    .Q(\line_cache[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23474_ (.CLK(clknet_leaf_290_clk_i),
    .D(net2548),
    .RESET_B(net196),
    .Q(\line_cache[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23475_ (.CLK(clknet_leaf_290_clk_i),
    .D(net696),
    .RESET_B(net196),
    .Q(\line_cache[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23476_ (.CLK(clknet_leaf_289_clk_i),
    .D(_00005_),
    .RESET_B(net197),
    .Q(\line_cache[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23477_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00006_),
    .RESET_B(net191),
    .Q(\line_cache[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23478_ (.CLK(clknet_leaf_30_clk_i),
    .D(net4296),
    .RESET_B(net191),
    .Q(\line_cache[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23479_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00888_),
    .RESET_B(net190),
    .Q(\line_cache[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23480_ (.CLK(clknet_leaf_30_clk_i),
    .D(net648),
    .RESET_B(net191),
    .Q(\line_cache[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23481_ (.CLK(clknet_leaf_30_clk_i),
    .D(net472),
    .RESET_B(net190),
    .Q(\line_cache[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23482_ (.CLK(clknet_leaf_294_clk_i),
    .D(net1360),
    .RESET_B(net191),
    .Q(\line_cache[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23483_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00892_),
    .RESET_B(net179),
    .Q(\line_cache[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23484_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00893_),
    .RESET_B(net190),
    .Q(\line_cache[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23485_ (.CLK(clknet_leaf_295_clk_i),
    .D(_00894_),
    .RESET_B(net191),
    .Q(\line_cache[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23486_ (.CLK(clknet_leaf_295_clk_i),
    .D(_00895_),
    .RESET_B(net191),
    .Q(\line_cache[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23487_ (.CLK(clknet_leaf_29_clk_i),
    .D(net444),
    .RESET_B(net190),
    .Q(\line_cache[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23488_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01777_),
    .RESET_B(net190),
    .Q(\line_cache[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23489_ (.CLK(clknet_leaf_29_clk_i),
    .D(_01778_),
    .RESET_B(net190),
    .Q(\line_cache[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23490_ (.CLK(clknet_leaf_295_clk_i),
    .D(net506),
    .RESET_B(net191),
    .Q(\line_cache[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23491_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01780_),
    .RESET_B(net190),
    .Q(\line_cache[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23492_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01781_),
    .RESET_B(net190),
    .Q(\line_cache[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23493_ (.CLK(clknet_leaf_29_clk_i),
    .D(_01782_),
    .RESET_B(net190),
    .Q(\line_cache[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23494_ (.CLK(clknet_leaf_30_clk_i),
    .D(net810),
    .RESET_B(net191),
    .Q(\line_cache[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23495_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02024_),
    .RESET_B(net190),
    .Q(\line_cache[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23496_ (.CLK(clknet_leaf_26_clk_i),
    .D(net766),
    .RESET_B(net170),
    .Q(\line_cache[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23497_ (.CLK(clknet_leaf_26_clk_i),
    .D(net492),
    .RESET_B(net170),
    .Q(\line_cache[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23498_ (.CLK(clknet_leaf_26_clk_i),
    .D(net930),
    .RESET_B(net170),
    .Q(\line_cache[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23499_ (.CLK(clknet_leaf_26_clk_i),
    .D(net1666),
    .RESET_B(net170),
    .Q(\line_cache[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23500_ (.CLK(clknet_leaf_26_clk_i),
    .D(net850),
    .RESET_B(net171),
    .Q(\line_cache[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23501_ (.CLK(clknet_leaf_29_clk_i),
    .D(net532),
    .RESET_B(net192),
    .Q(\line_cache[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23502_ (.CLK(clknet_leaf_29_clk_i),
    .D(net624),
    .RESET_B(net192),
    .Q(\line_cache[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23503_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02112_),
    .RESET_B(net192),
    .Q(\line_cache[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23504_ (.CLK(clknet_leaf_26_clk_i),
    .D(_02113_),
    .RESET_B(net171),
    .Q(\line_cache[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23505_ (.CLK(clknet_leaf_24_clk_i),
    .D(_02114_),
    .RESET_B(net173),
    .Q(\line_cache[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23506_ (.CLK(clknet_leaf_27_clk_i),
    .D(_02115_),
    .RESET_B(net170),
    .Q(\line_cache[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23507_ (.CLK(clknet_leaf_25_clk_i),
    .D(_02116_),
    .RESET_B(net171),
    .Q(\line_cache[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23508_ (.CLK(clknet_leaf_27_clk_i),
    .D(_02117_),
    .RESET_B(net170),
    .Q(\line_cache[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23509_ (.CLK(clknet_leaf_27_clk_i),
    .D(_02118_),
    .RESET_B(net170),
    .Q(\line_cache[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23510_ (.CLK(clknet_leaf_26_clk_i),
    .D(_02119_),
    .RESET_B(net171),
    .Q(\line_cache[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23511_ (.CLK(clknet_leaf_26_clk_i),
    .D(_02200_),
    .RESET_B(net171),
    .Q(\line_cache[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23512_ (.CLK(clknet_leaf_27_clk_i),
    .D(_02201_),
    .RESET_B(net170),
    .Q(\line_cache[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23513_ (.CLK(clknet_leaf_26_clk_i),
    .D(_02202_),
    .RESET_B(net171),
    .Q(\line_cache[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23514_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02203_),
    .RESET_B(net170),
    .Q(\line_cache[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23515_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02204_),
    .RESET_B(net170),
    .Q(\line_cache[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23516_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02205_),
    .RESET_B(net170),
    .Q(\line_cache[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23517_ (.CLK(clknet_leaf_28_clk_i),
    .D(_02206_),
    .RESET_B(net190),
    .Q(\line_cache[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23518_ (.CLK(clknet_leaf_28_clk_i),
    .D(_02207_),
    .RESET_B(net190),
    .Q(\line_cache[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23519_ (.CLK(clknet_leaf_25_clk_i),
    .D(_02288_),
    .RESET_B(net169),
    .Q(\line_cache[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23520_ (.CLK(clknet_leaf_10_clk_i),
    .D(_02289_),
    .RESET_B(net169),
    .Q(\line_cache[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23521_ (.CLK(clknet_leaf_24_clk_i),
    .D(_02290_),
    .RESET_B(net172),
    .Q(\line_cache[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23522_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02291_),
    .RESET_B(net169),
    .Q(\line_cache[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23523_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02292_),
    .RESET_B(net170),
    .Q(\line_cache[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23524_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02293_),
    .RESET_B(net170),
    .Q(\line_cache[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23525_ (.CLK(clknet_leaf_27_clk_i),
    .D(_02294_),
    .RESET_B(net170),
    .Q(\line_cache[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23526_ (.CLK(clknet_leaf_27_clk_i),
    .D(_02295_),
    .RESET_B(net170),
    .Q(\line_cache[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23527_ (.CLK(clknet_leaf_25_clk_i),
    .D(_02376_),
    .RESET_B(net169),
    .Q(\line_cache[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23528_ (.CLK(clknet_leaf_16_clk_i),
    .D(_02377_),
    .RESET_B(net164),
    .Q(\line_cache[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23529_ (.CLK(clknet_leaf_16_clk_i),
    .D(_02378_),
    .RESET_B(net164),
    .Q(\line_cache[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23530_ (.CLK(clknet_leaf_15_clk_i),
    .D(_02379_),
    .RESET_B(net163),
    .Q(\line_cache[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23531_ (.CLK(clknet_leaf_11_clk_i),
    .D(_02380_),
    .RESET_B(net169),
    .Q(\line_cache[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23532_ (.CLK(clknet_leaf_15_clk_i),
    .D(_02381_),
    .RESET_B(net163),
    .Q(\line_cache[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23533_ (.CLK(clknet_leaf_26_clk_i),
    .D(_02382_),
    .RESET_B(net169),
    .Q(\line_cache[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23534_ (.CLK(clknet_leaf_15_clk_i),
    .D(_02383_),
    .RESET_B(net163),
    .Q(\line_cache[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23535_ (.CLK(clknet_leaf_21_clk_i),
    .D(_02464_),
    .RESET_B(net172),
    .Q(\line_cache[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23536_ (.CLK(clknet_leaf_11_clk_i),
    .D(net1958),
    .RESET_B(net164),
    .Q(\line_cache[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23537_ (.CLK(clknet_leaf_16_clk_i),
    .D(_02466_),
    .RESET_B(net164),
    .Q(\line_cache[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23538_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02467_),
    .RESET_B(net167),
    .Q(\line_cache[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23539_ (.CLK(clknet_leaf_25_clk_i),
    .D(_02468_),
    .RESET_B(net169),
    .Q(\line_cache[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23540_ (.CLK(clknet_leaf_11_clk_i),
    .D(net4106),
    .RESET_B(net165),
    .Q(\line_cache[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23541_ (.CLK(clknet_leaf_25_clk_i),
    .D(net4018),
    .RESET_B(net171),
    .Q(\line_cache[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23542_ (.CLK(clknet_leaf_16_clk_i),
    .D(net1677),
    .RESET_B(net165),
    .Q(\line_cache[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23543_ (.CLK(clknet_leaf_21_clk_i),
    .D(_02552_),
    .RESET_B(net168),
    .Q(\line_cache[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23544_ (.CLK(clknet_leaf_16_clk_i),
    .D(net1873),
    .RESET_B(net165),
    .Q(\line_cache[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23545_ (.CLK(clknet_leaf_16_clk_i),
    .D(net958),
    .RESET_B(net165),
    .Q(\line_cache[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23546_ (.CLK(clknet_leaf_15_clk_i),
    .D(_02555_),
    .RESET_B(net163),
    .Q(\line_cache[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23547_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02556_),
    .RESET_B(net167),
    .Q(\line_cache[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23548_ (.CLK(clknet_leaf_17_clk_i),
    .D(_02557_),
    .RESET_B(net167),
    .Q(\line_cache[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23549_ (.CLK(clknet_leaf_25_clk_i),
    .D(net1068),
    .RESET_B(net172),
    .Q(\line_cache[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23550_ (.CLK(clknet_leaf_15_clk_i),
    .D(_02559_),
    .RESET_B(net163),
    .Q(\line_cache[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23551_ (.CLK(clknet_leaf_16_clk_i),
    .D(net1108),
    .RESET_B(net168),
    .Q(\line_cache[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23552_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00089_),
    .RESET_B(net168),
    .Q(\line_cache[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23553_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00090_),
    .RESET_B(net168),
    .Q(\line_cache[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23554_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00091_),
    .RESET_B(net163),
    .Q(\line_cache[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23555_ (.CLK(clknet_leaf_21_clk_i),
    .D(net640),
    .RESET_B(net168),
    .Q(\line_cache[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23556_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00093_),
    .RESET_B(net163),
    .Q(\line_cache[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23557_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00094_),
    .RESET_B(net171),
    .Q(\line_cache[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23558_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00095_),
    .RESET_B(net163),
    .Q(\line_cache[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23559_ (.CLK(clknet_leaf_10_clk_i),
    .D(net864),
    .RESET_B(net171),
    .Q(\line_cache[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23560_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00177_),
    .RESET_B(net164),
    .Q(\line_cache[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23561_ (.CLK(clknet_leaf_11_clk_i),
    .D(net1545),
    .RESET_B(net165),
    .Q(\line_cache[11][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23562_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00179_),
    .RESET_B(net164),
    .Q(\line_cache[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23563_ (.CLK(clknet_leaf_10_clk_i),
    .D(net1732),
    .RESET_B(net169),
    .Q(\line_cache[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23564_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00181_),
    .RESET_B(net163),
    .Q(\line_cache[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23565_ (.CLK(clknet_leaf_10_clk_i),
    .D(net1188),
    .RESET_B(net169),
    .Q(\line_cache[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23566_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00183_),
    .RESET_B(net163),
    .Q(\line_cache[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23567_ (.CLK(clknet_leaf_10_clk_i),
    .D(net1588),
    .RESET_B(net171),
    .Q(\line_cache[12][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23568_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00265_),
    .RESET_B(net164),
    .Q(\line_cache[12][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23569_ (.CLK(clknet_leaf_11_clk_i),
    .D(net1220),
    .RESET_B(net164),
    .Q(\line_cache[12][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23570_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00267_),
    .RESET_B(net162),
    .Q(\line_cache[12][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23571_ (.CLK(clknet_leaf_11_clk_i),
    .D(net618),
    .RESET_B(net164),
    .Q(\line_cache[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23572_ (.CLK(clknet_leaf_11_clk_i),
    .D(net836),
    .RESET_B(net165),
    .Q(\line_cache[12][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23573_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00270_),
    .RESET_B(net169),
    .Q(\line_cache[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23574_ (.CLK(clknet_leaf_14_clk_i),
    .D(net518),
    .RESET_B(net162),
    .Q(\line_cache[12][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23575_ (.CLK(clknet_leaf_11_clk_i),
    .D(net1833),
    .RESET_B(net171),
    .Q(\line_cache[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23576_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00353_),
    .RESET_B(net164),
    .Q(\line_cache[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23577_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00354_),
    .RESET_B(net162),
    .Q(\line_cache[13][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23578_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00355_),
    .RESET_B(net162),
    .Q(\line_cache[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23579_ (.CLK(clknet_leaf_11_clk_i),
    .D(net1488),
    .RESET_B(net164),
    .Q(\line_cache[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23580_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00357_),
    .RESET_B(net163),
    .Q(\line_cache[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23581_ (.CLK(clknet_leaf_10_clk_i),
    .D(net1785),
    .RESET_B(net169),
    .Q(\line_cache[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23582_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00359_),
    .RESET_B(net162),
    .Q(\line_cache[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23583_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00440_),
    .RESET_B(net164),
    .Q(\line_cache[14][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23584_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00441_),
    .RESET_B(net164),
    .Q(\line_cache[14][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23585_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00442_),
    .RESET_B(net162),
    .Q(\line_cache[14][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23586_ (.CLK(clknet_leaf_12_clk_i),
    .D(net2194),
    .RESET_B(net162),
    .Q(\line_cache[14][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23587_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00444_),
    .RESET_B(net164),
    .Q(\line_cache[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23588_ (.CLK(clknet_leaf_11_clk_i),
    .D(net1865),
    .RESET_B(net165),
    .Q(\line_cache[14][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23589_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00446_),
    .RESET_B(net169),
    .Q(\line_cache[14][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23590_ (.CLK(clknet_leaf_14_clk_i),
    .D(net1538),
    .RESET_B(net162),
    .Q(\line_cache[14][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23591_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00528_),
    .RESET_B(net171),
    .Q(\line_cache[15][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23592_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00529_),
    .RESET_B(net192),
    .Q(\line_cache[15][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23593_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00530_),
    .RESET_B(net192),
    .Q(\line_cache[15][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23594_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00531_),
    .RESET_B(net190),
    .Q(\line_cache[15][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23595_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00532_),
    .RESET_B(net190),
    .Q(\line_cache[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23596_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00533_),
    .RESET_B(net190),
    .Q(\line_cache[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23597_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00534_),
    .RESET_B(net169),
    .Q(\line_cache[15][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23598_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00535_),
    .RESET_B(net190),
    .Q(\line_cache[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23599_ (.CLK(clknet_leaf_332_clk_i),
    .D(net2138),
    .RESET_B(net148),
    .Q(\line_cache[16][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23600_ (.CLK(clknet_leaf_331_clk_i),
    .D(net1490),
    .RESET_B(net147),
    .Q(\line_cache[16][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23601_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00618_),
    .RESET_B(net147),
    .Q(\line_cache[16][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23602_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00619_),
    .RESET_B(net147),
    .Q(\line_cache[16][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23603_ (.CLK(clknet_leaf_332_clk_i),
    .D(net2519),
    .RESET_B(net148),
    .Q(\line_cache[16][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23604_ (.CLK(clknet_leaf_0_clk_i),
    .D(net2501),
    .RESET_B(net150),
    .Q(\line_cache[16][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23605_ (.CLK(clknet_leaf_332_clk_i),
    .D(net3515),
    .RESET_B(net149),
    .Q(\line_cache[16][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23606_ (.CLK(clknet_leaf_332_clk_i),
    .D(net3961),
    .RESET_B(net149),
    .Q(\line_cache[16][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23607_ (.CLK(clknet_leaf_0_clk_i),
    .D(net1748),
    .RESET_B(net149),
    .Q(\line_cache[17][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23608_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00705_),
    .RESET_B(net147),
    .Q(\line_cache[17][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23609_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00706_),
    .RESET_B(net147),
    .Q(\line_cache[17][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23610_ (.CLK(clknet_leaf_331_clk_i),
    .D(net1880),
    .RESET_B(net147),
    .Q(\line_cache[17][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23611_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00708_),
    .RESET_B(net147),
    .Q(\line_cache[17][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23612_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00709_),
    .RESET_B(net147),
    .Q(\line_cache[17][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23613_ (.CLK(clknet_leaf_332_clk_i),
    .D(_00710_),
    .RESET_B(net149),
    .Q(\line_cache[17][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23614_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00711_),
    .RESET_B(net147),
    .Q(\line_cache[17][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23615_ (.CLK(clknet_leaf_0_clk_i),
    .D(net1632),
    .RESET_B(net152),
    .Q(\line_cache[18][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23616_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00793_),
    .RESET_B(net147),
    .Q(\line_cache[18][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23617_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00794_),
    .RESET_B(net147),
    .Q(\line_cache[18][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23618_ (.CLK(clknet_leaf_330_clk_i),
    .D(net1258),
    .RESET_B(net148),
    .Q(\line_cache[18][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23619_ (.CLK(clknet_leaf_328_clk_i),
    .D(net1050),
    .RESET_B(net149),
    .Q(\line_cache[18][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23620_ (.CLK(clknet_leaf_0_clk_i),
    .D(net2153),
    .RESET_B(net150),
    .Q(\line_cache[18][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23621_ (.CLK(clknet_leaf_327_clk_i),
    .D(net1980),
    .RESET_B(net149),
    .Q(\line_cache[18][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23622_ (.CLK(clknet_leaf_331_clk_i),
    .D(net1266),
    .RESET_B(net154),
    .Q(\line_cache[18][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23623_ (.CLK(clknet_leaf_321_clk_i),
    .D(net758),
    .RESET_B(net152),
    .Q(\line_cache[19][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23624_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00881_),
    .RESET_B(net147),
    .Q(\line_cache[19][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23625_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00882_),
    .RESET_B(net147),
    .Q(\line_cache[19][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23626_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00883_),
    .RESET_B(net147),
    .Q(\line_cache[19][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23627_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00884_),
    .RESET_B(net154),
    .Q(\line_cache[19][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23628_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00885_),
    .RESET_B(net150),
    .Q(\line_cache[19][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23629_ (.CLK(clknet_leaf_327_clk_i),
    .D(_00886_),
    .RESET_B(net149),
    .Q(\line_cache[19][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23630_ (.CLK(clknet_leaf_331_clk_i),
    .D(_00887_),
    .RESET_B(net154),
    .Q(\line_cache[19][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23631_ (.CLK(clknet_leaf_326_clk_i),
    .D(net2482),
    .RESET_B(net155),
    .Q(\line_cache[20][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23632_ (.CLK(clknet_leaf_329_clk_i),
    .D(net1923),
    .RESET_B(net148),
    .Q(\line_cache[20][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23633_ (.CLK(clknet_leaf_327_clk_i),
    .D(net634),
    .RESET_B(net149),
    .Q(\line_cache[20][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23634_ (.CLK(clknet_leaf_330_clk_i),
    .D(_00979_),
    .RESET_B(net147),
    .Q(\line_cache[20][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23635_ (.CLK(clknet_leaf_327_clk_i),
    .D(net678),
    .RESET_B(net155),
    .Q(\line_cache[20][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23636_ (.CLK(clknet_leaf_321_clk_i),
    .D(_00981_),
    .RESET_B(net155),
    .Q(\line_cache[20][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23637_ (.CLK(clknet_leaf_327_clk_i),
    .D(_00982_),
    .RESET_B(net156),
    .Q(\line_cache[20][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23638_ (.CLK(clknet_leaf_327_clk_i),
    .D(_00983_),
    .RESET_B(net149),
    .Q(\line_cache[20][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23639_ (.CLK(clknet_leaf_326_clk_i),
    .D(_01064_),
    .RESET_B(net155),
    .Q(\line_cache[21][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23640_ (.CLK(clknet_leaf_329_clk_i),
    .D(net2318),
    .RESET_B(net148),
    .Q(\line_cache[21][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23641_ (.CLK(clknet_leaf_328_clk_i),
    .D(net434),
    .RESET_B(net148),
    .Q(\line_cache[21][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23642_ (.CLK(clknet_leaf_329_clk_i),
    .D(net2407),
    .RESET_B(net148),
    .Q(\line_cache[21][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23643_ (.CLK(clknet_leaf_326_clk_i),
    .D(net888),
    .RESET_B(net155),
    .Q(\line_cache[21][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23644_ (.CLK(clknet_leaf_327_clk_i),
    .D(_01069_),
    .RESET_B(net149),
    .Q(\line_cache[21][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23645_ (.CLK(clknet_leaf_327_clk_i),
    .D(_01070_),
    .RESET_B(net156),
    .Q(\line_cache[21][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23646_ (.CLK(clknet_leaf_330_clk_i),
    .D(_01071_),
    .RESET_B(net147),
    .Q(\line_cache[21][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23647_ (.CLK(clknet_leaf_326_clk_i),
    .D(_01152_),
    .RESET_B(net155),
    .Q(\line_cache[22][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23648_ (.CLK(clknet_leaf_329_clk_i),
    .D(_01153_),
    .RESET_B(net148),
    .Q(\line_cache[22][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23649_ (.CLK(clknet_leaf_329_clk_i),
    .D(_01154_),
    .RESET_B(net148),
    .Q(\line_cache[22][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23650_ (.CLK(clknet_leaf_329_clk_i),
    .D(net2063),
    .RESET_B(net148),
    .Q(\line_cache[22][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23651_ (.CLK(clknet_leaf_328_clk_i),
    .D(net1206),
    .RESET_B(net148),
    .Q(\line_cache[22][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23652_ (.CLK(clknet_leaf_326_clk_i),
    .D(_01157_),
    .RESET_B(net155),
    .Q(\line_cache[22][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23653_ (.CLK(clknet_leaf_326_clk_i),
    .D(net2447),
    .RESET_B(net155),
    .Q(\line_cache[22][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23654_ (.CLK(clknet_leaf_329_clk_i),
    .D(_01159_),
    .RESET_B(net148),
    .Q(\line_cache[22][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23655_ (.CLK(clknet_leaf_326_clk_i),
    .D(net1893),
    .RESET_B(net155),
    .Q(\line_cache[23][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23656_ (.CLK(clknet_leaf_329_clk_i),
    .D(net1598),
    .RESET_B(net148),
    .Q(\line_cache[23][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23657_ (.CLK(clknet_leaf_329_clk_i),
    .D(net1326),
    .RESET_B(net148),
    .Q(\line_cache[23][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23658_ (.CLK(clknet_leaf_329_clk_i),
    .D(net1992),
    .RESET_B(net148),
    .Q(\line_cache[23][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23659_ (.CLK(clknet_leaf_328_clk_i),
    .D(_01244_),
    .RESET_B(net148),
    .Q(\line_cache[23][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23660_ (.CLK(clknet_leaf_326_clk_i),
    .D(net2573),
    .RESET_B(net155),
    .Q(\line_cache[23][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23661_ (.CLK(clknet_leaf_326_clk_i),
    .D(_01246_),
    .RESET_B(net155),
    .Q(\line_cache[23][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23662_ (.CLK(clknet_leaf_326_clk_i),
    .D(net2641),
    .RESET_B(net155),
    .Q(\line_cache[23][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23663_ (.CLK(clknet_leaf_326_clk_i),
    .D(net1386),
    .RESET_B(net156),
    .Q(\line_cache[24][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23664_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01329_),
    .RESET_B(net157),
    .Q(\line_cache[24][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23665_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01330_),
    .RESET_B(net157),
    .Q(\line_cache[24][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23666_ (.CLK(clknet_leaf_312_clk_i),
    .D(_01331_),
    .RESET_B(net157),
    .Q(\line_cache[24][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23667_ (.CLK(clknet_leaf_327_clk_i),
    .D(net1520),
    .RESET_B(net156),
    .Q(\line_cache[24][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23668_ (.CLK(clknet_leaf_322_clk_i),
    .D(net3790),
    .RESET_B(net157),
    .Q(\line_cache[24][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23669_ (.CLK(clknet_leaf_322_clk_i),
    .D(net3588),
    .RESET_B(net156),
    .Q(\line_cache[24][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23670_ (.CLK(clknet_leaf_323_clk_i),
    .D(net3805),
    .RESET_B(net157),
    .Q(\line_cache[24][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23671_ (.CLK(clknet_leaf_326_clk_i),
    .D(net808),
    .RESET_B(net155),
    .Q(\line_cache[25][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23672_ (.CLK(clknet_leaf_323_clk_i),
    .D(net1122),
    .RESET_B(net158),
    .Q(\line_cache[25][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23673_ (.CLK(clknet_leaf_326_clk_i),
    .D(net1843),
    .RESET_B(net155),
    .Q(\line_cache[25][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23674_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01419_),
    .RESET_B(net157),
    .Q(\line_cache[25][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23675_ (.CLK(clknet_leaf_322_clk_i),
    .D(net460),
    .RESET_B(net156),
    .Q(\line_cache[25][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23676_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01421_),
    .RESET_B(net157),
    .Q(\line_cache[25][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23677_ (.CLK(clknet_leaf_321_clk_i),
    .D(net784),
    .RESET_B(net156),
    .Q(\line_cache[25][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23678_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01423_),
    .RESET_B(net157),
    .Q(\line_cache[25][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23679_ (.CLK(clknet_leaf_326_clk_i),
    .D(_01504_),
    .RESET_B(net155),
    .Q(\line_cache[26][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23680_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01505_),
    .RESET_B(net157),
    .Q(\line_cache[26][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23681_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01506_),
    .RESET_B(net157),
    .Q(\line_cache[26][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23682_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01507_),
    .RESET_B(net157),
    .Q(\line_cache[26][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23683_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01508_),
    .RESET_B(net156),
    .Q(\line_cache[26][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23684_ (.CLK(clknet_leaf_322_clk_i),
    .D(_01509_),
    .RESET_B(net158),
    .Q(\line_cache[26][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23685_ (.CLK(clknet_leaf_321_clk_i),
    .D(net1730),
    .RESET_B(net156),
    .Q(\line_cache[26][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23686_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01511_),
    .RESET_B(net158),
    .Q(\line_cache[26][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23687_ (.CLK(clknet_leaf_326_clk_i),
    .D(_01592_),
    .RESET_B(net155),
    .Q(\line_cache[27][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23688_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01593_),
    .RESET_B(net157),
    .Q(\line_cache[27][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23689_ (.CLK(clknet_leaf_325_clk_i),
    .D(_01594_),
    .RESET_B(net157),
    .Q(\line_cache[27][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23690_ (.CLK(clknet_leaf_324_clk_i),
    .D(_01595_),
    .RESET_B(net157),
    .Q(\line_cache[27][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23691_ (.CLK(clknet_leaf_321_clk_i),
    .D(net2564),
    .RESET_B(net156),
    .Q(\line_cache[27][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23692_ (.CLK(clknet_leaf_322_clk_i),
    .D(net2606),
    .RESET_B(net158),
    .Q(\line_cache[27][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23693_ (.CLK(clknet_leaf_322_clk_i),
    .D(net1681),
    .RESET_B(net156),
    .Q(\line_cache[27][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23694_ (.CLK(clknet_leaf_323_clk_i),
    .D(_01599_),
    .RESET_B(net158),
    .Q(\line_cache[27][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23695_ (.CLK(clknet_leaf_318_clk_i),
    .D(net616),
    .RESET_B(net160),
    .Q(\line_cache[28][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23696_ (.CLK(clknet_leaf_319_clk_i),
    .D(_01681_),
    .RESET_B(net160),
    .Q(\line_cache[28][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23697_ (.CLK(clknet_leaf_318_clk_i),
    .D(net1781),
    .RESET_B(net160),
    .Q(\line_cache[28][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23698_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01683_),
    .RESET_B(net160),
    .Q(\line_cache[28][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23699_ (.CLK(clknet_leaf_316_clk_i),
    .D(net1464),
    .RESET_B(net160),
    .Q(\line_cache[28][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23700_ (.CLK(clknet_leaf_318_clk_i),
    .D(net1672),
    .RESET_B(net160),
    .Q(\line_cache[28][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23701_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01686_),
    .RESET_B(net160),
    .Q(\line_cache[28][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23702_ (.CLK(clknet_leaf_319_clk_i),
    .D(net1646),
    .RESET_B(net160),
    .Q(\line_cache[28][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23703_ (.CLK(clknet_leaf_319_clk_i),
    .D(net1430),
    .RESET_B(net160),
    .Q(\line_cache[29][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23704_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01769_),
    .RESET_B(net160),
    .Q(\line_cache[29][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23705_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01770_),
    .RESET_B(net160),
    .Q(\line_cache[29][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23706_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01771_),
    .RESET_B(net160),
    .Q(\line_cache[29][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23707_ (.CLK(clknet_leaf_319_clk_i),
    .D(net800),
    .RESET_B(net160),
    .Q(\line_cache[29][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23708_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01773_),
    .RESET_B(net179),
    .Q(\line_cache[29][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23709_ (.CLK(clknet_leaf_317_clk_i),
    .D(net1374),
    .RESET_B(net179),
    .Q(\line_cache[29][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23710_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01775_),
    .RESET_B(net160),
    .Q(\line_cache[29][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23711_ (.CLK(clknet_leaf_320_clk_i),
    .D(net498),
    .RESET_B(net160),
    .Q(\line_cache[30][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23712_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01865_),
    .RESET_B(net161),
    .Q(\line_cache[30][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23713_ (.CLK(clknet_leaf_318_clk_i),
    .D(_01866_),
    .RESET_B(net161),
    .Q(\line_cache[30][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23714_ (.CLK(clknet_leaf_319_clk_i),
    .D(net1110),
    .RESET_B(net159),
    .Q(\line_cache[30][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23715_ (.CLK(clknet_leaf_320_clk_i),
    .D(net2177),
    .RESET_B(net159),
    .Q(\line_cache[30][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23716_ (.CLK(clknet_leaf_320_clk_i),
    .D(net1352),
    .RESET_B(net159),
    .Q(\line_cache[30][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23717_ (.CLK(clknet_leaf_8_clk_i),
    .D(_01870_),
    .RESET_B(net159),
    .Q(\line_cache[30][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23718_ (.CLK(clknet_leaf_320_clk_i),
    .D(_01871_),
    .RESET_B(net160),
    .Q(\line_cache[30][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23719_ (.CLK(clknet_leaf_317_clk_i),
    .D(_01952_),
    .RESET_B(net179),
    .Q(\line_cache[31][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23720_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01953_),
    .RESET_B(net179),
    .Q(\line_cache[31][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23721_ (.CLK(clknet_leaf_317_clk_i),
    .D(net614),
    .RESET_B(net179),
    .Q(\line_cache[31][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23722_ (.CLK(clknet_leaf_317_clk_i),
    .D(_01955_),
    .RESET_B(net181),
    .Q(\line_cache[31][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23723_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01956_),
    .RESET_B(net181),
    .Q(\line_cache[31][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23724_ (.CLK(clknet_leaf_316_clk_i),
    .D(_01957_),
    .RESET_B(net181),
    .Q(\line_cache[31][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23725_ (.CLK(clknet_leaf_296_clk_i),
    .D(_01958_),
    .RESET_B(net181),
    .Q(\line_cache[31][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23726_ (.CLK(clknet_leaf_317_clk_i),
    .D(_01959_),
    .RESET_B(net181),
    .Q(\line_cache[31][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23727_ (.CLK(clknet_leaf_320_clk_i),
    .D(_01960_),
    .RESET_B(net159),
    .Q(\line_cache[32][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23728_ (.CLK(clknet_leaf_5_clk_i),
    .D(_01961_),
    .RESET_B(net152),
    .Q(\line_cache[32][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23729_ (.CLK(clknet_leaf_7_clk_i),
    .D(net2603),
    .RESET_B(net159),
    .Q(\line_cache[32][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23730_ (.CLK(clknet_leaf_7_clk_i),
    .D(_01963_),
    .RESET_B(net159),
    .Q(\line_cache[32][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23731_ (.CLK(clknet_leaf_320_clk_i),
    .D(_01964_),
    .RESET_B(net159),
    .Q(\line_cache[32][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23732_ (.CLK(clknet_leaf_7_clk_i),
    .D(net1590),
    .RESET_B(net159),
    .Q(\line_cache[32][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23733_ (.CLK(clknet_leaf_7_clk_i),
    .D(net3824),
    .RESET_B(net159),
    .Q(\line_cache[32][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23734_ (.CLK(clknet_leaf_7_clk_i),
    .D(net3830),
    .RESET_B(net159),
    .Q(\line_cache[32][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23735_ (.CLK(clknet_leaf_4_clk_i),
    .D(net876),
    .RESET_B(net152),
    .Q(\line_cache[33][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23736_ (.CLK(clknet_leaf_2_clk_i),
    .D(_01969_),
    .RESET_B(net151),
    .Q(\line_cache[33][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23737_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01970_),
    .RESET_B(net150),
    .Q(\line_cache[33][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23738_ (.CLK(clknet_leaf_5_clk_i),
    .D(net1310),
    .RESET_B(net153),
    .Q(\line_cache[33][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23739_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01972_),
    .RESET_B(net150),
    .Q(\line_cache[33][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23740_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01973_),
    .RESET_B(net150),
    .Q(\line_cache[33][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23741_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01974_),
    .RESET_B(net152),
    .Q(\line_cache[33][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23742_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01975_),
    .RESET_B(net152),
    .Q(\line_cache[33][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23743_ (.CLK(clknet_leaf_4_clk_i),
    .D(net1098),
    .RESET_B(net153),
    .Q(\line_cache[34][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23744_ (.CLK(clknet_leaf_2_clk_i),
    .D(_01977_),
    .RESET_B(net151),
    .Q(\line_cache[34][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23745_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01978_),
    .RESET_B(net150),
    .Q(\line_cache[34][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23746_ (.CLK(clknet_leaf_2_clk_i),
    .D(net1823),
    .RESET_B(net150),
    .Q(\line_cache[34][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23747_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01980_),
    .RESET_B(net150),
    .Q(\line_cache[34][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23748_ (.CLK(clknet_leaf_1_clk_i),
    .D(_01981_),
    .RESET_B(net150),
    .Q(\line_cache[34][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23749_ (.CLK(clknet_leaf_0_clk_i),
    .D(net2338),
    .RESET_B(net152),
    .Q(\line_cache[34][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23750_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01983_),
    .RESET_B(net152),
    .Q(\line_cache[34][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23751_ (.CLK(clknet_leaf_5_clk_i),
    .D(_01984_),
    .RESET_B(net153),
    .Q(\line_cache[35][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23752_ (.CLK(clknet_leaf_2_clk_i),
    .D(net1272),
    .RESET_B(net151),
    .Q(\line_cache[35][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23753_ (.CLK(clknet_leaf_6_clk_i),
    .D(net1648),
    .RESET_B(net152),
    .Q(\line_cache[35][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23754_ (.CLK(clknet_leaf_2_clk_i),
    .D(_01987_),
    .RESET_B(net151),
    .Q(\line_cache[35][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23755_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01988_),
    .RESET_B(net152),
    .Q(\line_cache[35][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23756_ (.CLK(clknet_leaf_0_clk_i),
    .D(_01989_),
    .RESET_B(net150),
    .Q(\line_cache[35][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23757_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01990_),
    .RESET_B(net152),
    .Q(\line_cache[35][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23758_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01991_),
    .RESET_B(net152),
    .Q(\line_cache[35][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23759_ (.CLK(clknet_leaf_7_clk_i),
    .D(net1408),
    .RESET_B(net159),
    .Q(\line_cache[36][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23760_ (.CLK(clknet_leaf_3_clk_i),
    .D(_01993_),
    .RESET_B(net151),
    .Q(\line_cache[36][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23761_ (.CLK(clknet_leaf_7_clk_i),
    .D(net1492),
    .RESET_B(net159),
    .Q(\line_cache[36][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23762_ (.CLK(clknet_leaf_2_clk_i),
    .D(_01995_),
    .RESET_B(net151),
    .Q(\line_cache[36][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23763_ (.CLK(clknet_leaf_0_clk_i),
    .D(net2326),
    .RESET_B(net152),
    .Q(\line_cache[36][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23764_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01997_),
    .RESET_B(net152),
    .Q(\line_cache[36][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23765_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01998_),
    .RESET_B(net152),
    .Q(\line_cache[36][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23766_ (.CLK(clknet_leaf_6_clk_i),
    .D(_01999_),
    .RESET_B(net152),
    .Q(\line_cache[36][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23767_ (.CLK(clknet_leaf_4_clk_i),
    .D(_02000_),
    .RESET_B(net153),
    .Q(\line_cache[37][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23768_ (.CLK(clknet_leaf_7_clk_i),
    .D(net2257),
    .RESET_B(net159),
    .Q(\line_cache[37][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23769_ (.CLK(clknet_leaf_12_clk_i),
    .D(net656),
    .RESET_B(net164),
    .Q(\line_cache[37][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23770_ (.CLK(clknet_leaf_8_clk_i),
    .D(net1754),
    .RESET_B(net159),
    .Q(\line_cache[37][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23771_ (.CLK(clknet_leaf_4_clk_i),
    .D(net778),
    .RESET_B(net153),
    .Q(\line_cache[37][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23772_ (.CLK(clknet_leaf_3_clk_i),
    .D(_02005_),
    .RESET_B(net151),
    .Q(\line_cache[37][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23773_ (.CLK(clknet_leaf_4_clk_i),
    .D(_02006_),
    .RESET_B(net153),
    .Q(\line_cache[37][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23774_ (.CLK(clknet_leaf_13_clk_i),
    .D(_02007_),
    .RESET_B(net151),
    .Q(\line_cache[37][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23775_ (.CLK(clknet_leaf_4_clk_i),
    .D(_02008_),
    .RESET_B(net153),
    .Q(\line_cache[38][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23776_ (.CLK(clknet_leaf_3_clk_i),
    .D(_02009_),
    .RESET_B(net151),
    .Q(\line_cache[38][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23777_ (.CLK(clknet_leaf_13_clk_i),
    .D(_02010_),
    .RESET_B(net162),
    .Q(\line_cache[38][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23778_ (.CLK(clknet_leaf_4_clk_i),
    .D(_02011_),
    .RESET_B(net153),
    .Q(\line_cache[38][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23779_ (.CLK(clknet_leaf_3_clk_i),
    .D(_02012_),
    .RESET_B(net151),
    .Q(\line_cache[38][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23780_ (.CLK(clknet_leaf_4_clk_i),
    .D(net882),
    .RESET_B(net151),
    .Q(\line_cache[38][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23781_ (.CLK(clknet_leaf_10_clk_i),
    .D(net1400),
    .RESET_B(net169),
    .Q(\line_cache[38][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23782_ (.CLK(clknet_leaf_13_clk_i),
    .D(net856),
    .RESET_B(net162),
    .Q(\line_cache[38][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23783_ (.CLK(clknet_leaf_8_clk_i),
    .D(net1534),
    .RESET_B(net159),
    .Q(\line_cache[39][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23784_ (.CLK(clknet_leaf_8_clk_i),
    .D(net1216),
    .RESET_B(net161),
    .Q(\line_cache[39][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23785_ (.CLK(clknet_leaf_12_clk_i),
    .D(net796),
    .RESET_B(net164),
    .Q(\line_cache[39][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23786_ (.CLK(clknet_leaf_8_clk_i),
    .D(net1891),
    .RESET_B(net161),
    .Q(\line_cache[39][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23787_ (.CLK(clknet_leaf_5_clk_i),
    .D(_02020_),
    .RESET_B(net153),
    .Q(\line_cache[39][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23788_ (.CLK(clknet_leaf_9_clk_i),
    .D(net2149),
    .RESET_B(net169),
    .Q(\line_cache[39][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23789_ (.CLK(clknet_leaf_9_clk_i),
    .D(net1198),
    .RESET_B(net169),
    .Q(\line_cache[39][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23790_ (.CLK(clknet_leaf_9_clk_i),
    .D(net2349),
    .RESET_B(net170),
    .Q(\line_cache[39][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23791_ (.CLK(clknet_leaf_5_clk_i),
    .D(net500),
    .RESET_B(net153),
    .Q(\line_cache[40][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23792_ (.CLK(clknet_leaf_317_clk_i),
    .D(_02033_),
    .RESET_B(net161),
    .Q(\line_cache[40][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23793_ (.CLK(clknet_leaf_12_clk_i),
    .D(net1330),
    .RESET_B(net161),
    .Q(\line_cache[40][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23794_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02035_),
    .RESET_B(net161),
    .Q(\line_cache[40][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23795_ (.CLK(clknet_leaf_5_clk_i),
    .D(net1478),
    .RESET_B(net153),
    .Q(\line_cache[40][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23796_ (.CLK(clknet_leaf_8_clk_i),
    .D(net3800),
    .RESET_B(net161),
    .Q(\line_cache[40][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23797_ (.CLK(clknet_leaf_8_clk_i),
    .D(net3996),
    .RESET_B(net161),
    .Q(\line_cache[40][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23798_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02039_),
    .RESET_B(net161),
    .Q(\line_cache[40][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23799_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02040_),
    .RESET_B(net175),
    .Q(\line_cache[41][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23800_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02041_),
    .RESET_B(net175),
    .Q(\line_cache[41][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23801_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02042_),
    .RESET_B(net175),
    .Q(\line_cache[41][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23802_ (.CLK(clknet_leaf_324_clk_i),
    .D(_02043_),
    .RESET_B(net157),
    .Q(\line_cache[41][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23803_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02044_),
    .RESET_B(net158),
    .Q(\line_cache[41][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23804_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02045_),
    .RESET_B(net175),
    .Q(\line_cache[41][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23805_ (.CLK(clknet_leaf_316_clk_i),
    .D(net1270),
    .RESET_B(net179),
    .Q(\line_cache[41][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23806_ (.CLK(clknet_leaf_319_clk_i),
    .D(_02047_),
    .RESET_B(net179),
    .Q(\line_cache[41][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23807_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02048_),
    .RESET_B(net175),
    .Q(\line_cache[42][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23808_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02049_),
    .RESET_B(net175),
    .Q(\line_cache[42][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23809_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02050_),
    .RESET_B(net175),
    .Q(\line_cache[42][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23810_ (.CLK(clknet_leaf_324_clk_i),
    .D(_02051_),
    .RESET_B(net157),
    .Q(\line_cache[42][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23811_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02052_),
    .RESET_B(net176),
    .Q(\line_cache[42][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23812_ (.CLK(clknet_leaf_313_clk_i),
    .D(net820),
    .RESET_B(net176),
    .Q(\line_cache[42][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23813_ (.CLK(clknet_leaf_316_clk_i),
    .D(net1072),
    .RESET_B(net179),
    .Q(\line_cache[42][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23814_ (.CLK(clknet_leaf_316_clk_i),
    .D(net1118),
    .RESET_B(net176),
    .Q(\line_cache[42][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23815_ (.CLK(clknet_leaf_313_clk_i),
    .D(net1368),
    .RESET_B(net176),
    .Q(\line_cache[43][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23816_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02057_),
    .RESET_B(net175),
    .Q(\line_cache[43][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23817_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02058_),
    .RESET_B(net175),
    .Q(\line_cache[43][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23818_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02059_),
    .RESET_B(net175),
    .Q(\line_cache[43][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23819_ (.CLK(clknet_leaf_315_clk_i),
    .D(net2433),
    .RESET_B(net179),
    .Q(\line_cache[43][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23820_ (.CLK(clknet_leaf_316_clk_i),
    .D(net1086),
    .RESET_B(net179),
    .Q(\line_cache[43][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23821_ (.CLK(clknet_leaf_315_clk_i),
    .D(net1500),
    .RESET_B(net176),
    .Q(\line_cache[43][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23822_ (.CLK(clknet_leaf_316_clk_i),
    .D(net1390),
    .RESET_B(net179),
    .Q(\line_cache[43][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23823_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02064_),
    .RESET_B(net176),
    .Q(\line_cache[44][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23824_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02065_),
    .RESET_B(net175),
    .Q(\line_cache[44][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23825_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02066_),
    .RESET_B(net175),
    .Q(\line_cache[44][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23826_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02067_),
    .RESET_B(net175),
    .Q(\line_cache[44][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23827_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02068_),
    .RESET_B(net176),
    .Q(\line_cache[44][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23828_ (.CLK(clknet_leaf_315_clk_i),
    .D(_02069_),
    .RESET_B(net179),
    .Q(\line_cache[44][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23829_ (.CLK(clknet_leaf_315_clk_i),
    .D(_02070_),
    .RESET_B(net179),
    .Q(\line_cache[44][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23830_ (.CLK(clknet_leaf_315_clk_i),
    .D(_02071_),
    .RESET_B(net179),
    .Q(\line_cache[44][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23831_ (.CLK(clknet_leaf_314_clk_i),
    .D(_02072_),
    .RESET_B(net177),
    .Q(\line_cache[45][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23832_ (.CLK(clknet_leaf_314_clk_i),
    .D(_02073_),
    .RESET_B(net180),
    .Q(\line_cache[45][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23833_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02074_),
    .RESET_B(net176),
    .Q(\line_cache[45][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23834_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02075_),
    .RESET_B(net176),
    .Q(\line_cache[45][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23835_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02076_),
    .RESET_B(net176),
    .Q(\line_cache[45][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23836_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02077_),
    .RESET_B(net180),
    .Q(\line_cache[45][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23837_ (.CLK(clknet_leaf_315_clk_i),
    .D(_02078_),
    .RESET_B(net180),
    .Q(\line_cache[45][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23838_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02079_),
    .RESET_B(net180),
    .Q(\line_cache[45][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23839_ (.CLK(clknet_leaf_314_clk_i),
    .D(_02080_),
    .RESET_B(net177),
    .Q(\line_cache[46][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23840_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02081_),
    .RESET_B(net180),
    .Q(\line_cache[46][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23841_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02082_),
    .RESET_B(net176),
    .Q(\line_cache[46][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23842_ (.CLK(clknet_leaf_314_clk_i),
    .D(_02083_),
    .RESET_B(net177),
    .Q(\line_cache[46][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23843_ (.CLK(clknet_leaf_315_clk_i),
    .D(_02084_),
    .RESET_B(net179),
    .Q(\line_cache[46][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23844_ (.CLK(clknet_leaf_314_clk_i),
    .D(_02085_),
    .RESET_B(net180),
    .Q(\line_cache[46][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23845_ (.CLK(clknet_leaf_315_clk_i),
    .D(_02086_),
    .RESET_B(net180),
    .Q(\line_cache[46][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23846_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02087_),
    .RESET_B(net180),
    .Q(\line_cache[46][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23847_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02088_),
    .RESET_B(net181),
    .Q(\line_cache[47][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23848_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02089_),
    .RESET_B(net180),
    .Q(\line_cache[47][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23849_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02090_),
    .RESET_B(net180),
    .Q(\line_cache[47][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23850_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02091_),
    .RESET_B(net180),
    .Q(\line_cache[47][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23851_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02092_),
    .RESET_B(net180),
    .Q(\line_cache[47][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23852_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02093_),
    .RESET_B(net180),
    .Q(\line_cache[47][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23853_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02094_),
    .RESET_B(net180),
    .Q(\line_cache[47][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23854_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02095_),
    .RESET_B(net181),
    .Q(\line_cache[47][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23855_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02096_),
    .RESET_B(net177),
    .Q(\line_cache[48][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23856_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02097_),
    .RESET_B(net175),
    .Q(\line_cache[48][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23857_ (.CLK(clknet_leaf_310_clk_i),
    .D(net2216),
    .RESET_B(net177),
    .Q(\line_cache[48][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23858_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02099_),
    .RESET_B(net177),
    .Q(\line_cache[48][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23859_ (.CLK(clknet_leaf_313_clk_i),
    .D(net2239),
    .RESET_B(net178),
    .Q(\line_cache[48][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23860_ (.CLK(clknet_leaf_314_clk_i),
    .D(net1965),
    .RESET_B(net178),
    .Q(\line_cache[48][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23861_ (.CLK(clknet_leaf_314_clk_i),
    .D(net3766),
    .RESET_B(net178),
    .Q(\line_cache[48][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23862_ (.CLK(clknet_leaf_314_clk_i),
    .D(net3749),
    .RESET_B(net178),
    .Q(\line_cache[48][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23863_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02104_),
    .RESET_B(net177),
    .Q(\line_cache[49][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23864_ (.CLK(clknet_leaf_311_clk_i),
    .D(net2271),
    .RESET_B(net177),
    .Q(\line_cache[49][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23865_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02106_),
    .RESET_B(net175),
    .Q(\line_cache[49][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23866_ (.CLK(clknet_leaf_311_clk_i),
    .D(net1918),
    .RESET_B(net177),
    .Q(\line_cache[49][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23867_ (.CLK(clknet_leaf_313_clk_i),
    .D(net1016),
    .RESET_B(net175),
    .Q(\line_cache[49][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23868_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02109_),
    .RESET_B(net178),
    .Q(\line_cache[49][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23869_ (.CLK(clknet_leaf_309_clk_i),
    .D(net2305),
    .RESET_B(net178),
    .Q(\line_cache[49][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23870_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02111_),
    .RESET_B(net180),
    .Q(\line_cache[49][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23871_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02120_),
    .RESET_B(net182),
    .Q(\line_cache[50][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23872_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02121_),
    .RESET_B(net177),
    .Q(\line_cache[50][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23873_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02122_),
    .RESET_B(net182),
    .Q(\line_cache[50][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23874_ (.CLK(clknet_leaf_310_clk_i),
    .D(net1322),
    .RESET_B(net177),
    .Q(\line_cache[50][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23875_ (.CLK(clknet_leaf_309_clk_i),
    .D(net1178),
    .RESET_B(net178),
    .Q(\line_cache[50][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23876_ (.CLK(clknet_leaf_310_clk_i),
    .D(net1384),
    .RESET_B(net177),
    .Q(\line_cache[50][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23877_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02126_),
    .RESET_B(net186),
    .Q(\line_cache[50][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23878_ (.CLK(clknet_leaf_309_clk_i),
    .D(net1264),
    .RESET_B(net182),
    .Q(\line_cache[50][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23879_ (.CLK(clknet_leaf_307_clk_i),
    .D(net1250),
    .RESET_B(net182),
    .Q(\line_cache[51][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23880_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02129_),
    .RESET_B(net177),
    .Q(\line_cache[51][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23881_ (.CLK(clknet_leaf_310_clk_i),
    .D(net1046),
    .RESET_B(net182),
    .Q(\line_cache[51][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23882_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02131_),
    .RESET_B(net177),
    .Q(\line_cache[51][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23883_ (.CLK(clknet_leaf_310_clk_i),
    .D(net2560),
    .RESET_B(net177),
    .Q(\line_cache[51][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23884_ (.CLK(clknet_leaf_309_clk_i),
    .D(net2084),
    .RESET_B(net177),
    .Q(\line_cache[51][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23885_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02134_),
    .RESET_B(net178),
    .Q(\line_cache[51][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23886_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02135_),
    .RESET_B(net182),
    .Q(\line_cache[51][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23887_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02136_),
    .RESET_B(net184),
    .Q(\line_cache[52][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23888_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02137_),
    .RESET_B(net184),
    .Q(\line_cache[52][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23889_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02138_),
    .RESET_B(net184),
    .Q(\line_cache[52][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23890_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02139_),
    .RESET_B(net182),
    .Q(\line_cache[52][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23891_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02140_),
    .RESET_B(net184),
    .Q(\line_cache[52][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23892_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02141_),
    .RESET_B(net183),
    .Q(\line_cache[52][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23893_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02142_),
    .RESET_B(net183),
    .Q(\line_cache[52][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23894_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02143_),
    .RESET_B(net183),
    .Q(\line_cache[52][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23895_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02144_),
    .RESET_B(net184),
    .Q(\line_cache[53][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23896_ (.CLK(clknet_leaf_307_clk_i),
    .D(net2020),
    .RESET_B(net182),
    .Q(\line_cache[53][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23897_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02146_),
    .RESET_B(net184),
    .Q(\line_cache[53][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23898_ (.CLK(clknet_leaf_307_clk_i),
    .D(net1846),
    .RESET_B(net182),
    .Q(\line_cache[53][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23899_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02148_),
    .RESET_B(net184),
    .Q(\line_cache[53][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23900_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02149_),
    .RESET_B(net182),
    .Q(\line_cache[53][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23901_ (.CLK(clknet_leaf_309_clk_i),
    .D(net2244),
    .RESET_B(net183),
    .Q(\line_cache[53][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23902_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02151_),
    .RESET_B(net182),
    .Q(\line_cache[53][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23903_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02152_),
    .RESET_B(net184),
    .Q(\line_cache[54][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23904_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02153_),
    .RESET_B(net184),
    .Q(\line_cache[54][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23905_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02154_),
    .RESET_B(net184),
    .Q(\line_cache[54][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23906_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02155_),
    .RESET_B(net182),
    .Q(\line_cache[54][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23907_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02156_),
    .RESET_B(net184),
    .Q(\line_cache[54][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23908_ (.CLK(clknet_leaf_304_clk_i),
    .D(net1202),
    .RESET_B(net183),
    .Q(\line_cache[54][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23909_ (.CLK(clknet_leaf_307_clk_i),
    .D(net1762),
    .RESET_B(net182),
    .Q(\line_cache[54][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23910_ (.CLK(clknet_leaf_308_clk_i),
    .D(net662),
    .RESET_B(net183),
    .Q(\line_cache[54][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23911_ (.CLK(clknet_leaf_306_clk_i),
    .D(net1542),
    .RESET_B(net184),
    .Q(\line_cache[55][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23912_ (.CLK(clknet_leaf_306_clk_i),
    .D(net1644),
    .RESET_B(net184),
    .Q(\line_cache[55][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23913_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02162_),
    .RESET_B(net184),
    .Q(\line_cache[55][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23914_ (.CLK(clknet_leaf_307_clk_i),
    .D(net2179),
    .RESET_B(net182),
    .Q(\line_cache[55][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23915_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02164_),
    .RESET_B(net184),
    .Q(\line_cache[55][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23916_ (.CLK(clknet_leaf_304_clk_i),
    .D(net1734),
    .RESET_B(net183),
    .Q(\line_cache[55][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23917_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02166_),
    .RESET_B(net182),
    .Q(\line_cache[55][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23918_ (.CLK(clknet_leaf_308_clk_i),
    .D(net1563),
    .RESET_B(net182),
    .Q(\line_cache[55][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23919_ (.CLK(clknet_leaf_304_clk_i),
    .D(net2403),
    .RESET_B(net185),
    .Q(\line_cache[56][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23920_ (.CLK(clknet_leaf_304_clk_i),
    .D(net1042),
    .RESET_B(net185),
    .Q(\line_cache[56][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23921_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02170_),
    .RESET_B(net185),
    .Q(\line_cache[56][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23922_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02171_),
    .RESET_B(net186),
    .Q(\line_cache[56][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23923_ (.CLK(clknet_leaf_304_clk_i),
    .D(net2387),
    .RESET_B(net183),
    .Q(\line_cache[56][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23924_ (.CLK(clknet_leaf_298_clk_i),
    .D(net3848),
    .RESET_B(net186),
    .Q(\line_cache[56][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23925_ (.CLK(clknet_leaf_303_clk_i),
    .D(net3706),
    .RESET_B(net186),
    .Q(\line_cache[56][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23926_ (.CLK(clknet_leaf_303_clk_i),
    .D(net3733),
    .RESET_B(net183),
    .Q(\line_cache[56][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23927_ (.CLK(clknet_leaf_305_clk_i),
    .D(net1809),
    .RESET_B(net185),
    .Q(\line_cache[57][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23928_ (.CLK(clknet_leaf_302_clk_i),
    .D(net2523),
    .RESET_B(net187),
    .Q(\line_cache[57][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23929_ (.CLK(clknet_leaf_305_clk_i),
    .D(net2330),
    .RESET_B(net185),
    .Q(\line_cache[57][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23930_ (.CLK(clknet_leaf_302_clk_i),
    .D(net2492),
    .RESET_B(net186),
    .Q(\line_cache[57][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23931_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02180_),
    .RESET_B(net183),
    .Q(\line_cache[57][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23932_ (.CLK(clknet_leaf_303_clk_i),
    .D(_02181_),
    .RESET_B(net186),
    .Q(\line_cache[57][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23933_ (.CLK(clknet_leaf_302_clk_i),
    .D(net2202),
    .RESET_B(net185),
    .Q(\line_cache[57][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23934_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02183_),
    .RESET_B(net183),
    .Q(\line_cache[57][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23935_ (.CLK(clknet_leaf_302_clk_i),
    .D(_02184_),
    .RESET_B(net187),
    .Q(\line_cache[58][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23936_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02185_),
    .RESET_B(net186),
    .Q(\line_cache[58][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23937_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02186_),
    .RESET_B(net180),
    .Q(\line_cache[58][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23938_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02187_),
    .RESET_B(net186),
    .Q(\line_cache[58][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23939_ (.CLK(clknet_leaf_303_clk_i),
    .D(_02188_),
    .RESET_B(net187),
    .Q(\line_cache[58][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23940_ (.CLK(clknet_leaf_303_clk_i),
    .D(net1284),
    .RESET_B(net187),
    .Q(\line_cache[58][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23941_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02190_),
    .RESET_B(net186),
    .Q(\line_cache[58][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23942_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02191_),
    .RESET_B(net186),
    .Q(\line_cache[58][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23943_ (.CLK(clknet_leaf_301_clk_i),
    .D(net1094),
    .RESET_B(net187),
    .Q(\line_cache[59][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23944_ (.CLK(clknet_leaf_298_clk_i),
    .D(net1102),
    .RESET_B(net186),
    .Q(\line_cache[59][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23945_ (.CLK(clknet_leaf_297_clk_i),
    .D(net1998),
    .RESET_B(net181),
    .Q(\line_cache[59][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23946_ (.CLK(clknet_leaf_299_clk_i),
    .D(net2204),
    .RESET_B(net186),
    .Q(\line_cache[59][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23947_ (.CLK(clknet_leaf_299_clk_i),
    .D(net2091),
    .RESET_B(net187),
    .Q(\line_cache[59][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23948_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02197_),
    .RESET_B(net186),
    .Q(\line_cache[59][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23949_ (.CLK(clknet_leaf_303_clk_i),
    .D(net1536),
    .RESET_B(net186),
    .Q(\line_cache[59][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23950_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02199_),
    .RESET_B(net186),
    .Q(\line_cache[59][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23951_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02208_),
    .RESET_B(net187),
    .Q(\line_cache[60][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23952_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02209_),
    .RESET_B(net186),
    .Q(\line_cache[60][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23953_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02210_),
    .RESET_B(net181),
    .Q(\line_cache[60][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23954_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02211_),
    .RESET_B(net188),
    .Q(\line_cache[60][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23955_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02212_),
    .RESET_B(net187),
    .Q(\line_cache[60][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23956_ (.CLK(clknet_leaf_292_clk_i),
    .D(_02213_),
    .RESET_B(net188),
    .Q(\line_cache[60][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23957_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02214_),
    .RESET_B(net187),
    .Q(\line_cache[60][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23958_ (.CLK(clknet_leaf_299_clk_i),
    .D(net1884),
    .RESET_B(net188),
    .Q(\line_cache[60][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23959_ (.CLK(clknet_leaf_299_clk_i),
    .D(net2104),
    .RESET_B(net187),
    .Q(\line_cache[61][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23960_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02217_),
    .RESET_B(net188),
    .Q(\line_cache[61][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23961_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02218_),
    .RESET_B(net181),
    .Q(\line_cache[61][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23962_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02219_),
    .RESET_B(net188),
    .Q(\line_cache[61][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23963_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02220_),
    .RESET_B(net188),
    .Q(\line_cache[61][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23964_ (.CLK(clknet_leaf_292_clk_i),
    .D(_02221_),
    .RESET_B(net195),
    .Q(\line_cache[61][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23965_ (.CLK(clknet_leaf_291_clk_i),
    .D(net1434),
    .RESET_B(net196),
    .Q(\line_cache[61][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23966_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02223_),
    .RESET_B(net188),
    .Q(\line_cache[61][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23967_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02224_),
    .RESET_B(net188),
    .Q(\line_cache[62][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23968_ (.CLK(clknet_leaf_292_clk_i),
    .D(_02225_),
    .RESET_B(net195),
    .Q(\line_cache[62][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23969_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02226_),
    .RESET_B(net181),
    .Q(\line_cache[62][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23970_ (.CLK(clknet_leaf_292_clk_i),
    .D(net954),
    .RESET_B(net195),
    .Q(\line_cache[62][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23971_ (.CLK(clknet_leaf_290_clk_i),
    .D(net1398),
    .RESET_B(net196),
    .Q(\line_cache[62][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23972_ (.CLK(clknet_leaf_291_clk_i),
    .D(net1010),
    .RESET_B(net196),
    .Q(\line_cache[62][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23973_ (.CLK(clknet_leaf_291_clk_i),
    .D(net1496),
    .RESET_B(net196),
    .Q(\line_cache[62][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23974_ (.CLK(clknet_leaf_291_clk_i),
    .D(net1002),
    .RESET_B(net196),
    .Q(\line_cache[62][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23975_ (.CLK(clknet_leaf_292_clk_i),
    .D(_02232_),
    .RESET_B(net195),
    .Q(\line_cache[63][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23976_ (.CLK(clknet_leaf_295_clk_i),
    .D(_02233_),
    .RESET_B(net191),
    .Q(\line_cache[63][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23977_ (.CLK(clknet_leaf_292_clk_i),
    .D(_02234_),
    .RESET_B(net195),
    .Q(\line_cache[63][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23978_ (.CLK(clknet_leaf_292_clk_i),
    .D(_02235_),
    .RESET_B(net195),
    .Q(\line_cache[63][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23979_ (.CLK(clknet_leaf_295_clk_i),
    .D(_02236_),
    .RESET_B(net191),
    .Q(\line_cache[63][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23980_ (.CLK(clknet_leaf_293_clk_i),
    .D(_02237_),
    .RESET_B(net195),
    .Q(\line_cache[63][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23981_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02238_),
    .RESET_B(net181),
    .Q(\line_cache[63][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23982_ (.CLK(clknet_leaf_293_clk_i),
    .D(_02239_),
    .RESET_B(net191),
    .Q(\line_cache[63][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23983_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02240_),
    .RESET_B(net188),
    .Q(\line_cache[64][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23984_ (.CLK(clknet_leaf_267_clk_i),
    .D(_02241_),
    .RESET_B(net257),
    .Q(\line_cache[64][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23985_ (.CLK(clknet_leaf_267_clk_i),
    .D(_02242_),
    .RESET_B(net257),
    .Q(\line_cache[64][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23986_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02243_),
    .RESET_B(net257),
    .Q(\line_cache[64][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23987_ (.CLK(clknet_leaf_302_clk_i),
    .D(net1685),
    .RESET_B(net187),
    .Q(\line_cache[64][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23988_ (.CLK(clknet_leaf_304_clk_i),
    .D(net2307),
    .RESET_B(net185),
    .Q(\line_cache[64][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23989_ (.CLK(clknet_leaf_264_clk_i),
    .D(net3785),
    .RESET_B(net253),
    .Q(\line_cache[64][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23990_ (.CLK(clknet_leaf_263_clk_i),
    .D(_02247_),
    .RESET_B(net254),
    .Q(\line_cache[64][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23991_ (.CLK(clknet_leaf_302_clk_i),
    .D(_02248_),
    .RESET_B(net187),
    .Q(\line_cache[65][0] ));
 sky130_fd_sc_hd__dfrtp_1 _23992_ (.CLK(clknet_leaf_305_clk_i),
    .D(net2532),
    .RESET_B(net254),
    .Q(\line_cache[65][1] ));
 sky130_fd_sc_hd__dfrtp_1 _23993_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02250_),
    .RESET_B(net257),
    .Q(\line_cache[65][2] ));
 sky130_fd_sc_hd__dfrtp_1 _23994_ (.CLK(clknet_leaf_302_clk_i),
    .D(net2545),
    .RESET_B(net254),
    .Q(\line_cache[65][3] ));
 sky130_fd_sc_hd__dfrtp_1 _23995_ (.CLK(clknet_leaf_302_clk_i),
    .D(net504),
    .RESET_B(net187),
    .Q(\line_cache[65][4] ));
 sky130_fd_sc_hd__dfrtp_1 _23996_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02253_),
    .RESET_B(net185),
    .Q(\line_cache[65][5] ));
 sky130_fd_sc_hd__dfrtp_1 _23997_ (.CLK(clknet_leaf_305_clk_i),
    .D(net2659),
    .RESET_B(net185),
    .Q(\line_cache[65][6] ));
 sky130_fd_sc_hd__dfrtp_1 _23998_ (.CLK(clknet_leaf_264_clk_i),
    .D(_02255_),
    .RESET_B(net254),
    .Q(\line_cache[65][7] ));
 sky130_fd_sc_hd__dfrtp_1 _23999_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02256_),
    .RESET_B(net187),
    .Q(\line_cache[66][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24000_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02257_),
    .RESET_B(net259),
    .Q(\line_cache[66][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24001_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02258_),
    .RESET_B(net259),
    .Q(\line_cache[66][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24002_ (.CLK(clknet_leaf_267_clk_i),
    .D(net1096),
    .RESET_B(net257),
    .Q(\line_cache[66][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24003_ (.CLK(clknet_leaf_301_clk_i),
    .D(net960),
    .RESET_B(net187),
    .Q(\line_cache[66][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24004_ (.CLK(clknet_leaf_267_clk_i),
    .D(net896),
    .RESET_B(net257),
    .Q(\line_cache[66][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24005_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02262_),
    .RESET_B(net257),
    .Q(\line_cache[66][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24006_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02263_),
    .RESET_B(net257),
    .Q(\line_cache[66][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24007_ (.CLK(clknet_leaf_301_clk_i),
    .D(net774),
    .RESET_B(net188),
    .Q(\line_cache[67][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24008_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02265_),
    .RESET_B(net259),
    .Q(\line_cache[67][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24009_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02266_),
    .RESET_B(net259),
    .Q(\line_cache[67][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24010_ (.CLK(clknet_leaf_266_clk_i),
    .D(net2095),
    .RESET_B(net257),
    .Q(\line_cache[67][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24011_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02268_),
    .RESET_B(net187),
    .Q(\line_cache[67][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24012_ (.CLK(clknet_leaf_270_clk_i),
    .D(_02269_),
    .RESET_B(net259),
    .Q(\line_cache[67][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24013_ (.CLK(clknet_leaf_266_clk_i),
    .D(net1551),
    .RESET_B(net257),
    .Q(\line_cache[67][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24014_ (.CLK(clknet_leaf_267_clk_i),
    .D(net1935),
    .RESET_B(net257),
    .Q(\line_cache[67][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24015_ (.CLK(clknet_leaf_300_clk_i),
    .D(net676),
    .RESET_B(net188),
    .Q(\line_cache[68][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24016_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02273_),
    .RESET_B(net188),
    .Q(\line_cache[68][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24017_ (.CLK(clknet_leaf_290_clk_i),
    .D(_02274_),
    .RESET_B(net196),
    .Q(\line_cache[68][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24018_ (.CLK(clknet_leaf_281_clk_i),
    .D(_02275_),
    .RESET_B(net272),
    .Q(\line_cache[68][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24019_ (.CLK(clknet_leaf_280_clk_i),
    .D(_02276_),
    .RESET_B(net272),
    .Q(\line_cache[68][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24020_ (.CLK(clknet_leaf_290_clk_i),
    .D(_02277_),
    .RESET_B(net196),
    .Q(\line_cache[68][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24021_ (.CLK(clknet_leaf_267_clk_i),
    .D(_02278_),
    .RESET_B(net257),
    .Q(\line_cache[68][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24022_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02279_),
    .RESET_B(net257),
    .Q(\line_cache[68][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24023_ (.CLK(clknet_leaf_300_clk_i),
    .D(net752),
    .RESET_B(net188),
    .Q(\line_cache[69][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24024_ (.CLK(clknet_leaf_291_clk_i),
    .D(_02281_),
    .RESET_B(net196),
    .Q(\line_cache[69][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24025_ (.CLK(clknet_leaf_290_clk_i),
    .D(net990),
    .RESET_B(net196),
    .Q(\line_cache[69][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24026_ (.CLK(clknet_leaf_280_clk_i),
    .D(net650),
    .RESET_B(net272),
    .Q(\line_cache[69][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24027_ (.CLK(clknet_leaf_291_clk_i),
    .D(net870),
    .RESET_B(net272),
    .Q(\line_cache[69][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24028_ (.CLK(clknet_leaf_290_clk_i),
    .D(_02285_),
    .RESET_B(net197),
    .Q(\line_cache[69][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24029_ (.CLK(clknet_leaf_300_clk_i),
    .D(net2221),
    .RESET_B(net257),
    .Q(\line_cache[69][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24030_ (.CLK(clknet_leaf_281_clk_i),
    .D(_02287_),
    .RESET_B(net272),
    .Q(\line_cache[69][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24031_ (.CLK(clknet_leaf_291_clk_i),
    .D(_02296_),
    .RESET_B(net196),
    .Q(\line_cache[70][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24032_ (.CLK(clknet_leaf_279_clk_i),
    .D(_02297_),
    .RESET_B(net272),
    .Q(\line_cache[70][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24033_ (.CLK(clknet_leaf_280_clk_i),
    .D(_02298_),
    .RESET_B(net272),
    .Q(\line_cache[70][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24034_ (.CLK(clknet_leaf_268_clk_i),
    .D(net906),
    .RESET_B(net257),
    .Q(\line_cache[70][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24035_ (.CLK(clknet_leaf_280_clk_i),
    .D(_02300_),
    .RESET_B(net257),
    .Q(\line_cache[70][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24036_ (.CLK(clknet_leaf_281_clk_i),
    .D(_02301_),
    .RESET_B(net272),
    .Q(\line_cache[70][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24037_ (.CLK(clknet_leaf_268_clk_i),
    .D(net914),
    .RESET_B(net258),
    .Q(\line_cache[70][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24038_ (.CLK(clknet_leaf_267_clk_i),
    .D(net1344),
    .RESET_B(net258),
    .Q(\line_cache[70][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24039_ (.CLK(clknet_leaf_281_clk_i),
    .D(_02304_),
    .RESET_B(net272),
    .Q(\line_cache[71][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24040_ (.CLK(clknet_leaf_279_clk_i),
    .D(net600),
    .RESET_B(net272),
    .Q(\line_cache[71][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24041_ (.CLK(clknet_leaf_280_clk_i),
    .D(net832),
    .RESET_B(net272),
    .Q(\line_cache[71][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24042_ (.CLK(clknet_leaf_278_clk_i),
    .D(_02307_),
    .RESET_B(net258),
    .Q(\line_cache[71][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24043_ (.CLK(clknet_leaf_279_clk_i),
    .D(net782),
    .RESET_B(net258),
    .Q(\line_cache[71][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24044_ (.CLK(clknet_leaf_281_clk_i),
    .D(_02309_),
    .RESET_B(net272),
    .Q(\line_cache[71][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24045_ (.CLK(clknet_leaf_267_clk_i),
    .D(net1432),
    .RESET_B(net258),
    .Q(\line_cache[71][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24046_ (.CLK(clknet_leaf_268_clk_i),
    .D(net1578),
    .RESET_B(net258),
    .Q(\line_cache[71][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24047_ (.CLK(clknet_leaf_281_clk_i),
    .D(_02312_),
    .RESET_B(net272),
    .Q(\line_cache[72][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24048_ (.CLK(clknet_leaf_270_clk_i),
    .D(_02313_),
    .RESET_B(net259),
    .Q(\line_cache[72][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24049_ (.CLK(clknet_leaf_278_clk_i),
    .D(net2207),
    .RESET_B(net270),
    .Q(\line_cache[72][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24050_ (.CLK(clknet_leaf_282_clk_i),
    .D(_02315_),
    .RESET_B(net270),
    .Q(\line_cache[72][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24051_ (.CLK(clknet_leaf_269_clk_i),
    .D(net2609),
    .RESET_B(net260),
    .Q(\line_cache[72][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24052_ (.CLK(clknet_leaf_279_clk_i),
    .D(net974),
    .RESET_B(net270),
    .Q(\line_cache[72][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24053_ (.CLK(clknet_leaf_269_clk_i),
    .D(_02318_),
    .RESET_B(net260),
    .Q(\line_cache[72][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24054_ (.CLK(clknet_leaf_277_clk_i),
    .D(net1502),
    .RESET_B(net270),
    .Q(\line_cache[72][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24055_ (.CLK(clknet_leaf_269_clk_i),
    .D(_02320_),
    .RESET_B(net260),
    .Q(\line_cache[73][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24056_ (.CLK(clknet_leaf_270_clk_i),
    .D(net2124),
    .RESET_B(net259),
    .Q(\line_cache[73][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24057_ (.CLK(clknet_leaf_277_clk_i),
    .D(_02322_),
    .RESET_B(net270),
    .Q(\line_cache[73][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24058_ (.CLK(clknet_leaf_268_clk_i),
    .D(net1324),
    .RESET_B(net258),
    .Q(\line_cache[73][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24059_ (.CLK(clknet_leaf_278_clk_i),
    .D(_02324_),
    .RESET_B(net260),
    .Q(\line_cache[73][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24060_ (.CLK(clknet_leaf_282_clk_i),
    .D(_02325_),
    .RESET_B(net270),
    .Q(\line_cache[73][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24061_ (.CLK(clknet_leaf_268_clk_i),
    .D(net1565),
    .RESET_B(net258),
    .Q(\line_cache[73][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24062_ (.CLK(clknet_leaf_276_clk_i),
    .D(_02327_),
    .RESET_B(net270),
    .Q(\line_cache[73][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24063_ (.CLK(clknet_leaf_269_clk_i),
    .D(_02328_),
    .RESET_B(net260),
    .Q(\line_cache[74][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24064_ (.CLK(clknet_leaf_279_clk_i),
    .D(_02329_),
    .RESET_B(net272),
    .Q(\line_cache[74][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24065_ (.CLK(clknet_leaf_277_clk_i),
    .D(_02330_),
    .RESET_B(net270),
    .Q(\line_cache[74][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24066_ (.CLK(clknet_leaf_268_clk_i),
    .D(net452),
    .RESET_B(net258),
    .Q(\line_cache[74][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24067_ (.CLK(clknet_leaf_278_clk_i),
    .D(_02332_),
    .RESET_B(net270),
    .Q(\line_cache[74][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24068_ (.CLK(clknet_leaf_278_clk_i),
    .D(_02333_),
    .RESET_B(net270),
    .Q(\line_cache[74][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24069_ (.CLK(clknet_leaf_268_clk_i),
    .D(_02334_),
    .RESET_B(net260),
    .Q(\line_cache[74][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24070_ (.CLK(clknet_leaf_269_clk_i),
    .D(net2131),
    .RESET_B(net260),
    .Q(\line_cache[74][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24071_ (.CLK(clknet_leaf_270_clk_i),
    .D(_02336_),
    .RESET_B(net259),
    .Q(\line_cache[75][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24072_ (.CLK(clknet_leaf_278_clk_i),
    .D(_02337_),
    .RESET_B(net270),
    .Q(\line_cache[75][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24073_ (.CLK(clknet_leaf_279_clk_i),
    .D(_02338_),
    .RESET_B(net270),
    .Q(\line_cache[75][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24074_ (.CLK(clknet_leaf_270_clk_i),
    .D(net2591),
    .RESET_B(net259),
    .Q(\line_cache[75][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24075_ (.CLK(clknet_leaf_269_clk_i),
    .D(net2200),
    .RESET_B(net260),
    .Q(\line_cache[75][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24076_ (.CLK(clknet_leaf_277_clk_i),
    .D(_02341_),
    .RESET_B(net270),
    .Q(\line_cache[75][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24077_ (.CLK(clknet_leaf_269_clk_i),
    .D(net1348),
    .RESET_B(net260),
    .Q(\line_cache[75][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24078_ (.CLK(clknet_leaf_269_clk_i),
    .D(net1172),
    .RESET_B(net260),
    .Q(\line_cache[75][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24079_ (.CLK(clknet_leaf_265_clk_i),
    .D(net1282),
    .RESET_B(net255),
    .Q(\line_cache[76][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24080_ (.CLK(clknet_leaf_261_clk_i),
    .D(_02345_),
    .RESET_B(net255),
    .Q(\line_cache[76][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24081_ (.CLK(clknet_leaf_262_clk_i),
    .D(net1254),
    .RESET_B(net253),
    .Q(\line_cache[76][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24082_ (.CLK(clknet_leaf_264_clk_i),
    .D(_02347_),
    .RESET_B(net254),
    .Q(\line_cache[76][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24083_ (.CLK(clknet_leaf_263_clk_i),
    .D(net1907),
    .RESET_B(net253),
    .Q(\line_cache[76][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24084_ (.CLK(clknet_leaf_263_clk_i),
    .D(net1764),
    .RESET_B(net254),
    .Q(\line_cache[76][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24085_ (.CLK(clknet_leaf_263_clk_i),
    .D(net3108),
    .RESET_B(net254),
    .Q(\line_cache[76][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24086_ (.CLK(clknet_leaf_305_clk_i),
    .D(net3642),
    .RESET_B(net185),
    .Q(\line_cache[76][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24087_ (.CLK(clknet_leaf_262_clk_i),
    .D(_02352_),
    .RESET_B(net253),
    .Q(\line_cache[77][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24088_ (.CLK(clknet_leaf_260_clk_i),
    .D(net2167),
    .RESET_B(net255),
    .Q(\line_cache[77][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24089_ (.CLK(clknet_leaf_262_clk_i),
    .D(net1100),
    .RESET_B(net253),
    .Q(\line_cache[77][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24090_ (.CLK(clknet_leaf_264_clk_i),
    .D(net2248),
    .RESET_B(net255),
    .Q(\line_cache[77][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24091_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02356_),
    .RESET_B(net253),
    .Q(\line_cache[77][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24092_ (.CLK(clknet_leaf_262_clk_i),
    .D(_02357_),
    .RESET_B(net253),
    .Q(\line_cache[77][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24093_ (.CLK(clknet_leaf_264_clk_i),
    .D(net804),
    .RESET_B(net254),
    .Q(\line_cache[77][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24094_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02359_),
    .RESET_B(net185),
    .Q(\line_cache[77][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24095_ (.CLK(clknet_leaf_262_clk_i),
    .D(net768),
    .RESET_B(net253),
    .Q(\line_cache[78][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24096_ (.CLK(clknet_leaf_262_clk_i),
    .D(_02361_),
    .RESET_B(net253),
    .Q(\line_cache[78][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24097_ (.CLK(clknet_leaf_262_clk_i),
    .D(_02362_),
    .RESET_B(net253),
    .Q(\line_cache[78][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24098_ (.CLK(clknet_leaf_264_clk_i),
    .D(_02363_),
    .RESET_B(net254),
    .Q(\line_cache[78][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24099_ (.CLK(clknet_leaf_263_clk_i),
    .D(net2010),
    .RESET_B(net253),
    .Q(\line_cache[78][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24100_ (.CLK(clknet_leaf_260_clk_i),
    .D(net1522),
    .RESET_B(net255),
    .Q(\line_cache[78][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24101_ (.CLK(clknet_leaf_263_clk_i),
    .D(net2366),
    .RESET_B(net254),
    .Q(\line_cache[78][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24102_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02367_),
    .RESET_B(net253),
    .Q(\line_cache[78][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24103_ (.CLK(clknet_leaf_261_clk_i),
    .D(net1116),
    .RESET_B(net255),
    .Q(\line_cache[79][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24104_ (.CLK(clknet_leaf_262_clk_i),
    .D(net1138),
    .RESET_B(net253),
    .Q(\line_cache[79][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24105_ (.CLK(clknet_leaf_262_clk_i),
    .D(_02370_),
    .RESET_B(net253),
    .Q(\line_cache[79][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24106_ (.CLK(clknet_leaf_265_clk_i),
    .D(net1424),
    .RESET_B(net255),
    .Q(\line_cache[79][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24107_ (.CLK(clknet_leaf_263_clk_i),
    .D(net2280),
    .RESET_B(net184),
    .Q(\line_cache[79][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24108_ (.CLK(clknet_leaf_265_clk_i),
    .D(net1346),
    .RESET_B(net256),
    .Q(\line_cache[79][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24109_ (.CLK(clknet_leaf_262_clk_i),
    .D(_02374_),
    .RESET_B(net253),
    .Q(\line_cache[79][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24110_ (.CLK(clknet_leaf_263_clk_i),
    .D(_02375_),
    .RESET_B(net254),
    .Q(\line_cache[79][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24111_ (.CLK(clknet_leaf_261_clk_i),
    .D(_02384_),
    .RESET_B(net255),
    .Q(\line_cache[80][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24112_ (.CLK(clknet_leaf_257_clk_i),
    .D(net1334),
    .RESET_B(net262),
    .Q(\line_cache[80][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24113_ (.CLK(clknet_leaf_261_clk_i),
    .D(_02386_),
    .RESET_B(net262),
    .Q(\line_cache[80][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24114_ (.CLK(clknet_leaf_259_clk_i),
    .D(_02387_),
    .RESET_B(net255),
    .Q(\line_cache[80][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24115_ (.CLK(clknet_leaf_260_clk_i),
    .D(_02388_),
    .RESET_B(net255),
    .Q(\line_cache[80][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24116_ (.CLK(clknet_leaf_265_clk_i),
    .D(net2261),
    .RESET_B(net256),
    .Q(\line_cache[80][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24117_ (.CLK(clknet_leaf_258_clk_i),
    .D(_02390_),
    .RESET_B(net262),
    .Q(\line_cache[80][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24118_ (.CLK(clknet_leaf_258_clk_i),
    .D(_02391_),
    .RESET_B(net262),
    .Q(\line_cache[80][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24119_ (.CLK(clknet_leaf_261_clk_i),
    .D(net948),
    .RESET_B(net255),
    .Q(\line_cache[81][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24120_ (.CLK(clknet_leaf_257_clk_i),
    .D(net1340),
    .RESET_B(net262),
    .Q(\line_cache[81][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24121_ (.CLK(clknet_leaf_260_clk_i),
    .D(net840),
    .RESET_B(net262),
    .Q(\line_cache[81][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24122_ (.CLK(clknet_leaf_259_clk_i),
    .D(_02395_),
    .RESET_B(net256),
    .Q(\line_cache[81][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24123_ (.CLK(clknet_leaf_260_clk_i),
    .D(net880),
    .RESET_B(net262),
    .Q(\line_cache[81][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24124_ (.CLK(clknet_leaf_259_clk_i),
    .D(_02397_),
    .RESET_B(net256),
    .Q(\line_cache[81][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24125_ (.CLK(clknet_leaf_253_clk_i),
    .D(net1555),
    .RESET_B(net263),
    .Q(\line_cache[81][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24126_ (.CLK(clknet_leaf_259_clk_i),
    .D(_02399_),
    .RESET_B(net256),
    .Q(\line_cache[81][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24127_ (.CLK(clknet_leaf_261_clk_i),
    .D(_02400_),
    .RESET_B(net255),
    .Q(\line_cache[82][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24128_ (.CLK(clknet_leaf_257_clk_i),
    .D(_02401_),
    .RESET_B(net262),
    .Q(\line_cache[82][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24129_ (.CLK(clknet_leaf_261_clk_i),
    .D(_02402_),
    .RESET_B(net255),
    .Q(\line_cache[82][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24130_ (.CLK(clknet_leaf_265_clk_i),
    .D(net632),
    .RESET_B(net256),
    .Q(\line_cache[82][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24131_ (.CLK(clknet_leaf_260_clk_i),
    .D(_02404_),
    .RESET_B(net255),
    .Q(\line_cache[82][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24132_ (.CLK(clknet_leaf_265_clk_i),
    .D(net610),
    .RESET_B(net256),
    .Q(\line_cache[82][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24133_ (.CLK(clknet_leaf_259_clk_i),
    .D(net1170),
    .RESET_B(net263),
    .Q(\line_cache[82][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24134_ (.CLK(clknet_leaf_259_clk_i),
    .D(net654),
    .RESET_B(net263),
    .Q(\line_cache[82][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24135_ (.CLK(clknet_leaf_266_clk_i),
    .D(_02408_),
    .RESET_B(net259),
    .Q(\line_cache[83][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24136_ (.CLK(clknet_leaf_256_clk_i),
    .D(net1744),
    .RESET_B(net262),
    .Q(\line_cache[83][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24137_ (.CLK(clknet_leaf_261_clk_i),
    .D(net1222),
    .RESET_B(net255),
    .Q(\line_cache[83][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24138_ (.CLK(clknet_leaf_258_clk_i),
    .D(net2251),
    .RESET_B(net256),
    .Q(\line_cache[83][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24139_ (.CLK(clknet_leaf_260_clk_i),
    .D(_02412_),
    .RESET_B(net255),
    .Q(\line_cache[83][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24140_ (.CLK(clknet_leaf_253_clk_i),
    .D(net1512),
    .RESET_B(net256),
    .Q(\line_cache[83][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24141_ (.CLK(clknet_leaf_258_clk_i),
    .D(_02414_),
    .RESET_B(net263),
    .Q(\line_cache[83][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24142_ (.CLK(clknet_leaf_258_clk_i),
    .D(net1298),
    .RESET_B(net262),
    .Q(\line_cache[83][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24143_ (.CLK(clknet_leaf_271_clk_i),
    .D(net1064),
    .RESET_B(net259),
    .Q(\line_cache[84][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24144_ (.CLK(clknet_leaf_271_clk_i),
    .D(net822),
    .RESET_B(net266),
    .Q(\line_cache[84][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24145_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02418_),
    .RESET_B(net266),
    .Q(\line_cache[84][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24146_ (.CLK(clknet_leaf_270_clk_i),
    .D(_02419_),
    .RESET_B(net259),
    .Q(\line_cache[84][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24147_ (.CLK(clknet_leaf_266_clk_i),
    .D(net2428),
    .RESET_B(net259),
    .Q(\line_cache[84][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24148_ (.CLK(clknet_leaf_271_clk_i),
    .D(net884),
    .RESET_B(net266),
    .Q(\line_cache[84][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24149_ (.CLK(clknet_leaf_269_clk_i),
    .D(_02422_),
    .RESET_B(net260),
    .Q(\line_cache[84][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24150_ (.CLK(clknet_leaf_269_clk_i),
    .D(_02423_),
    .RESET_B(net266),
    .Q(\line_cache[84][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24151_ (.CLK(clknet_leaf_252_clk_i),
    .D(net1553),
    .RESET_B(net266),
    .Q(\line_cache[85][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24152_ (.CLK(clknet_leaf_252_clk_i),
    .D(net2253),
    .RESET_B(net266),
    .Q(\line_cache[85][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24153_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02426_),
    .RESET_B(net266),
    .Q(\line_cache[85][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24154_ (.CLK(clknet_leaf_270_clk_i),
    .D(net842),
    .RESET_B(net259),
    .Q(\line_cache[85][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24155_ (.CLK(clknet_leaf_270_clk_i),
    .D(net984),
    .RESET_B(net259),
    .Q(\line_cache[85][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24156_ (.CLK(clknet_leaf_271_clk_i),
    .D(_02429_),
    .RESET_B(net266),
    .Q(\line_cache[85][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24157_ (.CLK(clknet_leaf_270_clk_i),
    .D(net2411),
    .RESET_B(net259),
    .Q(\line_cache[85][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24158_ (.CLK(clknet_leaf_269_clk_i),
    .D(_02431_),
    .RESET_B(net266),
    .Q(\line_cache[85][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24159_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02432_),
    .RESET_B(net267),
    .Q(\line_cache[86][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24160_ (.CLK(clknet_leaf_274_clk_i),
    .D(_02433_),
    .RESET_B(net276),
    .Q(\line_cache[86][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24161_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02434_),
    .RESET_B(net267),
    .Q(\line_cache[86][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24162_ (.CLK(clknet_leaf_271_clk_i),
    .D(net854),
    .RESET_B(net266),
    .Q(\line_cache[86][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24163_ (.CLK(clknet_leaf_271_clk_i),
    .D(_02436_),
    .RESET_B(net266),
    .Q(\line_cache[86][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24164_ (.CLK(clknet_leaf_252_clk_i),
    .D(net900),
    .RESET_B(net266),
    .Q(\line_cache[86][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24165_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02438_),
    .RESET_B(net267),
    .Q(\line_cache[86][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24166_ (.CLK(clknet_leaf_272_clk_i),
    .D(net1561),
    .RESET_B(net267),
    .Q(\line_cache[86][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24167_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02440_),
    .RESET_B(net267),
    .Q(\line_cache[87][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24168_ (.CLK(clknet_leaf_278_clk_i),
    .D(_02441_),
    .RESET_B(net276),
    .Q(\line_cache[87][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24169_ (.CLK(clknet_leaf_278_clk_i),
    .D(_02442_),
    .RESET_B(net276),
    .Q(\line_cache[87][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24170_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02443_),
    .RESET_B(net266),
    .Q(\line_cache[87][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24171_ (.CLK(clknet_leaf_271_clk_i),
    .D(_02444_),
    .RESET_B(net266),
    .Q(\line_cache[87][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24172_ (.CLK(clknet_leaf_274_clk_i),
    .D(_02445_),
    .RESET_B(net276),
    .Q(\line_cache[87][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24173_ (.CLK(clknet_leaf_269_clk_i),
    .D(_02446_),
    .RESET_B(net267),
    .Q(\line_cache[87][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24174_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02447_),
    .RESET_B(net267),
    .Q(\line_cache[87][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24175_ (.CLK(clknet_leaf_273_clk_i),
    .D(_02448_),
    .RESET_B(net268),
    .Q(\line_cache[88][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24176_ (.CLK(clknet_leaf_251_clk_i),
    .D(_02449_),
    .RESET_B(net268),
    .Q(\line_cache[88][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24177_ (.CLK(clknet_leaf_250_clk_i),
    .D(net1802),
    .RESET_B(net268),
    .Q(\line_cache[88][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24178_ (.CLK(clknet_leaf_250_clk_i),
    .D(_02451_),
    .RESET_B(net268),
    .Q(\line_cache[88][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24179_ (.CLK(clknet_leaf_251_clk_i),
    .D(net1362),
    .RESET_B(net268),
    .Q(\line_cache[88][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24180_ (.CLK(clknet_leaf_251_clk_i),
    .D(net1120),
    .RESET_B(net268),
    .Q(\line_cache[88][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24181_ (.CLK(clknet_leaf_252_clk_i),
    .D(_02454_),
    .RESET_B(net266),
    .Q(\line_cache[88][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24182_ (.CLK(clknet_leaf_250_clk_i),
    .D(_02455_),
    .RESET_B(net268),
    .Q(\line_cache[88][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24183_ (.CLK(clknet_leaf_273_clk_i),
    .D(_02456_),
    .RESET_B(net277),
    .Q(\line_cache[89][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24184_ (.CLK(clknet_leaf_251_clk_i),
    .D(net2069),
    .RESET_B(net268),
    .Q(\line_cache[89][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24185_ (.CLK(clknet_leaf_273_clk_i),
    .D(_02458_),
    .RESET_B(net269),
    .Q(\line_cache[89][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24186_ (.CLK(clknet_leaf_252_clk_i),
    .D(net598),
    .RESET_B(net268),
    .Q(\line_cache[89][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24187_ (.CLK(clknet_leaf_251_clk_i),
    .D(net1925),
    .RESET_B(net268),
    .Q(\line_cache[89][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24188_ (.CLK(clknet_leaf_250_clk_i),
    .D(_02461_),
    .RESET_B(net268),
    .Q(\line_cache[89][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24189_ (.CLK(clknet_leaf_272_clk_i),
    .D(net1889),
    .RESET_B(net267),
    .Q(\line_cache[89][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24190_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02463_),
    .RESET_B(net269),
    .Q(\line_cache[89][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24191_ (.CLK(clknet_leaf_272_clk_i),
    .D(_02472_),
    .RESET_B(net268),
    .Q(\line_cache[90][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24192_ (.CLK(clknet_leaf_251_clk_i),
    .D(_02473_),
    .RESET_B(net268),
    .Q(\line_cache[90][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24193_ (.CLK(clknet_leaf_273_clk_i),
    .D(_02474_),
    .RESET_B(net269),
    .Q(\line_cache[90][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24194_ (.CLK(clknet_leaf_254_clk_i),
    .D(_02475_),
    .RESET_B(net265),
    .Q(\line_cache[90][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24195_ (.CLK(clknet_leaf_251_clk_i),
    .D(net1078),
    .RESET_B(net268),
    .Q(\line_cache[90][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24196_ (.CLK(clknet_leaf_251_clk_i),
    .D(_02477_),
    .RESET_B(net289),
    .Q(\line_cache[90][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24197_ (.CLK(clknet_leaf_252_clk_i),
    .D(net1194),
    .RESET_B(net266),
    .Q(\line_cache[90][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24198_ (.CLK(clknet_leaf_250_clk_i),
    .D(_02479_),
    .RESET_B(net269),
    .Q(\line_cache[90][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24199_ (.CLK(clknet_leaf_244_clk_i),
    .D(net2035),
    .RESET_B(net285),
    .Q(\line_cache[91][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24200_ (.CLK(clknet_leaf_248_clk_i),
    .D(net980),
    .RESET_B(net289),
    .Q(\line_cache[91][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24201_ (.CLK(clknet_leaf_250_clk_i),
    .D(_02482_),
    .RESET_B(net269),
    .Q(\line_cache[91][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24202_ (.CLK(clknet_leaf_253_clk_i),
    .D(net1044),
    .RESET_B(net265),
    .Q(\line_cache[91][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24203_ (.CLK(clknet_leaf_250_clk_i),
    .D(_02484_),
    .RESET_B(net269),
    .Q(\line_cache[91][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24204_ (.CLK(clknet_leaf_251_clk_i),
    .D(net1328),
    .RESET_B(net268),
    .Q(\line_cache[91][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24205_ (.CLK(clknet_leaf_251_clk_i),
    .D(net1252),
    .RESET_B(net268),
    .Q(\line_cache[91][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24206_ (.CLK(clknet_leaf_273_clk_i),
    .D(_02487_),
    .RESET_B(net269),
    .Q(\line_cache[91][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24207_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2265),
    .RESET_B(net265),
    .Q(\line_cache[92][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24208_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2000),
    .RESET_B(net285),
    .Q(\line_cache[92][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24209_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2370),
    .RESET_B(net264),
    .Q(\line_cache[92][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24210_ (.CLK(clknet_leaf_255_clk_i),
    .D(_02491_),
    .RESET_B(net264),
    .Q(\line_cache[92][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24211_ (.CLK(clknet_leaf_258_clk_i),
    .D(net1783),
    .RESET_B(net264),
    .Q(\line_cache[92][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24212_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2528),
    .RESET_B(net265),
    .Q(\line_cache[92][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24213_ (.CLK(clknet_leaf_253_clk_i),
    .D(_02494_),
    .RESET_B(net263),
    .Q(\line_cache[92][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24214_ (.CLK(clknet_leaf_258_clk_i),
    .D(_02495_),
    .RESET_B(net263),
    .Q(\line_cache[92][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24215_ (.CLK(clknet_leaf_255_clk_i),
    .D(_02496_),
    .RESET_B(net264),
    .Q(\line_cache[93][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24216_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2430),
    .RESET_B(net265),
    .Q(\line_cache[93][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24217_ (.CLK(clknet_leaf_254_clk_i),
    .D(net1937),
    .RESET_B(net264),
    .Q(\line_cache[93][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24218_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2078),
    .RESET_B(net265),
    .Q(\line_cache[93][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24219_ (.CLK(clknet_leaf_256_clk_i),
    .D(_02500_),
    .RESET_B(net264),
    .Q(\line_cache[93][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24220_ (.CLK(clknet_leaf_255_clk_i),
    .D(_02501_),
    .RESET_B(net264),
    .Q(\line_cache[93][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24221_ (.CLK(clknet_leaf_258_clk_i),
    .D(_02502_),
    .RESET_B(net263),
    .Q(\line_cache[93][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24222_ (.CLK(clknet_leaf_257_clk_i),
    .D(_02503_),
    .RESET_B(net262),
    .Q(\line_cache[93][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24223_ (.CLK(clknet_leaf_255_clk_i),
    .D(net1192),
    .RESET_B(net285),
    .Q(\line_cache[94][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24224_ (.CLK(clknet_leaf_244_clk_i),
    .D(_02505_),
    .RESET_B(net286),
    .Q(\line_cache[94][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24225_ (.CLK(clknet_leaf_255_clk_i),
    .D(_02506_),
    .RESET_B(net264),
    .Q(\line_cache[94][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24226_ (.CLK(clknet_leaf_254_clk_i),
    .D(_02507_),
    .RESET_B(net265),
    .Q(\line_cache[94][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24227_ (.CLK(clknet_leaf_256_clk_i),
    .D(net1617),
    .RESET_B(net264),
    .Q(\line_cache[94][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24228_ (.CLK(clknet_leaf_254_clk_i),
    .D(_02509_),
    .RESET_B(net265),
    .Q(\line_cache[94][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24229_ (.CLK(clknet_leaf_253_clk_i),
    .D(net1750),
    .RESET_B(net263),
    .Q(\line_cache[94][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24230_ (.CLK(clknet_leaf_257_clk_i),
    .D(_02511_),
    .RESET_B(net262),
    .Q(\line_cache[94][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24231_ (.CLK(clknet_leaf_243_clk_i),
    .D(net1768),
    .RESET_B(net285),
    .Q(\line_cache[95][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24232_ (.CLK(clknet_leaf_244_clk_i),
    .D(net1687),
    .RESET_B(net286),
    .Q(\line_cache[95][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24233_ (.CLK(clknet_leaf_243_clk_i),
    .D(_02514_),
    .RESET_B(net285),
    .Q(\line_cache[95][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24234_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2444),
    .RESET_B(net286),
    .Q(\line_cache[95][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24235_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2237),
    .RESET_B(net264),
    .Q(\line_cache[95][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24236_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2426),
    .RESET_B(net265),
    .Q(\line_cache[95][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24237_ (.CLK(clknet_leaf_254_clk_i),
    .D(_02518_),
    .RESET_B(net265),
    .Q(\line_cache[95][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24238_ (.CLK(clknet_leaf_254_clk_i),
    .D(net2486),
    .RESET_B(net263),
    .Q(\line_cache[95][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24239_ (.CLK(clknet_leaf_243_clk_i),
    .D(_02520_),
    .RESET_B(net285),
    .Q(\line_cache[96][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24240_ (.CLK(clknet_leaf_244_clk_i),
    .D(net1652),
    .RESET_B(net286),
    .Q(\line_cache[96][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24241_ (.CLK(clknet_leaf_244_clk_i),
    .D(net2631),
    .RESET_B(net286),
    .Q(\line_cache[96][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24242_ (.CLK(clknet_leaf_241_clk_i),
    .D(_02523_),
    .RESET_B(net287),
    .Q(\line_cache[96][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24243_ (.CLK(clknet_leaf_245_clk_i),
    .D(_02524_),
    .RESET_B(net287),
    .Q(\line_cache[96][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24244_ (.CLK(clknet_leaf_246_clk_i),
    .D(_02525_),
    .RESET_B(net291),
    .Q(\line_cache[96][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24245_ (.CLK(clknet_leaf_248_clk_i),
    .D(_02526_),
    .RESET_B(net289),
    .Q(\line_cache[96][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24246_ (.CLK(clknet_leaf_248_clk_i),
    .D(_02527_),
    .RESET_B(net289),
    .Q(\line_cache[96][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24247_ (.CLK(clknet_leaf_243_clk_i),
    .D(net1640),
    .RESET_B(net285),
    .Q(\line_cache[97][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24248_ (.CLK(clknet_leaf_244_clk_i),
    .D(net2510),
    .RESET_B(net286),
    .Q(\line_cache[97][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24249_ (.CLK(clknet_leaf_241_clk_i),
    .D(net1080),
    .RESET_B(net287),
    .Q(\line_cache[97][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24250_ (.CLK(clknet_leaf_242_clk_i),
    .D(_02531_),
    .RESET_B(net287),
    .Q(\line_cache[97][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24251_ (.CLK(clknet_leaf_245_clk_i),
    .D(net1292),
    .RESET_B(net287),
    .Q(\line_cache[97][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24252_ (.CLK(clknet_leaf_245_clk_i),
    .D(_02533_),
    .RESET_B(net287),
    .Q(\line_cache[97][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24253_ (.CLK(clknet_leaf_247_clk_i),
    .D(_02534_),
    .RESET_B(net289),
    .Q(\line_cache[97][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24254_ (.CLK(clknet_leaf_247_clk_i),
    .D(_02535_),
    .RESET_B(net291),
    .Q(\line_cache[97][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24255_ (.CLK(clknet_leaf_244_clk_i),
    .D(_02536_),
    .RESET_B(net286),
    .Q(\line_cache[98][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24256_ (.CLK(clknet_leaf_243_clk_i),
    .D(_02537_),
    .RESET_B(net285),
    .Q(\line_cache[98][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24257_ (.CLK(clknet_leaf_241_clk_i),
    .D(_02538_),
    .RESET_B(net287),
    .Q(\line_cache[98][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24258_ (.CLK(clknet_leaf_244_clk_i),
    .D(_02539_),
    .RESET_B(net288),
    .Q(\line_cache[98][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24259_ (.CLK(clknet_leaf_240_clk_i),
    .D(net834),
    .RESET_B(net288),
    .Q(\line_cache[98][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24260_ (.CLK(clknet_leaf_246_clk_i),
    .D(_02541_),
    .RESET_B(net291),
    .Q(\line_cache[98][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24261_ (.CLK(clknet_leaf_244_clk_i),
    .D(net2209),
    .RESET_B(net286),
    .Q(\line_cache[98][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24262_ (.CLK(clknet_leaf_247_clk_i),
    .D(_02543_),
    .RESET_B(net286),
    .Q(\line_cache[98][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24263_ (.CLK(clknet_leaf_240_clk_i),
    .D(_02544_),
    .RESET_B(net287),
    .Q(\line_cache[99][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24264_ (.CLK(clknet_leaf_243_clk_i),
    .D(net970),
    .RESET_B(net285),
    .Q(\line_cache[99][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24265_ (.CLK(clknet_leaf_241_clk_i),
    .D(net1714),
    .RESET_B(net287),
    .Q(\line_cache[99][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24266_ (.CLK(clknet_leaf_244_clk_i),
    .D(net2400),
    .RESET_B(net288),
    .Q(\line_cache[99][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24267_ (.CLK(clknet_leaf_245_clk_i),
    .D(net1082),
    .RESET_B(net288),
    .Q(\line_cache[99][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24268_ (.CLK(clknet_leaf_246_clk_i),
    .D(net1901),
    .RESET_B(net288),
    .Q(\line_cache[99][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24269_ (.CLK(clknet_leaf_244_clk_i),
    .D(_02550_),
    .RESET_B(net286),
    .Q(\line_cache[99][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24270_ (.CLK(clknet_leaf_244_clk_i),
    .D(_02551_),
    .RESET_B(net286),
    .Q(\line_cache[99][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24271_ (.CLK(clknet_leaf_240_clk_i),
    .D(net724),
    .RESET_B(net288),
    .Q(\line_cache[100][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24272_ (.CLK(clknet_leaf_246_clk_i),
    .D(net1929),
    .RESET_B(net291),
    .Q(\line_cache[100][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24273_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00010_),
    .RESET_B(net295),
    .Q(\line_cache[100][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24274_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00011_),
    .RESET_B(net291),
    .Q(\line_cache[100][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24275_ (.CLK(clknet_leaf_245_clk_i),
    .D(net1584),
    .RESET_B(net288),
    .Q(\line_cache[100][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24276_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00013_),
    .RESET_B(net291),
    .Q(\line_cache[100][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24277_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00014_),
    .RESET_B(net293),
    .Q(\line_cache[100][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24278_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00015_),
    .RESET_B(net291),
    .Q(\line_cache[100][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24279_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00016_),
    .RESET_B(net293),
    .Q(\line_cache[101][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24280_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00017_),
    .RESET_B(net295),
    .Q(\line_cache[101][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24281_ (.CLK(clknet_leaf_241_clk_i),
    .D(_00018_),
    .RESET_B(net287),
    .Q(\line_cache[101][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24282_ (.CLK(clknet_leaf_246_clk_i),
    .D(net770),
    .RESET_B(net288),
    .Q(\line_cache[101][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24283_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00020_),
    .RESET_B(net295),
    .Q(\line_cache[101][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24284_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00021_),
    .RESET_B(net295),
    .Q(\line_cache[101][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24285_ (.CLK(clknet_leaf_240_clk_i),
    .D(net1304),
    .RESET_B(net288),
    .Q(\line_cache[101][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24286_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00023_),
    .RESET_B(net291),
    .Q(\line_cache[101][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24287_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00024_),
    .RESET_B(net293),
    .Q(\line_cache[102][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24288_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00025_),
    .RESET_B(net295),
    .Q(\line_cache[102][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24289_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00026_),
    .RESET_B(net295),
    .Q(\line_cache[102][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24290_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00027_),
    .RESET_B(net293),
    .Q(\line_cache[102][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24291_ (.CLK(clknet_leaf_239_clk_i),
    .D(net924),
    .RESET_B(net293),
    .Q(\line_cache[102][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24292_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00029_),
    .RESET_B(net295),
    .Q(\line_cache[102][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24293_ (.CLK(clknet_leaf_240_clk_i),
    .D(net938),
    .RESET_B(net293),
    .Q(\line_cache[102][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24294_ (.CLK(clknet_leaf_236_clk_i),
    .D(net868),
    .RESET_B(net295),
    .Q(\line_cache[102][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24295_ (.CLK(clknet_leaf_239_clk_i),
    .D(net1903),
    .RESET_B(net293),
    .Q(\line_cache[103][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24296_ (.CLK(clknet_leaf_230_clk_i),
    .D(net1160),
    .RESET_B(net295),
    .Q(\line_cache[103][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24297_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00034_),
    .RESET_B(net293),
    .Q(\line_cache[103][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24298_ (.CLK(clknet_leaf_236_clk_i),
    .D(net702),
    .RESET_B(net293),
    .Q(\line_cache[103][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24299_ (.CLK(clknet_leaf_239_clk_i),
    .D(net764),
    .RESET_B(net293),
    .Q(\line_cache[103][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24300_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00037_),
    .RESET_B(net295),
    .Q(\line_cache[103][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24301_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00038_),
    .RESET_B(net294),
    .Q(\line_cache[103][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24302_ (.CLK(clknet_leaf_236_clk_i),
    .D(net1758),
    .RESET_B(net294),
    .Q(\line_cache[103][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24303_ (.CLK(clknet_leaf_237_clk_i),
    .D(net1858),
    .RESET_B(net294),
    .Q(\line_cache[104][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24304_ (.CLK(clknet_leaf_237_clk_i),
    .D(net942),
    .RESET_B(net294),
    .Q(\line_cache[104][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24305_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00042_),
    .RESET_B(net297),
    .Q(\line_cache[104][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24306_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00043_),
    .RESET_B(net297),
    .Q(\line_cache[104][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24307_ (.CLK(clknet_leaf_237_clk_i),
    .D(net540),
    .RESET_B(net294),
    .Q(\line_cache[104][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24308_ (.CLK(clknet_leaf_235_clk_i),
    .D(net1168),
    .RESET_B(net297),
    .Q(\line_cache[104][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24309_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00046_),
    .RESET_B(net295),
    .Q(\line_cache[104][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24310_ (.CLK(clknet_leaf_235_clk_i),
    .D(net1602),
    .RESET_B(net297),
    .Q(\line_cache[104][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24311_ (.CLK(clknet_leaf_239_clk_i),
    .D(net626),
    .RESET_B(net294),
    .Q(\line_cache[105][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24312_ (.CLK(clknet_leaf_237_clk_i),
    .D(net2438),
    .RESET_B(net294),
    .Q(\line_cache[105][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24313_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00050_),
    .RESET_B(net297),
    .Q(\line_cache[105][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24314_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00051_),
    .RESET_B(net297),
    .Q(\line_cache[105][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24315_ (.CLK(clknet_leaf_237_clk_i),
    .D(net1278),
    .RESET_B(net294),
    .Q(\line_cache[105][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24316_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00053_),
    .RESET_B(net297),
    .Q(\line_cache[105][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24317_ (.CLK(clknet_leaf_235_clk_i),
    .D(net2100),
    .RESET_B(net295),
    .Q(\line_cache[105][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24318_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00055_),
    .RESET_B(net297),
    .Q(\line_cache[105][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24319_ (.CLK(clknet_leaf_236_clk_i),
    .D(net508),
    .RESET_B(net294),
    .Q(\line_cache[106][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24320_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00057_),
    .RESET_B(net297),
    .Q(\line_cache[106][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24321_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00058_),
    .RESET_B(net297),
    .Q(\line_cache[106][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24322_ (.CLK(clknet_leaf_230_clk_i),
    .D(net1611),
    .RESET_B(net295),
    .Q(\line_cache[106][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24323_ (.CLK(clknet_leaf_237_clk_i),
    .D(net744),
    .RESET_B(net294),
    .Q(\line_cache[106][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24324_ (.CLK(clknet_leaf_235_clk_i),
    .D(net1230),
    .RESET_B(net295),
    .Q(\line_cache[106][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24325_ (.CLK(clknet_leaf_230_clk_i),
    .D(net1136),
    .RESET_B(net295),
    .Q(\line_cache[106][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24326_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00063_),
    .RESET_B(net297),
    .Q(\line_cache[106][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24327_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00064_),
    .RESET_B(net295),
    .Q(\line_cache[107][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24328_ (.CLK(clknet_leaf_235_clk_i),
    .D(net1444),
    .RESET_B(net297),
    .Q(\line_cache[107][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24329_ (.CLK(clknet_leaf_234_clk_i),
    .D(net1320),
    .RESET_B(net297),
    .Q(\line_cache[107][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24330_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00067_),
    .RESET_B(net296),
    .Q(\line_cache[107][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24331_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00068_),
    .RESET_B(net297),
    .Q(\line_cache[107][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24332_ (.CLK(clknet_leaf_235_clk_i),
    .D(net1342),
    .RESET_B(net297),
    .Q(\line_cache[107][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24333_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00070_),
    .RESET_B(net296),
    .Q(\line_cache[107][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24334_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00071_),
    .RESET_B(net297),
    .Q(\line_cache[107][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24335_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1248),
    .RESET_B(net296),
    .Q(\line_cache[108][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24336_ (.CLK(clknet_leaf_222_clk_i),
    .D(net996),
    .RESET_B(net309),
    .Q(\line_cache[108][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24337_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00074_),
    .RESET_B(net298),
    .Q(\line_cache[108][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24338_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00075_),
    .RESET_B(net309),
    .Q(\line_cache[108][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24339_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00076_),
    .RESET_B(net309),
    .Q(\line_cache[108][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24340_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1690),
    .RESET_B(net298),
    .Q(\line_cache[108][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24341_ (.CLK(clknet_leaf_226_clk_i),
    .D(net2684),
    .RESET_B(net301),
    .Q(\line_cache[108][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24342_ (.CLK(clknet_leaf_233_clk_i),
    .D(net898),
    .RESET_B(net298),
    .Q(\line_cache[108][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24343_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00080_),
    .RESET_B(net308),
    .Q(\line_cache[109][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24344_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00081_),
    .RESET_B(net309),
    .Q(\line_cache[109][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24345_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00082_),
    .RESET_B(net298),
    .Q(\line_cache[109][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24346_ (.CLK(clknet_leaf_233_clk_i),
    .D(net908),
    .RESET_B(net298),
    .Q(\line_cache[109][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24347_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00084_),
    .RESET_B(net309),
    .Q(\line_cache[109][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24348_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00085_),
    .RESET_B(net298),
    .Q(\line_cache[109][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24349_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1152),
    .RESET_B(net296),
    .Q(\line_cache[109][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24350_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00087_),
    .RESET_B(net298),
    .Q(\line_cache[109][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24351_ (.CLK(clknet_leaf_223_clk_i),
    .D(net1829),
    .RESET_B(net308),
    .Q(\line_cache[110][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24352_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00097_),
    .RESET_B(net308),
    .Q(\line_cache[110][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24353_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00098_),
    .RESET_B(net298),
    .Q(\line_cache[110][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24354_ (.CLK(clknet_leaf_223_clk_i),
    .D(net1242),
    .RESET_B(net296),
    .Q(\line_cache[110][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24355_ (.CLK(clknet_leaf_223_clk_i),
    .D(net1869),
    .RESET_B(net309),
    .Q(\line_cache[110][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24356_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00101_),
    .RESET_B(net298),
    .Q(\line_cache[110][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24357_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1670),
    .RESET_B(net296),
    .Q(\line_cache[110][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24358_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1316),
    .RESET_B(net296),
    .Q(\line_cache[110][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24359_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00104_),
    .RESET_B(net291),
    .Q(\line_cache[111][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24360_ (.CLK(clknet_leaf_225_clk_i),
    .D(net754),
    .RESET_B(net308),
    .Q(\line_cache[111][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24361_ (.CLK(clknet_leaf_233_clk_i),
    .D(net684),
    .RESET_B(net298),
    .Q(\line_cache[111][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24362_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1557),
    .RESET_B(net296),
    .Q(\line_cache[111][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24363_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00108_),
    .RESET_B(net309),
    .Q(\line_cache[111][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24364_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1166),
    .RESET_B(net298),
    .Q(\line_cache[111][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24365_ (.CLK(clknet_leaf_232_clk_i),
    .D(net1364),
    .RESET_B(net296),
    .Q(\line_cache[111][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24366_ (.CLK(clknet_leaf_232_clk_i),
    .D(net2230),
    .RESET_B(net296),
    .Q(\line_cache[111][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24367_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00112_),
    .RESET_B(net291),
    .Q(\line_cache[112][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24368_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00113_),
    .RESET_B(net289),
    .Q(\line_cache[112][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24369_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00114_),
    .RESET_B(net289),
    .Q(\line_cache[112][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24370_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00115_),
    .RESET_B(net291),
    .Q(\line_cache[112][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24371_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00116_),
    .RESET_B(net292),
    .Q(\line_cache[112][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24372_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00117_),
    .RESET_B(net289),
    .Q(\line_cache[112][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24373_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00118_),
    .RESET_B(net289),
    .Q(\line_cache[112][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24374_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00119_),
    .RESET_B(net290),
    .Q(\line_cache[112][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24375_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00120_),
    .RESET_B(net292),
    .Q(\line_cache[113][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24376_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00121_),
    .RESET_B(net290),
    .Q(\line_cache[113][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24377_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00122_),
    .RESET_B(net290),
    .Q(\line_cache[113][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24378_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00123_),
    .RESET_B(net292),
    .Q(\line_cache[113][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24379_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00124_),
    .RESET_B(net292),
    .Q(\line_cache[113][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24380_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00125_),
    .RESET_B(net290),
    .Q(\line_cache[113][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24381_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00126_),
    .RESET_B(net290),
    .Q(\line_cache[113][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24382_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00127_),
    .RESET_B(net290),
    .Q(\line_cache[113][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24383_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00128_),
    .RESET_B(net292),
    .Q(\line_cache[114][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24384_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00129_),
    .RESET_B(net289),
    .Q(\line_cache[114][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24385_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00130_),
    .RESET_B(net289),
    .Q(\line_cache[114][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24386_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00131_),
    .RESET_B(net291),
    .Q(\line_cache[114][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24387_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00132_),
    .RESET_B(net291),
    .Q(\line_cache[114][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24388_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00133_),
    .RESET_B(net289),
    .Q(\line_cache[114][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24389_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00134_),
    .RESET_B(net289),
    .Q(\line_cache[114][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24390_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00135_),
    .RESET_B(net290),
    .Q(\line_cache[114][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24391_ (.CLK(clknet_leaf_228_clk_i),
    .D(_00136_),
    .RESET_B(net292),
    .Q(\line_cache[115][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24392_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00137_),
    .RESET_B(net289),
    .Q(\line_cache[115][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24393_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00138_),
    .RESET_B(net291),
    .Q(\line_cache[115][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24394_ (.CLK(clknet_leaf_229_clk_i),
    .D(_00139_),
    .RESET_B(net291),
    .Q(\line_cache[115][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24395_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00140_),
    .RESET_B(net291),
    .Q(\line_cache[115][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24396_ (.CLK(clknet_leaf_251_clk_i),
    .D(_00141_),
    .RESET_B(net289),
    .Q(\line_cache[115][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24397_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00142_),
    .RESET_B(net289),
    .Q(\line_cache[115][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24398_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00143_),
    .RESET_B(net290),
    .Q(\line_cache[115][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24399_ (.CLK(clknet_leaf_226_clk_i),
    .D(net2006),
    .RESET_B(net301),
    .Q(\line_cache[116][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24400_ (.CLK(clknet_leaf_225_clk_i),
    .D(net1710),
    .RESET_B(net301),
    .Q(\line_cache[116][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24401_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00146_),
    .RESET_B(net300),
    .Q(\line_cache[116][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24402_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00147_),
    .RESET_B(net300),
    .Q(\line_cache[116][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24403_ (.CLK(clknet_leaf_226_clk_i),
    .D(net1766),
    .RESET_B(net301),
    .Q(\line_cache[116][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24404_ (.CLK(clknet_leaf_226_clk_i),
    .D(net1863),
    .RESET_B(net300),
    .Q(\line_cache[116][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24405_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00150_),
    .RESET_B(net300),
    .Q(\line_cache[116][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24406_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00151_),
    .RESET_B(net300),
    .Q(\line_cache[116][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24407_ (.CLK(clknet_leaf_225_clk_i),
    .D(net1792),
    .RESET_B(net301),
    .Q(\line_cache[117][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24408_ (.CLK(clknet_leaf_226_clk_i),
    .D(net2218),
    .RESET_B(net301),
    .Q(\line_cache[117][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24409_ (.CLK(clknet_leaf_227_clk_i),
    .D(_00154_),
    .RESET_B(net300),
    .Q(\line_cache[117][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24410_ (.CLK(clknet_leaf_206_clk_i),
    .D(net2286),
    .RESET_B(net300),
    .Q(\line_cache[117][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24411_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00156_),
    .RESET_B(net301),
    .Q(\line_cache[117][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24412_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00157_),
    .RESET_B(net300),
    .Q(\line_cache[117][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24413_ (.CLK(clknet_leaf_206_clk_i),
    .D(net1668),
    .RESET_B(net300),
    .Q(\line_cache[117][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24414_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00159_),
    .RESET_B(net277),
    .Q(\line_cache[117][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24415_ (.CLK(clknet_leaf_226_clk_i),
    .D(_00160_),
    .RESET_B(net301),
    .Q(\line_cache[118][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24416_ (.CLK(clknet_leaf_225_clk_i),
    .D(_00161_),
    .RESET_B(net301),
    .Q(\line_cache[118][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24417_ (.CLK(clknet_leaf_225_clk_i),
    .D(_00162_),
    .RESET_B(net301),
    .Q(\line_cache[118][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24418_ (.CLK(clknet_leaf_206_clk_i),
    .D(net1854),
    .RESET_B(net300),
    .Q(\line_cache[118][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24419_ (.CLK(clknet_leaf_225_clk_i),
    .D(_00164_),
    .RESET_B(net301),
    .Q(\line_cache[118][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24420_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00165_),
    .RESET_B(net277),
    .Q(\line_cache[118][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24421_ (.CLK(clknet_leaf_205_clk_i),
    .D(net2363),
    .RESET_B(net277),
    .Q(\line_cache[118][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24422_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00167_),
    .RESET_B(net290),
    .Q(\line_cache[118][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24423_ (.CLK(clknet_leaf_205_clk_i),
    .D(net2398),
    .RESET_B(net277),
    .Q(\line_cache[119][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24424_ (.CLK(clknet_leaf_226_clk_i),
    .D(net1204),
    .RESET_B(net301),
    .Q(\line_cache[119][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24425_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00170_),
    .RESET_B(net300),
    .Q(\line_cache[119][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24426_ (.CLK(clknet_leaf_205_clk_i),
    .D(net2589),
    .RESET_B(net277),
    .Q(\line_cache[119][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24427_ (.CLK(clknet_leaf_225_clk_i),
    .D(_00172_),
    .RESET_B(net301),
    .Q(\line_cache[119][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24428_ (.CLK(clknet_leaf_273_clk_i),
    .D(net1772),
    .RESET_B(net277),
    .Q(\line_cache[119][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24429_ (.CLK(clknet_leaf_205_clk_i),
    .D(net1705),
    .RESET_B(net277),
    .Q(\line_cache[119][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24430_ (.CLK(clknet_leaf_273_clk_i),
    .D(net2568),
    .RESET_B(net277),
    .Q(\line_cache[119][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24431_ (.CLK(clknet_leaf_274_clk_i),
    .D(net2314),
    .RESET_B(net276),
    .Q(\line_cache[120][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24432_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00185_),
    .RESET_B(net270),
    .Q(\line_cache[120][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24433_ (.CLK(clknet_leaf_203_clk_i),
    .D(net2151),
    .RESET_B(net277),
    .Q(\line_cache[120][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24434_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00187_),
    .RESET_B(net271),
    .Q(\line_cache[120][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24435_ (.CLK(clknet_leaf_273_clk_i),
    .D(net2008),
    .RESET_B(net277),
    .Q(\line_cache[120][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24436_ (.CLK(clknet_leaf_277_clk_i),
    .D(net2277),
    .RESET_B(net276),
    .Q(\line_cache[120][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24437_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00190_),
    .RESET_B(net276),
    .Q(\line_cache[120][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24438_ (.CLK(clknet_leaf_204_clk_i),
    .D(net694),
    .RESET_B(net278),
    .Q(\line_cache[120][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24439_ (.CLK(clknet_leaf_275_clk_i),
    .D(net1807),
    .RESET_B(net276),
    .Q(\line_cache[121][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24440_ (.CLK(clknet_leaf_277_clk_i),
    .D(net2031),
    .RESET_B(net276),
    .Q(\line_cache[121][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24441_ (.CLK(clknet_leaf_203_clk_i),
    .D(net416),
    .RESET_B(net278),
    .Q(\line_cache[121][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24442_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00195_),
    .RESET_B(net271),
    .Q(\line_cache[121][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24443_ (.CLK(clknet_leaf_274_clk_i),
    .D(net490),
    .RESET_B(net277),
    .Q(\line_cache[121][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24444_ (.CLK(clknet_leaf_277_clk_i),
    .D(_00197_),
    .RESET_B(net270),
    .Q(\line_cache[121][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24445_ (.CLK(clknet_leaf_275_clk_i),
    .D(net1446),
    .RESET_B(net276),
    .Q(\line_cache[121][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24446_ (.CLK(clknet_leaf_275_clk_i),
    .D(_00199_),
    .RESET_B(net276),
    .Q(\line_cache[121][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24447_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00200_),
    .RESET_B(net276),
    .Q(\line_cache[122][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24448_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00201_),
    .RESET_B(net271),
    .Q(\line_cache[122][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24449_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00202_),
    .RESET_B(net279),
    .Q(\line_cache[122][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24450_ (.CLK(clknet_leaf_275_clk_i),
    .D(net736),
    .RESET_B(net276),
    .Q(\line_cache[122][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24451_ (.CLK(clknet_leaf_205_clk_i),
    .D(net1841),
    .RESET_B(net277),
    .Q(\line_cache[122][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24452_ (.CLK(clknet_leaf_274_clk_i),
    .D(net1897),
    .RESET_B(net276),
    .Q(\line_cache[122][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24453_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00206_),
    .RESET_B(net271),
    .Q(\line_cache[122][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24454_ (.CLK(clknet_leaf_205_clk_i),
    .D(net2012),
    .RESET_B(net277),
    .Q(\line_cache[122][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24455_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00208_),
    .RESET_B(net279),
    .Q(\line_cache[123][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24456_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00209_),
    .RESET_B(net271),
    .Q(\line_cache[123][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24457_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00210_),
    .RESET_B(net278),
    .Q(\line_cache[123][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24458_ (.CLK(clknet_leaf_274_clk_i),
    .D(net2175),
    .RESET_B(net276),
    .Q(\line_cache[123][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24459_ (.CLK(clknet_leaf_205_clk_i),
    .D(net1634),
    .RESET_B(net277),
    .Q(\line_cache[123][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24460_ (.CLK(clknet_leaf_274_clk_i),
    .D(net1658),
    .RESET_B(net276),
    .Q(\line_cache[123][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24461_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00214_),
    .RESET_B(net271),
    .Q(\line_cache[123][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24462_ (.CLK(clknet_leaf_275_clk_i),
    .D(_00215_),
    .RESET_B(net277),
    .Q(\line_cache[123][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24463_ (.CLK(clknet_leaf_202_clk_i),
    .D(net1276),
    .RESET_B(net279),
    .Q(\line_cache[124][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24464_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00217_),
    .RESET_B(net280),
    .Q(\line_cache[124][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24465_ (.CLK(clknet_leaf_202_clk_i),
    .D(net1412),
    .RESET_B(net280),
    .Q(\line_cache[124][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24466_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00219_),
    .RESET_B(net280),
    .Q(\line_cache[124][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24467_ (.CLK(clknet_leaf_202_clk_i),
    .D(net1567),
    .RESET_B(net279),
    .Q(\line_cache[124][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24468_ (.CLK(clknet_leaf_202_clk_i),
    .D(net1989),
    .RESET_B(net279),
    .Q(\line_cache[124][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24469_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00222_),
    .RESET_B(net278),
    .Q(\line_cache[124][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24470_ (.CLK(clknet_leaf_198_clk_i),
    .D(net786),
    .RESET_B(net281),
    .Q(\line_cache[124][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24471_ (.CLK(clknet_leaf_203_clk_i),
    .D(net920),
    .RESET_B(net281),
    .Q(\line_cache[125][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24472_ (.CLK(clknet_leaf_201_clk_i),
    .D(net918),
    .RESET_B(net280),
    .Q(\line_cache[125][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24473_ (.CLK(clknet_leaf_202_clk_i),
    .D(net976),
    .RESET_B(net280),
    .Q(\line_cache[125][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24474_ (.CLK(clknet_leaf_197_clk_i),
    .D(net562),
    .RESET_B(net280),
    .Q(\line_cache[125][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24475_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00228_),
    .RESET_B(net279),
    .Q(\line_cache[125][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24476_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00229_),
    .RESET_B(net280),
    .Q(\line_cache[125][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24477_ (.CLK(clknet_leaf_203_clk_i),
    .D(net994),
    .RESET_B(net278),
    .Q(\line_cache[125][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24478_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00231_),
    .RESET_B(net281),
    .Q(\line_cache[125][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24479_ (.CLK(clknet_leaf_201_clk_i),
    .D(net1468),
    .RESET_B(net281),
    .Q(\line_cache[126][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24480_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00233_),
    .RESET_B(net280),
    .Q(\line_cache[126][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24481_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00234_),
    .RESET_B(net281),
    .Q(\line_cache[126][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24482_ (.CLK(clknet_leaf_197_clk_i),
    .D(net410),
    .RESET_B(net280),
    .Q(\line_cache[126][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24483_ (.CLK(clknet_leaf_197_clk_i),
    .D(net408),
    .RESET_B(net280),
    .Q(\line_cache[126][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24484_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00237_),
    .RESET_B(net274),
    .Q(\line_cache[126][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24485_ (.CLK(clknet_leaf_201_clk_i),
    .D(net478),
    .RESET_B(net281),
    .Q(\line_cache[126][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24486_ (.CLK(clknet_leaf_200_clk_i),
    .D(net582),
    .RESET_B(net281),
    .Q(\line_cache[126][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24487_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00240_),
    .RESET_B(net281),
    .Q(\line_cache[127][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24488_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00241_),
    .RESET_B(net280),
    .Q(\line_cache[127][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24489_ (.CLK(clknet_leaf_201_clk_i),
    .D(net1308),
    .RESET_B(net281),
    .Q(\line_cache[127][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24490_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00243_),
    .RESET_B(net280),
    .Q(\line_cache[127][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24491_ (.CLK(clknet_leaf_196_clk_i),
    .D(net2756),
    .RESET_B(net280),
    .Q(\line_cache[127][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24492_ (.CLK(clknet_leaf_202_clk_i),
    .D(net1296),
    .RESET_B(net280),
    .Q(\line_cache[127][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24493_ (.CLK(clknet_leaf_201_clk_i),
    .D(net1466),
    .RESET_B(net281),
    .Q(\line_cache[127][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24494_ (.CLK(clknet_leaf_201_clk_i),
    .D(net2145),
    .RESET_B(net281),
    .Q(\line_cache[127][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24495_ (.CLK(clknet_leaf_201_clk_i),
    .D(net2049),
    .RESET_B(net281),
    .Q(\line_cache[128][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24496_ (.CLK(clknet_leaf_208_clk_i),
    .D(net1104),
    .RESET_B(net305),
    .Q(\line_cache[128][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24497_ (.CLK(clknet_leaf_207_clk_i),
    .D(net2117),
    .RESET_B(net300),
    .Q(\line_cache[128][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24498_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00251_),
    .RESET_B(net278),
    .Q(\line_cache[128][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24499_ (.CLK(clknet_leaf_207_clk_i),
    .D(net2497),
    .RESET_B(net301),
    .Q(\line_cache[128][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24500_ (.CLK(clknet_leaf_207_clk_i),
    .D(net2455),
    .RESET_B(net300),
    .Q(\line_cache[128][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24501_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00254_),
    .RESET_B(net278),
    .Q(\line_cache[128][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24502_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00255_),
    .RESET_B(net278),
    .Q(\line_cache[128][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24503_ (.CLK(clknet_leaf_201_clk_i),
    .D(net1788),
    .RESET_B(net281),
    .Q(\line_cache[129][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24504_ (.CLK(clknet_leaf_209_clk_i),
    .D(net2494),
    .RESET_B(net303),
    .Q(\line_cache[129][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24505_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00258_),
    .RESET_B(net300),
    .Q(\line_cache[129][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24506_ (.CLK(clknet_leaf_210_clk_i),
    .D(net2484),
    .RESET_B(net303),
    .Q(\line_cache[129][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24507_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00260_),
    .RESET_B(net301),
    .Q(\line_cache[129][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24508_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00261_),
    .RESET_B(net302),
    .Q(\line_cache[129][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24509_ (.CLK(clknet_leaf_203_clk_i),
    .D(net574),
    .RESET_B(net278),
    .Q(\line_cache[129][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24510_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00263_),
    .RESET_B(net278),
    .Q(\line_cache[129][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24511_ (.CLK(clknet_leaf_210_clk_i),
    .D(net436),
    .RESET_B(net303),
    .Q(\line_cache[130][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24512_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00273_),
    .RESET_B(net302),
    .Q(\line_cache[130][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24513_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00274_),
    .RESET_B(net300),
    .Q(\line_cache[130][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24514_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00275_),
    .RESET_B(net300),
    .Q(\line_cache[130][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24515_ (.CLK(clknet_leaf_207_clk_i),
    .D(net2110),
    .RESET_B(net302),
    .Q(\line_cache[130][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24516_ (.CLK(clknet_leaf_207_clk_i),
    .D(net1851),
    .RESET_B(net307),
    .Q(\line_cache[130][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24517_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00278_),
    .RESET_B(net307),
    .Q(\line_cache[130][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24518_ (.CLK(clknet_leaf_224_clk_i),
    .D(net1356),
    .RESET_B(net302),
    .Q(\line_cache[130][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24519_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00280_),
    .RESET_B(net302),
    .Q(\line_cache[131][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24520_ (.CLK(clknet_leaf_207_clk_i),
    .D(net1228),
    .RESET_B(net302),
    .Q(\line_cache[131][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24521_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00282_),
    .RESET_B(net307),
    .Q(\line_cache[131][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24522_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00283_),
    .RESET_B(net307),
    .Q(\line_cache[131][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24523_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00284_),
    .RESET_B(net302),
    .Q(\line_cache[131][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24524_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00285_),
    .RESET_B(net302),
    .Q(\line_cache[131][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24525_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00286_),
    .RESET_B(net303),
    .Q(\line_cache[131][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24526_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00287_),
    .RESET_B(net302),
    .Q(\line_cache[131][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24527_ (.CLK(clknet_leaf_219_clk_i),
    .D(net946),
    .RESET_B(net308),
    .Q(\line_cache[132][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24528_ (.CLK(clknet_leaf_222_clk_i),
    .D(net612),
    .RESET_B(net309),
    .Q(\line_cache[132][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24529_ (.CLK(clknet_leaf_220_clk_i),
    .D(net464),
    .RESET_B(net309),
    .Q(\line_cache[132][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24530_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00291_),
    .RESET_B(net309),
    .Q(\line_cache[132][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24531_ (.CLK(clknet_leaf_224_clk_i),
    .D(net486),
    .RESET_B(net308),
    .Q(\line_cache[132][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24532_ (.CLK(clknet_leaf_224_clk_i),
    .D(net1586),
    .RESET_B(net308),
    .Q(\line_cache[132][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24533_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00294_),
    .RESET_B(net301),
    .Q(\line_cache[132][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24534_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00295_),
    .RESET_B(net302),
    .Q(\line_cache[132][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24535_ (.CLK(clknet_leaf_224_clk_i),
    .D(net1835),
    .RESET_B(net308),
    .Q(\line_cache[133][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24536_ (.CLK(clknet_leaf_222_clk_i),
    .D(net578),
    .RESET_B(net309),
    .Q(\line_cache[133][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24537_ (.CLK(clknet_leaf_220_clk_i),
    .D(net628),
    .RESET_B(net309),
    .Q(\line_cache[133][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24538_ (.CLK(clknet_leaf_223_clk_i),
    .D(net516),
    .RESET_B(net309),
    .Q(\line_cache[133][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24539_ (.CLK(clknet_leaf_220_clk_i),
    .D(net462),
    .RESET_B(net309),
    .Q(\line_cache[133][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24540_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00301_),
    .RESET_B(net308),
    .Q(\line_cache[133][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24541_ (.CLK(clknet_leaf_225_clk_i),
    .D(net1140),
    .RESET_B(net308),
    .Q(\line_cache[133][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24542_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00303_),
    .RESET_B(net308),
    .Q(\line_cache[133][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24543_ (.CLK(clknet_leaf_219_clk_i),
    .D(net1088),
    .RESET_B(net308),
    .Q(\line_cache[134][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24544_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00305_),
    .RESET_B(net310),
    .Q(\line_cache[134][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24545_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00306_),
    .RESET_B(net310),
    .Q(\line_cache[134][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24546_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00307_),
    .RESET_B(net309),
    .Q(\line_cache[134][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24547_ (.CLK(clknet_leaf_219_clk_i),
    .D(net1032),
    .RESET_B(net310),
    .Q(\line_cache[134][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24548_ (.CLK(clknet_leaf_220_clk_i),
    .D(net792),
    .RESET_B(net308),
    .Q(\line_cache[134][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24549_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00310_),
    .RESET_B(net308),
    .Q(\line_cache[134][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24550_ (.CLK(clknet_leaf_224_clk_i),
    .D(net1396),
    .RESET_B(net315),
    .Q(\line_cache[134][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24551_ (.CLK(clknet_leaf_221_clk_i),
    .D(net1186),
    .RESET_B(net310),
    .Q(\line_cache[135][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24552_ (.CLK(clknet_leaf_221_clk_i),
    .D(net828),
    .RESET_B(net310),
    .Q(\line_cache[135][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24553_ (.CLK(clknet_leaf_221_clk_i),
    .D(net1438),
    .RESET_B(net310),
    .Q(\line_cache[135][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24554_ (.CLK(clknet_leaf_220_clk_i),
    .D(net742),
    .RESET_B(net310),
    .Q(\line_cache[135][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24555_ (.CLK(clknet_leaf_219_clk_i),
    .D(net630),
    .RESET_B(net315),
    .Q(\line_cache[135][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24556_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00317_),
    .RESET_B(net309),
    .Q(\line_cache[135][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24557_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00318_),
    .RESET_B(net308),
    .Q(\line_cache[135][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24558_ (.CLK(clknet_leaf_223_clk_i),
    .D(net2029),
    .RESET_B(net308),
    .Q(\line_cache[135][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24559_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00320_),
    .RESET_B(net310),
    .Q(\line_cache[136][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24560_ (.CLK(clknet_leaf_216_clk_i),
    .D(net1569),
    .RESET_B(net313),
    .Q(\line_cache[136][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24561_ (.CLK(clknet_leaf_220_clk_i),
    .D(net858),
    .RESET_B(net310),
    .Q(\line_cache[136][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24562_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00323_),
    .RESET_B(net313),
    .Q(\line_cache[136][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24563_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00324_),
    .RESET_B(net313),
    .Q(\line_cache[136][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24564_ (.CLK(clknet_leaf_216_clk_i),
    .D(net1394),
    .RESET_B(net313),
    .Q(\line_cache[136][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24565_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00326_),
    .RESET_B(net311),
    .Q(\line_cache[136][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24566_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00327_),
    .RESET_B(net311),
    .Q(\line_cache[136][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24567_ (.CLK(clknet_leaf_217_clk_i),
    .D(net680),
    .RESET_B(net313),
    .Q(\line_cache[137][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24568_ (.CLK(clknet_leaf_217_clk_i),
    .D(net414),
    .RESET_B(net313),
    .Q(\line_cache[137][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24569_ (.CLK(clknet_leaf_220_clk_i),
    .D(net474),
    .RESET_B(net310),
    .Q(\line_cache[137][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24570_ (.CLK(clknet_leaf_218_clk_i),
    .D(net664),
    .RESET_B(net313),
    .Q(\line_cache[137][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24571_ (.CLK(clknet_leaf_218_clk_i),
    .D(net1516),
    .RESET_B(net313),
    .Q(\line_cache[137][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24572_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00333_),
    .RESET_B(net313),
    .Q(\line_cache[137][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24573_ (.CLK(clknet_leaf_218_clk_i),
    .D(net718),
    .RESET_B(net311),
    .Q(\line_cache[137][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24574_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00335_),
    .RESET_B(net313),
    .Q(\line_cache[137][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24575_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00336_),
    .RESET_B(net313),
    .Q(\line_cache[138][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24576_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00337_),
    .RESET_B(net313),
    .Q(\line_cache[138][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24577_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00338_),
    .RESET_B(net310),
    .Q(\line_cache[138][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24578_ (.CLK(clknet_leaf_218_clk_i),
    .D(net1518),
    .RESET_B(net311),
    .Q(\line_cache[138][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24579_ (.CLK(clknet_leaf_218_clk_i),
    .D(net1062),
    .RESET_B(net311),
    .Q(\line_cache[138][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24580_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00341_),
    .RESET_B(net313),
    .Q(\line_cache[138][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24581_ (.CLK(clknet_leaf_219_clk_i),
    .D(net2074),
    .RESET_B(net310),
    .Q(\line_cache[138][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24582_ (.CLK(clknet_leaf_218_clk_i),
    .D(net1018),
    .RESET_B(net311),
    .Q(\line_cache[138][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24583_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00344_),
    .RESET_B(net311),
    .Q(\line_cache[139][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24584_ (.CLK(clknet_leaf_216_clk_i),
    .D(net750),
    .RESET_B(net313),
    .Q(\line_cache[139][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24585_ (.CLK(clknet_leaf_221_clk_i),
    .D(net1238),
    .RESET_B(net310),
    .Q(\line_cache[139][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24586_ (.CLK(clknet_leaf_213_clk_i),
    .D(net1724),
    .RESET_B(net311),
    .Q(\line_cache[139][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24587_ (.CLK(clknet_leaf_218_clk_i),
    .D(net1636),
    .RESET_B(net313),
    .Q(\line_cache[139][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24588_ (.CLK(clknet_leaf_217_clk_i),
    .D(net652),
    .RESET_B(net313),
    .Q(\line_cache[139][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24589_ (.CLK(clknet_leaf_219_clk_i),
    .D(net622),
    .RESET_B(net315),
    .Q(\line_cache[139][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24590_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00351_),
    .RESET_B(net311),
    .Q(\line_cache[139][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24591_ (.CLK(clknet_leaf_214_clk_i),
    .D(net2097),
    .RESET_B(net311),
    .Q(\line_cache[140][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24592_ (.CLK(clknet_leaf_212_clk_i),
    .D(net1510),
    .RESET_B(net305),
    .Q(\line_cache[140][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24593_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00362_),
    .RESET_B(net305),
    .Q(\line_cache[140][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24594_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00363_),
    .RESET_B(net305),
    .Q(\line_cache[140][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24595_ (.CLK(clknet_leaf_213_clk_i),
    .D(net2332),
    .RESET_B(net311),
    .Q(\line_cache[140][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24596_ (.CLK(clknet_leaf_212_clk_i),
    .D(net2512),
    .RESET_B(net305),
    .Q(\line_cache[140][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24597_ (.CLK(clknet_leaf_210_clk_i),
    .D(net3807),
    .RESET_B(net303),
    .Q(\line_cache[140][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24598_ (.CLK(clknet_leaf_208_clk_i),
    .D(net1124),
    .RESET_B(net305),
    .Q(\line_cache[140][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24599_ (.CLK(clknet_leaf_213_clk_i),
    .D(net1148),
    .RESET_B(net311),
    .Q(\line_cache[141][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24600_ (.CLK(clknet_leaf_212_clk_i),
    .D(net2440),
    .RESET_B(net305),
    .Q(\line_cache[141][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24601_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00370_),
    .RESET_B(net303),
    .Q(\line_cache[141][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24602_ (.CLK(clknet_leaf_212_clk_i),
    .D(net2558),
    .RESET_B(net306),
    .Q(\line_cache[141][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24603_ (.CLK(clknet_leaf_213_clk_i),
    .D(net1028),
    .RESET_B(net311),
    .Q(\line_cache[141][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24604_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00373_),
    .RESET_B(net305),
    .Q(\line_cache[141][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24605_ (.CLK(clknet_leaf_210_clk_i),
    .D(net2347),
    .RESET_B(net303),
    .Q(\line_cache[141][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24606_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00375_),
    .RESET_B(net305),
    .Q(\line_cache[141][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24607_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00376_),
    .RESET_B(net305),
    .Q(\line_cache[142][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24608_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00377_),
    .RESET_B(net305),
    .Q(\line_cache[142][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24609_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00378_),
    .RESET_B(net305),
    .Q(\line_cache[142][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24610_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00379_),
    .RESET_B(net306),
    .Q(\line_cache[142][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24611_ (.CLK(clknet_leaf_213_clk_i),
    .D(net1996),
    .RESET_B(net311),
    .Q(\line_cache[142][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24612_ (.CLK(clknet_leaf_213_clk_i),
    .D(net1200),
    .RESET_B(net305),
    .Q(\line_cache[142][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24613_ (.CLK(clknet_leaf_210_clk_i),
    .D(net1905),
    .RESET_B(net303),
    .Q(\line_cache[142][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24614_ (.CLK(clknet_leaf_208_clk_i),
    .D(net1460),
    .RESET_B(net305),
    .Q(\line_cache[142][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24615_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00384_),
    .RESET_B(net306),
    .Q(\line_cache[143][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24616_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00385_),
    .RESET_B(net311),
    .Q(\line_cache[143][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24617_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00386_),
    .RESET_B(net306),
    .Q(\line_cache[143][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24618_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00387_),
    .RESET_B(net306),
    .Q(\line_cache[143][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24619_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00388_),
    .RESET_B(net311),
    .Q(\line_cache[143][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24620_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00389_),
    .RESET_B(net305),
    .Q(\line_cache[143][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24621_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00390_),
    .RESET_B(net303),
    .Q(\line_cache[143][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24622_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00391_),
    .RESET_B(net305),
    .Q(\line_cache[143][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24623_ (.CLK(clknet_leaf_211_clk_i),
    .D(net2039),
    .RESET_B(net303),
    .Q(\line_cache[144][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24624_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00393_),
    .RESET_B(net345),
    .Q(\line_cache[144][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24625_ (.CLK(clknet_leaf_177_clk_i),
    .D(net2016),
    .RESET_B(net345),
    .Q(\line_cache[144][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24626_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00395_),
    .RESET_B(net303),
    .Q(\line_cache[144][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24627_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00396_),
    .RESET_B(net303),
    .Q(\line_cache[144][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24628_ (.CLK(clknet_leaf_211_clk_i),
    .D(net2617),
    .RESET_B(net303),
    .Q(\line_cache[144][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24629_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00398_),
    .RESET_B(net303),
    .Q(\line_cache[144][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24630_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00399_),
    .RESET_B(net304),
    .Q(\line_cache[144][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24631_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00400_),
    .RESET_B(net304),
    .Q(\line_cache[145][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24632_ (.CLK(clknet_leaf_177_clk_i),
    .D(net2600),
    .RESET_B(net345),
    .Q(\line_cache[145][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24633_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00402_),
    .RESET_B(net306),
    .Q(\line_cache[145][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24634_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00403_),
    .RESET_B(net304),
    .Q(\line_cache[145][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24635_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00404_),
    .RESET_B(net306),
    .Q(\line_cache[145][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24636_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00405_),
    .RESET_B(net303),
    .Q(\line_cache[145][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24637_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00406_),
    .RESET_B(net345),
    .Q(\line_cache[145][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24638_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00407_),
    .RESET_B(net303),
    .Q(\line_cache[145][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24639_ (.CLK(clknet_leaf_211_clk_i),
    .D(net1162),
    .RESET_B(net304),
    .Q(\line_cache[146][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24640_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00409_),
    .RESET_B(net281),
    .Q(\line_cache[146][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24641_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00410_),
    .RESET_B(net325),
    .Q(\line_cache[146][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24642_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00411_),
    .RESET_B(net281),
    .Q(\line_cache[146][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24643_ (.CLK(clknet_leaf_211_clk_i),
    .D(net1532),
    .RESET_B(net304),
    .Q(\line_cache[146][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24644_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00413_),
    .RESET_B(net282),
    .Q(\line_cache[146][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24645_ (.CLK(clknet_leaf_211_clk_i),
    .D(net2033),
    .RESET_B(net304),
    .Q(\line_cache[146][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24646_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00415_),
    .RESET_B(net282),
    .Q(\line_cache[146][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24647_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00416_),
    .RESET_B(net306),
    .Q(\line_cache[147][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24648_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00417_),
    .RESET_B(net282),
    .Q(\line_cache[147][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24649_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00418_),
    .RESET_B(net304),
    .Q(\line_cache[147][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24650_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00419_),
    .RESET_B(net281),
    .Q(\line_cache[147][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24651_ (.CLK(clknet_leaf_211_clk_i),
    .D(net2356),
    .RESET_B(net304),
    .Q(\line_cache[147][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24652_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00421_),
    .RESET_B(net282),
    .Q(\line_cache[147][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24653_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00422_),
    .RESET_B(net282),
    .Q(\line_cache[147][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24654_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00423_),
    .RESET_B(net282),
    .Q(\line_cache[147][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24655_ (.CLK(clknet_leaf_212_clk_i),
    .D(net1224),
    .RESET_B(net312),
    .Q(\line_cache[148][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24656_ (.CLK(clknet_leaf_171_clk_i),
    .D(net1126),
    .RESET_B(net355),
    .Q(\line_cache[148][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24657_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00426_),
    .RESET_B(net355),
    .Q(\line_cache[148][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24658_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00427_),
    .RESET_B(net355),
    .Q(\line_cache[148][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24659_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00428_),
    .RESET_B(net353),
    .Q(\line_cache[148][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24660_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00429_),
    .RESET_B(net314),
    .Q(\line_cache[148][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24661_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00430_),
    .RESET_B(net312),
    .Q(\line_cache[148][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24662_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00431_),
    .RESET_B(net314),
    .Q(\line_cache[148][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24663_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00432_),
    .RESET_B(net314),
    .Q(\line_cache[149][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24664_ (.CLK(clknet_leaf_171_clk_i),
    .D(net1406),
    .RESET_B(net355),
    .Q(\line_cache[149][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24665_ (.CLK(clknet_leaf_171_clk_i),
    .D(net1182),
    .RESET_B(net355),
    .Q(\line_cache[149][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24666_ (.CLK(clknet_leaf_172_clk_i),
    .D(net756),
    .RESET_B(net312),
    .Q(\line_cache[149][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24667_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00436_),
    .RESET_B(net312),
    .Q(\line_cache[149][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24668_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00437_),
    .RESET_B(net314),
    .Q(\line_cache[149][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24669_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00438_),
    .RESET_B(net312),
    .Q(\line_cache[149][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24670_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00439_),
    .RESET_B(net314),
    .Q(\line_cache[149][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24671_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00448_),
    .RESET_B(net314),
    .Q(\line_cache[150][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24672_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00449_),
    .RESET_B(net355),
    .Q(\line_cache[150][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24673_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00450_),
    .RESET_B(net355),
    .Q(\line_cache[150][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24674_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00451_),
    .RESET_B(net353),
    .Q(\line_cache[150][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24675_ (.CLK(clknet_leaf_173_clk_i),
    .D(net844),
    .RESET_B(net353),
    .Q(\line_cache[150][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24676_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00453_),
    .RESET_B(net314),
    .Q(\line_cache[150][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24677_ (.CLK(clknet_leaf_215_clk_i),
    .D(net968),
    .RESET_B(net312),
    .Q(\line_cache[150][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24678_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00455_),
    .RESET_B(net314),
    .Q(\line_cache[150][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24679_ (.CLK(clknet_leaf_171_clk_i),
    .D(net1720),
    .RESET_B(net355),
    .Q(\line_cache[151][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24680_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00457_),
    .RESET_B(net355),
    .Q(\line_cache[151][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24681_ (.CLK(clknet_leaf_171_clk_i),
    .D(_00458_),
    .RESET_B(net355),
    .Q(\line_cache[151][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24682_ (.CLK(clknet_leaf_171_clk_i),
    .D(net2556),
    .RESET_B(net355),
    .Q(\line_cache[151][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24683_ (.CLK(clknet_leaf_172_clk_i),
    .D(net992),
    .RESET_B(net353),
    .Q(\line_cache[151][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24684_ (.CLK(clknet_leaf_215_clk_i),
    .D(net2543),
    .RESET_B(net314),
    .Q(\line_cache[151][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24685_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00462_),
    .RESET_B(net312),
    .Q(\line_cache[151][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24686_ (.CLK(clknet_leaf_215_clk_i),
    .D(net2526),
    .RESET_B(net314),
    .Q(\line_cache[151][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24687_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00464_),
    .RESET_B(net355),
    .Q(\line_cache[152][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24688_ (.CLK(clknet_leaf_169_clk_i),
    .D(net1722),
    .RESET_B(net355),
    .Q(\line_cache[152][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24689_ (.CLK(clknet_leaf_169_clk_i),
    .D(net1236),
    .RESET_B(net356),
    .Q(\line_cache[152][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24690_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00467_),
    .RESET_B(net356),
    .Q(\line_cache[152][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24691_ (.CLK(clknet_leaf_174_clk_i),
    .D(net1708),
    .RESET_B(net356),
    .Q(\line_cache[152][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24692_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00469_),
    .RESET_B(net356),
    .Q(\line_cache[152][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24693_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00470_),
    .RESET_B(net353),
    .Q(\line_cache[152][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24694_ (.CLK(clknet_leaf_170_clk_i),
    .D(net1621),
    .RESET_B(net355),
    .Q(\line_cache[152][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24695_ (.CLK(clknet_leaf_172_clk_i),
    .D(net802),
    .RESET_B(net355),
    .Q(\line_cache[153][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24696_ (.CLK(clknet_leaf_169_clk_i),
    .D(net1882),
    .RESET_B(net356),
    .Q(\line_cache[153][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24697_ (.CLK(clknet_leaf_170_clk_i),
    .D(net1916),
    .RESET_B(net356),
    .Q(\line_cache[153][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24698_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00475_),
    .RESET_B(net358),
    .Q(\line_cache[153][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24699_ (.CLK(clknet_leaf_168_clk_i),
    .D(net1164),
    .RESET_B(net353),
    .Q(\line_cache[153][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24700_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00477_),
    .RESET_B(net356),
    .Q(\line_cache[153][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24701_ (.CLK(clknet_leaf_172_clk_i),
    .D(net1134),
    .RESET_B(net353),
    .Q(\line_cache[153][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24702_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00479_),
    .RESET_B(net355),
    .Q(\line_cache[153][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24703_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00480_),
    .RESET_B(net353),
    .Q(\line_cache[154][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24704_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00481_),
    .RESET_B(net358),
    .Q(\line_cache[154][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24705_ (.CLK(clknet_leaf_169_clk_i),
    .D(_00482_),
    .RESET_B(net356),
    .Q(\line_cache[154][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24706_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00483_),
    .RESET_B(net357),
    .Q(\line_cache[154][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24707_ (.CLK(clknet_leaf_168_clk_i),
    .D(net1660),
    .RESET_B(net353),
    .Q(\line_cache[154][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24708_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00485_),
    .RESET_B(net358),
    .Q(\line_cache[154][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24709_ (.CLK(clknet_leaf_174_clk_i),
    .D(net2372),
    .RESET_B(net353),
    .Q(\line_cache[154][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24710_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00487_),
    .RESET_B(net356),
    .Q(\line_cache[154][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24711_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00488_),
    .RESET_B(net357),
    .Q(\line_cache[155][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24712_ (.CLK(clknet_leaf_169_clk_i),
    .D(net1582),
    .RESET_B(net356),
    .Q(\line_cache[155][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24713_ (.CLK(clknet_leaf_169_clk_i),
    .D(net1462),
    .RESET_B(net356),
    .Q(\line_cache[155][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24714_ (.CLK(clknet_leaf_168_clk_i),
    .D(net1480),
    .RESET_B(net353),
    .Q(\line_cache[155][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24715_ (.CLK(clknet_leaf_168_clk_i),
    .D(net1623),
    .RESET_B(net353),
    .Q(\line_cache[155][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24716_ (.CLK(clknet_leaf_169_clk_i),
    .D(net940),
    .RESET_B(net356),
    .Q(\line_cache[155][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24717_ (.CLK(clknet_leaf_174_clk_i),
    .D(net1486),
    .RESET_B(net354),
    .Q(\line_cache[155][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24718_ (.CLK(clknet_leaf_170_clk_i),
    .D(_00495_),
    .RESET_B(net356),
    .Q(\line_cache[155][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24719_ (.CLK(clknet_leaf_174_clk_i),
    .D(net2170),
    .RESET_B(net354),
    .Q(\line_cache[156][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24720_ (.CLK(clknet_leaf_175_clk_i),
    .D(net586),
    .RESET_B(net347),
    .Q(\line_cache[156][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24721_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00498_),
    .RESET_B(net347),
    .Q(\line_cache[156][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24722_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00499_),
    .RESET_B(net347),
    .Q(\line_cache[156][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24723_ (.CLK(clknet_leaf_174_clk_i),
    .D(net2321),
    .RESET_B(net354),
    .Q(\line_cache[156][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24724_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00501_),
    .RESET_B(net306),
    .Q(\line_cache[156][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24725_ (.CLK(clknet_leaf_179_clk_i),
    .D(net3840),
    .RESET_B(net347),
    .Q(\line_cache[156][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24726_ (.CLK(clknet_leaf_173_clk_i),
    .D(net688),
    .RESET_B(net353),
    .Q(\line_cache[156][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24727_ (.CLK(clknet_leaf_168_clk_i),
    .D(net1530),
    .RESET_B(net354),
    .Q(\line_cache[157][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24728_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00505_),
    .RESET_B(net347),
    .Q(\line_cache[157][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24729_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00506_),
    .RESET_B(net347),
    .Q(\line_cache[157][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24730_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00507_),
    .RESET_B(net347),
    .Q(\line_cache[157][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24731_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00508_),
    .RESET_B(net347),
    .Q(\line_cache[157][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24732_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00509_),
    .RESET_B(net347),
    .Q(\line_cache[157][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24733_ (.CLK(clknet_leaf_179_clk_i),
    .D(net2275),
    .RESET_B(net347),
    .Q(\line_cache[157][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24734_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00511_),
    .RESET_B(net347),
    .Q(\line_cache[157][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24735_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00512_),
    .RESET_B(net354),
    .Q(\line_cache[158][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24736_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00513_),
    .RESET_B(net347),
    .Q(\line_cache[158][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24737_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00514_),
    .RESET_B(net306),
    .Q(\line_cache[158][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24738_ (.CLK(clknet_leaf_174_clk_i),
    .D(net1952),
    .RESET_B(net348),
    .Q(\line_cache[158][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24739_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00516_),
    .RESET_B(net354),
    .Q(\line_cache[158][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24740_ (.CLK(clknet_leaf_176_clk_i),
    .D(net934),
    .RESET_B(net353),
    .Q(\line_cache[158][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24741_ (.CLK(clknet_leaf_179_clk_i),
    .D(net2129),
    .RESET_B(net348),
    .Q(\line_cache[158][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24742_ (.CLK(clknet_leaf_172_clk_i),
    .D(net966),
    .RESET_B(net353),
    .Q(\line_cache[158][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24743_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00520_),
    .RESET_B(net351),
    .Q(\line_cache[159][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24744_ (.CLK(clknet_leaf_173_clk_i),
    .D(net590),
    .RESET_B(net353),
    .Q(\line_cache[159][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24745_ (.CLK(clknet_leaf_173_clk_i),
    .D(net890),
    .RESET_B(net347),
    .Q(\line_cache[159][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24746_ (.CLK(clknet_leaf_179_clk_i),
    .D(net2354),
    .RESET_B(net348),
    .Q(\line_cache[159][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24747_ (.CLK(clknet_leaf_174_clk_i),
    .D(net2310),
    .RESET_B(net354),
    .Q(\line_cache[159][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24748_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00525_),
    .RESET_B(net347),
    .Q(\line_cache[159][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24749_ (.CLK(clknet_leaf_174_clk_i),
    .D(net1300),
    .RESET_B(net354),
    .Q(\line_cache[159][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24750_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00527_),
    .RESET_B(net306),
    .Q(\line_cache[159][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24751_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00536_),
    .RESET_B(net351),
    .Q(\line_cache[160][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24752_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00537_),
    .RESET_B(net351),
    .Q(\line_cache[160][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24753_ (.CLK(clknet_leaf_161_clk_i),
    .D(net1984),
    .RESET_B(net351),
    .Q(\line_cache[160][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24754_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00539_),
    .RESET_B(net351),
    .Q(\line_cache[160][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24755_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00540_),
    .RESET_B(net351),
    .Q(\line_cache[160][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24756_ (.CLK(clknet_leaf_160_clk_i),
    .D(net2065),
    .RESET_B(net351),
    .Q(\line_cache[160][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24757_ (.CLK(clknet_leaf_160_clk_i),
    .D(net4039),
    .RESET_B(net349),
    .Q(\line_cache[160][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24758_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00543_),
    .RESET_B(net349),
    .Q(\line_cache[160][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24759_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00544_),
    .RESET_B(net357),
    .Q(\line_cache[161][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24760_ (.CLK(clknet_leaf_161_clk_i),
    .D(net2267),
    .RESET_B(net357),
    .Q(\line_cache[161][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24761_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00546_),
    .RESET_B(net351),
    .Q(\line_cache[161][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24762_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00547_),
    .RESET_B(net351),
    .Q(\line_cache[161][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24763_ (.CLK(clknet_leaf_162_clk_i),
    .D(net732),
    .RESET_B(net357),
    .Q(\line_cache[161][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24764_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00549_),
    .RESET_B(net352),
    .Q(\line_cache[161][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24765_ (.CLK(clknet_leaf_161_clk_i),
    .D(net1895),
    .RESET_B(net352),
    .Q(\line_cache[161][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24766_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00551_),
    .RESET_B(net349),
    .Q(\line_cache[161][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24767_ (.CLK(clknet_leaf_162_clk_i),
    .D(net412),
    .RESET_B(net357),
    .Q(\line_cache[162][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24768_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00553_),
    .RESET_B(net351),
    .Q(\line_cache[162][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24769_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00554_),
    .RESET_B(net351),
    .Q(\line_cache[162][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24770_ (.CLK(clknet_leaf_161_clk_i),
    .D(net1594),
    .RESET_B(net352),
    .Q(\line_cache[162][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24771_ (.CLK(clknet_leaf_161_clk_i),
    .D(net1214),
    .RESET_B(net351),
    .Q(\line_cache[162][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24772_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00557_),
    .RESET_B(net352),
    .Q(\line_cache[162][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24773_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00558_),
    .RESET_B(net349),
    .Q(\line_cache[162][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24774_ (.CLK(clknet_leaf_163_clk_i),
    .D(net892),
    .RESET_B(net357),
    .Q(\line_cache[162][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24775_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00560_),
    .RESET_B(net357),
    .Q(\line_cache[163][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24776_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00561_),
    .RESET_B(net357),
    .Q(\line_cache[163][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24777_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00562_),
    .RESET_B(net351),
    .Q(\line_cache[163][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24778_ (.CLK(clknet_leaf_161_clk_i),
    .D(_00563_),
    .RESET_B(net351),
    .Q(\line_cache[163][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24779_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00564_),
    .RESET_B(net351),
    .Q(\line_cache[163][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24780_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00565_),
    .RESET_B(net352),
    .Q(\line_cache[163][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24781_ (.CLK(clknet_leaf_163_clk_i),
    .D(net1106),
    .RESET_B(net352),
    .Q(\line_cache[163][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24782_ (.CLK(clknet_leaf_163_clk_i),
    .D(net2165),
    .RESET_B(net357),
    .Q(\line_cache[163][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24783_ (.CLK(clknet_leaf_168_clk_i),
    .D(net1428),
    .RESET_B(net357),
    .Q(\line_cache[164][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24784_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00569_),
    .RESET_B(net358),
    .Q(\line_cache[164][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24785_ (.CLK(clknet_leaf_167_clk_i),
    .D(net1158),
    .RESET_B(net358),
    .Q(\line_cache[164][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24786_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00571_),
    .RESET_B(net358),
    .Q(\line_cache[164][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24787_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00572_),
    .RESET_B(net358),
    .Q(\line_cache[164][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24788_ (.CLK(clknet_leaf_165_clk_i),
    .D(net712),
    .RESET_B(net358),
    .Q(\line_cache[164][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24789_ (.CLK(clknet_leaf_163_clk_i),
    .D(_00574_),
    .RESET_B(net357),
    .Q(\line_cache[164][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24790_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00575_),
    .RESET_B(net357),
    .Q(\line_cache[164][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24791_ (.CLK(clknet_leaf_168_clk_i),
    .D(_00576_),
    .RESET_B(net357),
    .Q(\line_cache[165][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24792_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00577_),
    .RESET_B(net358),
    .Q(\line_cache[165][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24793_ (.CLK(clknet_leaf_166_clk_i),
    .D(net1190),
    .RESET_B(net358),
    .Q(\line_cache[165][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24794_ (.CLK(clknet_leaf_167_clk_i),
    .D(net922),
    .RESET_B(net358),
    .Q(\line_cache[165][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24795_ (.CLK(clknet_leaf_167_clk_i),
    .D(net1232),
    .RESET_B(net358),
    .Q(\line_cache[165][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24796_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00581_),
    .RESET_B(net358),
    .Q(\line_cache[165][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24797_ (.CLK(clknet_leaf_163_clk_i),
    .D(net2076),
    .RESET_B(net357),
    .Q(\line_cache[165][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24798_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00583_),
    .RESET_B(net358),
    .Q(\line_cache[165][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24799_ (.CLK(clknet_leaf_167_clk_i),
    .D(_00584_),
    .RESET_B(net357),
    .Q(\line_cache[166][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24800_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00585_),
    .RESET_B(net359),
    .Q(\line_cache[166][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24801_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00586_),
    .RESET_B(net359),
    .Q(\line_cache[166][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24802_ (.CLK(clknet_leaf_166_clk_i),
    .D(net904),
    .RESET_B(net359),
    .Q(\line_cache[166][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24803_ (.CLK(clknet_leaf_162_clk_i),
    .D(_00588_),
    .RESET_B(net358),
    .Q(\line_cache[166][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24804_ (.CLK(clknet_leaf_165_clk_i),
    .D(net1128),
    .RESET_B(net359),
    .Q(\line_cache[166][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24805_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00590_),
    .RESET_B(net360),
    .Q(\line_cache[166][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24806_ (.CLK(clknet_leaf_164_clk_i),
    .D(net722),
    .RESET_B(net360),
    .Q(\line_cache[166][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24807_ (.CLK(clknet_leaf_166_clk_i),
    .D(net1302),
    .RESET_B(net359),
    .Q(\line_cache[167][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24808_ (.CLK(clknet_leaf_165_clk_i),
    .D(net1008),
    .RESET_B(net359),
    .Q(\line_cache[167][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24809_ (.CLK(clknet_leaf_166_clk_i),
    .D(net1422),
    .RESET_B(net359),
    .Q(\line_cache[167][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24810_ (.CLK(clknet_leaf_166_clk_i),
    .D(_00595_),
    .RESET_B(net358),
    .Q(\line_cache[167][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24811_ (.CLK(clknet_leaf_163_clk_i),
    .D(net894),
    .RESET_B(net359),
    .Q(\line_cache[167][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24812_ (.CLK(clknet_leaf_165_clk_i),
    .D(net716),
    .RESET_B(net359),
    .Q(\line_cache[167][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24813_ (.CLK(clknet_leaf_164_clk_i),
    .D(_00598_),
    .RESET_B(net360),
    .Q(\line_cache[167][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24814_ (.CLK(clknet_leaf_164_clk_i),
    .D(net690),
    .RESET_B(net359),
    .Q(\line_cache[167][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24815_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00600_),
    .RESET_B(net368),
    .Q(\line_cache[168][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24816_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00601_),
    .RESET_B(net367),
    .Q(\line_cache[168][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24817_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00602_),
    .RESET_B(net368),
    .Q(\line_cache[168][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24818_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00603_),
    .RESET_B(net368),
    .Q(\line_cache[168][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24819_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00604_),
    .RESET_B(net359),
    .Q(\line_cache[168][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24820_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00605_),
    .RESET_B(net368),
    .Q(\line_cache[168][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24821_ (.CLK(clknet_leaf_158_clk_i),
    .D(_00606_),
    .RESET_B(net363),
    .Q(\line_cache[168][6] ));
 sky130_fd_sc_hd__dfrtp_2 _24822_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00607_),
    .RESET_B(net312),
    .Q(\line_cache[168][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24823_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00608_),
    .RESET_B(net368),
    .Q(\line_cache[169][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24824_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00609_),
    .RESET_B(net367),
    .Q(\line_cache[169][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24825_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00610_),
    .RESET_B(net368),
    .Q(\line_cache[169][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24826_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00611_),
    .RESET_B(net368),
    .Q(\line_cache[169][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24827_ (.CLK(clknet_leaf_164_clk_i),
    .D(_00612_),
    .RESET_B(net360),
    .Q(\line_cache[169][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24828_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00613_),
    .RESET_B(net368),
    .Q(\line_cache[169][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24829_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00614_),
    .RESET_B(net367),
    .Q(\line_cache[169][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24830_ (.CLK(clknet_leaf_165_clk_i),
    .D(_00615_),
    .RESET_B(net359),
    .Q(\line_cache[169][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24831_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00624_),
    .RESET_B(net368),
    .Q(\line_cache[170][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24832_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00625_),
    .RESET_B(net367),
    .Q(\line_cache[170][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24833_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00626_),
    .RESET_B(net367),
    .Q(\line_cache[170][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24834_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00627_),
    .RESET_B(net368),
    .Q(\line_cache[170][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24835_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00628_),
    .RESET_B(net368),
    .Q(\line_cache[170][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24836_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00629_),
    .RESET_B(net368),
    .Q(\line_cache[170][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24837_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00630_),
    .RESET_B(net367),
    .Q(\line_cache[170][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24838_ (.CLK(clknet_leaf_154_clk_i),
    .D(_00631_),
    .RESET_B(net368),
    .Q(\line_cache[170][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24839_ (.CLK(clknet_leaf_155_clk_i),
    .D(_00632_),
    .RESET_B(net367),
    .Q(\line_cache[171][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24840_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00633_),
    .RESET_B(net367),
    .Q(\line_cache[171][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24841_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00634_),
    .RESET_B(net367),
    .Q(\line_cache[171][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24842_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00635_),
    .RESET_B(net368),
    .Q(\line_cache[171][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24843_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00636_),
    .RESET_B(net369),
    .Q(\line_cache[171][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24844_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00637_),
    .RESET_B(net368),
    .Q(\line_cache[171][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24845_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00638_),
    .RESET_B(net368),
    .Q(\line_cache[171][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24846_ (.CLK(clknet_leaf_153_clk_i),
    .D(_00639_),
    .RESET_B(net369),
    .Q(\line_cache[171][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24847_ (.CLK(clknet_leaf_156_clk_i),
    .D(net1070),
    .RESET_B(net367),
    .Q(\line_cache[172][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24848_ (.CLK(clknet_leaf_158_clk_i),
    .D(net1280),
    .RESET_B(net363),
    .Q(\line_cache[172][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24849_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00642_),
    .RESET_B(net367),
    .Q(\line_cache[172][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24850_ (.CLK(clknet_leaf_157_clk_i),
    .D(_00643_),
    .RESET_B(net363),
    .Q(\line_cache[172][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24851_ (.CLK(clknet_leaf_158_clk_i),
    .D(net1886),
    .RESET_B(net363),
    .Q(\line_cache[172][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24852_ (.CLK(clknet_leaf_164_clk_i),
    .D(net1638),
    .RESET_B(net360),
    .Q(\line_cache[172][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24853_ (.CLK(clknet_leaf_160_clk_i),
    .D(net2676),
    .RESET_B(net352),
    .Q(\line_cache[172][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24854_ (.CLK(clknet_leaf_156_clk_i),
    .D(net1506),
    .RESET_B(net369),
    .Q(\line_cache[172][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24855_ (.CLK(clknet_leaf_157_clk_i),
    .D(net1514),
    .RESET_B(net363),
    .Q(\line_cache[173][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24856_ (.CLK(clknet_leaf_157_clk_i),
    .D(net1967),
    .RESET_B(net363),
    .Q(\line_cache[173][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24857_ (.CLK(clknet_leaf_156_clk_i),
    .D(net794),
    .RESET_B(net369),
    .Q(\line_cache[173][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24858_ (.CLK(clknet_leaf_158_clk_i),
    .D(net748),
    .RESET_B(net363),
    .Q(\line_cache[173][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24859_ (.CLK(clknet_leaf_159_clk_i),
    .D(net1482),
    .RESET_B(net363),
    .Q(\line_cache[173][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24860_ (.CLK(clknet_leaf_158_clk_i),
    .D(_00653_),
    .RESET_B(net367),
    .Q(\line_cache[173][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24861_ (.CLK(clknet_leaf_158_clk_i),
    .D(net952),
    .RESET_B(net363),
    .Q(\line_cache[173][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24862_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00655_),
    .RESET_B(net369),
    .Q(\line_cache[173][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24863_ (.CLK(clknet_leaf_150_clk_i),
    .D(_00656_),
    .RESET_B(net363),
    .Q(\line_cache[174][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24864_ (.CLK(clknet_leaf_157_clk_i),
    .D(_00657_),
    .RESET_B(net364),
    .Q(\line_cache[174][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24865_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00658_),
    .RESET_B(net369),
    .Q(\line_cache[174][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24866_ (.CLK(clknet_leaf_155_clk_i),
    .D(net1066),
    .RESET_B(net367),
    .Q(\line_cache[174][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24867_ (.CLK(clknet_leaf_158_clk_i),
    .D(net1600),
    .RESET_B(net363),
    .Q(\line_cache[174][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24868_ (.CLK(clknet_leaf_155_clk_i),
    .D(net1572),
    .RESET_B(net367),
    .Q(\line_cache[174][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24869_ (.CLK(clknet_leaf_161_clk_i),
    .D(net1752),
    .RESET_B(net352),
    .Q(\line_cache[174][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24870_ (.CLK(clknet_leaf_156_clk_i),
    .D(_00663_),
    .RESET_B(net369),
    .Q(\line_cache[174][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24871_ (.CLK(clknet_leaf_160_clk_i),
    .D(_00664_),
    .RESET_B(net352),
    .Q(\line_cache[175][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24872_ (.CLK(clknet_leaf_157_clk_i),
    .D(_00665_),
    .RESET_B(net364),
    .Q(\line_cache[175][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24873_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00666_),
    .RESET_B(net369),
    .Q(\line_cache[175][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24874_ (.CLK(clknet_leaf_158_clk_i),
    .D(net1290),
    .RESET_B(net367),
    .Q(\line_cache[175][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24875_ (.CLK(clknet_leaf_157_clk_i),
    .D(_00668_),
    .RESET_B(net369),
    .Q(\line_cache[175][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24876_ (.CLK(clknet_leaf_164_clk_i),
    .D(net1716),
    .RESET_B(net360),
    .Q(\line_cache[175][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24877_ (.CLK(clknet_leaf_155_clk_i),
    .D(net642),
    .RESET_B(net363),
    .Q(\line_cache[175][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24878_ (.CLK(clknet_leaf_155_clk_i),
    .D(net1092),
    .RESET_B(net367),
    .Q(\line_cache[175][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24879_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00672_),
    .RESET_B(net351),
    .Q(\line_cache[176][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24880_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00673_),
    .RESET_B(net345),
    .Q(\line_cache[176][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24881_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00674_),
    .RESET_B(net348),
    .Q(\line_cache[176][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24882_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00675_),
    .RESET_B(net345),
    .Q(\line_cache[176][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24883_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00676_),
    .RESET_B(net348),
    .Q(\line_cache[176][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24884_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00677_),
    .RESET_B(net345),
    .Q(\line_cache[176][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24885_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00678_),
    .RESET_B(net345),
    .Q(\line_cache[176][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24886_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00679_),
    .RESET_B(net345),
    .Q(\line_cache[176][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24887_ (.CLK(clknet_leaf_180_clk_i),
    .D(net928),
    .RESET_B(net345),
    .Q(\line_cache[177][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24888_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00681_),
    .RESET_B(net346),
    .Q(\line_cache[177][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24889_ (.CLK(clknet_leaf_178_clk_i),
    .D(net814),
    .RESET_B(net346),
    .Q(\line_cache[177][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24890_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00683_),
    .RESET_B(net346),
    .Q(\line_cache[177][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24891_ (.CLK(clknet_leaf_178_clk_i),
    .D(net1074),
    .RESET_B(net346),
    .Q(\line_cache[177][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24892_ (.CLK(clknet_leaf_176_clk_i),
    .D(_00685_),
    .RESET_B(net347),
    .Q(\line_cache[177][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24893_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00686_),
    .RESET_B(net346),
    .Q(\line_cache[177][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24894_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00687_),
    .RESET_B(net345),
    .Q(\line_cache[177][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24895_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00688_),
    .RESET_B(net349),
    .Q(\line_cache[178][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24896_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00689_),
    .RESET_B(net349),
    .Q(\line_cache[178][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24897_ (.CLK(clknet_leaf_178_clk_i),
    .D(_00690_),
    .RESET_B(net346),
    .Q(\line_cache[178][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24898_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00691_),
    .RESET_B(net325),
    .Q(\line_cache[178][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24899_ (.CLK(clknet_leaf_178_clk_i),
    .D(net1392),
    .RESET_B(net346),
    .Q(\line_cache[178][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24900_ (.CLK(clknet_leaf_177_clk_i),
    .D(net1034),
    .RESET_B(net345),
    .Q(\line_cache[178][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24901_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00694_),
    .RESET_B(net345),
    .Q(\line_cache[178][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24902_ (.CLK(clknet_leaf_187_clk_i),
    .D(net1494),
    .RESET_B(net345),
    .Q(\line_cache[178][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24903_ (.CLK(clknet_leaf_186_clk_i),
    .D(net1774),
    .RESET_B(net325),
    .Q(\line_cache[179][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24904_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00697_),
    .RESET_B(net349),
    .Q(\line_cache[179][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24905_ (.CLK(clknet_leaf_178_clk_i),
    .D(net1318),
    .RESET_B(net346),
    .Q(\line_cache[179][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24906_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00699_),
    .RESET_B(net325),
    .Q(\line_cache[179][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24907_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00700_),
    .RESET_B(net348),
    .Q(\line_cache[179][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24908_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00701_),
    .RESET_B(net347),
    .Q(\line_cache[179][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24909_ (.CLK(clknet_leaf_177_clk_i),
    .D(_00702_),
    .RESET_B(net345),
    .Q(\line_cache[179][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24910_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00703_),
    .RESET_B(net345),
    .Q(\line_cache[179][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24911_ (.CLK(clknet_leaf_184_clk_i),
    .D(net2508),
    .RESET_B(net326),
    .Q(\line_cache[180][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24912_ (.CLK(clknet_leaf_181_clk_i),
    .D(net726),
    .RESET_B(net349),
    .Q(\line_cache[180][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24913_ (.CLK(clknet_leaf_184_clk_i),
    .D(net2645),
    .RESET_B(net330),
    .Q(\line_cache[180][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24914_ (.CLK(clknet_leaf_128_clk_i),
    .D(_00715_),
    .RESET_B(net330),
    .Q(\line_cache[180][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24915_ (.CLK(clknet_leaf_183_clk_i),
    .D(net1613),
    .RESET_B(net330),
    .Q(\line_cache[180][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24916_ (.CLK(clknet_leaf_183_clk_i),
    .D(net1454),
    .RESET_B(net330),
    .Q(\line_cache[180][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24917_ (.CLK(clknet_leaf_184_clk_i),
    .D(net3885),
    .RESET_B(net330),
    .Q(\line_cache[180][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24918_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00719_),
    .RESET_B(net330),
    .Q(\line_cache[180][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24919_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00720_),
    .RESET_B(net349),
    .Q(\line_cache[181][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24920_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00721_),
    .RESET_B(net349),
    .Q(\line_cache[181][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24921_ (.CLK(clknet_leaf_184_clk_i),
    .D(net1370),
    .RESET_B(net349),
    .Q(\line_cache[181][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24922_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00723_),
    .RESET_B(net330),
    .Q(\line_cache[181][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24923_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00724_),
    .RESET_B(net331),
    .Q(\line_cache[181][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24924_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00725_),
    .RESET_B(net331),
    .Q(\line_cache[181][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24925_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00726_),
    .RESET_B(net328),
    .Q(\line_cache[181][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24926_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00727_),
    .RESET_B(net330),
    .Q(\line_cache[181][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24927_ (.CLK(clknet_leaf_180_clk_i),
    .D(net1184),
    .RESET_B(net349),
    .Q(\line_cache[182][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24928_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00729_),
    .RESET_B(net349),
    .Q(\line_cache[182][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24929_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00730_),
    .RESET_B(net349),
    .Q(\line_cache[182][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24930_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00731_),
    .RESET_B(net330),
    .Q(\line_cache[182][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24931_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00732_),
    .RESET_B(net330),
    .Q(\line_cache[182][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24932_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00733_),
    .RESET_B(net350),
    .Q(\line_cache[182][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24933_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00734_),
    .RESET_B(net330),
    .Q(\line_cache[182][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24934_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00735_),
    .RESET_B(net330),
    .Q(\line_cache[182][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24935_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00736_),
    .RESET_B(net326),
    .Q(\line_cache[183][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24936_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00737_),
    .RESET_B(net349),
    .Q(\line_cache[183][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24937_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00738_),
    .RESET_B(net349),
    .Q(\line_cache[183][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24938_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00739_),
    .RESET_B(net330),
    .Q(\line_cache[183][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24939_ (.CLK(clknet_leaf_184_clk_i),
    .D(net2450),
    .RESET_B(net330),
    .Q(\line_cache[183][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24940_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00741_),
    .RESET_B(net350),
    .Q(\line_cache[183][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24941_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00742_),
    .RESET_B(net330),
    .Q(\line_cache[183][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24942_ (.CLK(clknet_leaf_184_clk_i),
    .D(net2414),
    .RESET_B(net330),
    .Q(\line_cache[183][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24943_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00744_),
    .RESET_B(net326),
    .Q(\line_cache[184][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24944_ (.CLK(clknet_leaf_187_clk_i),
    .D(net2014),
    .RESET_B(net325),
    .Q(\line_cache[184][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24945_ (.CLK(clknet_leaf_186_clk_i),
    .D(net2284),
    .RESET_B(net326),
    .Q(\line_cache[184][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24946_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00747_),
    .RESET_B(net326),
    .Q(\line_cache[184][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24947_ (.CLK(clknet_leaf_186_clk_i),
    .D(net2067),
    .RESET_B(net325),
    .Q(\line_cache[184][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24948_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00749_),
    .RESET_B(net325),
    .Q(\line_cache[184][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24949_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00750_),
    .RESET_B(net324),
    .Q(\line_cache[184][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24950_ (.CLK(clknet_leaf_188_clk_i),
    .D(net806),
    .RESET_B(net325),
    .Q(\line_cache[184][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24951_ (.CLK(clknet_leaf_199_clk_i),
    .D(net1372),
    .RESET_B(net282),
    .Q(\line_cache[185][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24952_ (.CLK(clknet_leaf_188_clk_i),
    .D(net1811),
    .RESET_B(net325),
    .Q(\line_cache[185][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24953_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00754_),
    .RESET_B(net324),
    .Q(\line_cache[185][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24954_ (.CLK(clknet_leaf_186_clk_i),
    .D(net2246),
    .RESET_B(net326),
    .Q(\line_cache[185][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24955_ (.CLK(clknet_leaf_187_clk_i),
    .D(net1790),
    .RESET_B(net325),
    .Q(\line_cache[185][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24956_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00757_),
    .RESET_B(net325),
    .Q(\line_cache[185][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24957_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00758_),
    .RESET_B(net326),
    .Q(\line_cache[185][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24958_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00759_),
    .RESET_B(net325),
    .Q(\line_cache[185][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24959_ (.CLK(clknet_leaf_199_clk_i),
    .D(net468),
    .RESET_B(net280),
    .Q(\line_cache[186][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24960_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00761_),
    .RESET_B(net325),
    .Q(\line_cache[186][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24961_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00762_),
    .RESET_B(net324),
    .Q(\line_cache[186][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24962_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00763_),
    .RESET_B(net325),
    .Q(\line_cache[186][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24963_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00764_),
    .RESET_B(net326),
    .Q(\line_cache[186][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24964_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00765_),
    .RESET_B(net282),
    .Q(\line_cache[186][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24965_ (.CLK(clknet_leaf_186_clk_i),
    .D(net2112),
    .RESET_B(net326),
    .Q(\line_cache[186][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24966_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00767_),
    .RESET_B(net282),
    .Q(\line_cache[186][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24967_ (.CLK(clknet_leaf_190_clk_i),
    .D(net1498),
    .RESET_B(net324),
    .Q(\line_cache[187][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24968_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00769_),
    .RESET_B(net325),
    .Q(\line_cache[187][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24969_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00770_),
    .RESET_B(net280),
    .Q(\line_cache[187][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24970_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00771_),
    .RESET_B(net326),
    .Q(\line_cache[187][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24971_ (.CLK(clknet_leaf_186_clk_i),
    .D(net2214),
    .RESET_B(net326),
    .Q(\line_cache[187][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24972_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00773_),
    .RESET_B(net282),
    .Q(\line_cache[187][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24973_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00774_),
    .RESET_B(net325),
    .Q(\line_cache[187][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24974_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00775_),
    .RESET_B(net282),
    .Q(\line_cache[187][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24975_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00776_),
    .RESET_B(net324),
    .Q(\line_cache[188][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24976_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00777_),
    .RESET_B(net324),
    .Q(\line_cache[188][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24977_ (.CLK(clknet_leaf_189_clk_i),
    .D(net950),
    .RESET_B(net324),
    .Q(\line_cache[188][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24978_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00779_),
    .RESET_B(net317),
    .Q(\line_cache[188][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24979_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00780_),
    .RESET_B(net324),
    .Q(\line_cache[188][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24980_ (.CLK(clknet_leaf_191_clk_i),
    .D(net1592),
    .RESET_B(net324),
    .Q(\line_cache[188][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24981_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00782_),
    .RESET_B(net283),
    .Q(\line_cache[188][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24982_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00783_),
    .RESET_B(net283),
    .Q(\line_cache[188][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24983_ (.CLK(clknet_leaf_190_clk_i),
    .D(net1256),
    .RESET_B(net327),
    .Q(\line_cache[189][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24984_ (.CLK(clknet_leaf_190_clk_i),
    .D(net1150),
    .RESET_B(net317),
    .Q(\line_cache[189][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24985_ (.CLK(clknet_leaf_188_clk_i),
    .D(net420),
    .RESET_B(net324),
    .Q(\line_cache[189][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24986_ (.CLK(clknet_leaf_191_clk_i),
    .D(_00787_),
    .RESET_B(net327),
    .Q(\line_cache[189][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24987_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00788_),
    .RESET_B(net327),
    .Q(\line_cache[189][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24988_ (.CLK(clknet_leaf_191_clk_i),
    .D(_00789_),
    .RESET_B(net317),
    .Q(\line_cache[189][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24989_ (.CLK(clknet_leaf_189_clk_i),
    .D(net846),
    .RESET_B(net324),
    .Q(\line_cache[189][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24990_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00791_),
    .RESET_B(net324),
    .Q(\line_cache[189][7] ));
 sky130_fd_sc_hd__dfrtp_1 _24991_ (.CLK(clknet_leaf_190_clk_i),
    .D(net2055),
    .RESET_B(net318),
    .Q(\line_cache[190][0] ));
 sky130_fd_sc_hd__dfrtp_1 _24992_ (.CLK(clknet_leaf_121_clk_i),
    .D(_00801_),
    .RESET_B(net318),
    .Q(\line_cache[190][1] ));
 sky130_fd_sc_hd__dfrtp_1 _24993_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00802_),
    .RESET_B(net328),
    .Q(\line_cache[190][2] ));
 sky130_fd_sc_hd__dfrtp_1 _24994_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00803_),
    .RESET_B(net274),
    .Q(\line_cache[190][3] ));
 sky130_fd_sc_hd__dfrtp_1 _24995_ (.CLK(clknet_leaf_190_clk_i),
    .D(net1931),
    .RESET_B(net327),
    .Q(\line_cache[190][4] ));
 sky130_fd_sc_hd__dfrtp_1 _24996_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00805_),
    .RESET_B(net324),
    .Q(\line_cache[190][5] ));
 sky130_fd_sc_hd__dfrtp_1 _24997_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00806_),
    .RESET_B(net324),
    .Q(\line_cache[190][6] ));
 sky130_fd_sc_hd__dfrtp_1 _24998_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00807_),
    .RESET_B(net283),
    .Q(\line_cache[190][7] ));
 sky130_fd_sc_hd__dfrtp_2 _24999_ (.CLK(clknet_leaf_121_clk_i),
    .D(_00808_),
    .RESET_B(net321),
    .Q(\line_cache[191][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25000_ (.CLK(clknet_leaf_121_clk_i),
    .D(_00809_),
    .RESET_B(net318),
    .Q(\line_cache[191][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25001_ (.CLK(clknet_leaf_185_clk_i),
    .D(net1380),
    .RESET_B(net327),
    .Q(\line_cache[191][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25002_ (.CLK(clknet_leaf_191_clk_i),
    .D(net944),
    .RESET_B(net317),
    .Q(\line_cache[191][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25003_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00812_),
    .RESET_B(net327),
    .Q(\line_cache[191][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25004_ (.CLK(clknet_leaf_191_clk_i),
    .D(_00813_),
    .RESET_B(net317),
    .Q(\line_cache[191][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25005_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00814_),
    .RESET_B(net324),
    .Q(\line_cache[191][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25006_ (.CLK(clknet_leaf_189_clk_i),
    .D(net2045),
    .RESET_B(net324),
    .Q(\line_cache[191][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25007_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00816_),
    .RESET_B(net247),
    .Q(\line_cache[192][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25008_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00817_),
    .RESET_B(net249),
    .Q(\line_cache[192][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25009_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00818_),
    .RESET_B(net249),
    .Q(\line_cache[192][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25010_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00819_),
    .RESET_B(net249),
    .Q(\line_cache[192][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25011_ (.CLK(clknet_leaf_99_clk_i),
    .D(_00820_),
    .RESET_B(net245),
    .Q(\line_cache[192][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25012_ (.CLK(clknet_leaf_99_clk_i),
    .D(_00821_),
    .RESET_B(net246),
    .Q(\line_cache[192][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25013_ (.CLK(clknet_leaf_97_clk_i),
    .D(net3236),
    .RESET_B(net250),
    .Q(\line_cache[192][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25014_ (.CLK(clknet_leaf_96_clk_i),
    .D(net3252),
    .RESET_B(net250),
    .Q(\line_cache[192][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25015_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00824_),
    .RESET_B(net247),
    .Q(\line_cache[193][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25016_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00825_),
    .RESET_B(net249),
    .Q(\line_cache[193][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25017_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00826_),
    .RESET_B(net249),
    .Q(\line_cache[193][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25018_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00827_),
    .RESET_B(net249),
    .Q(\line_cache[193][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25019_ (.CLK(clknet_leaf_99_clk_i),
    .D(_00828_),
    .RESET_B(net246),
    .Q(\line_cache[193][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25020_ (.CLK(clknet_leaf_95_clk_i),
    .D(_00829_),
    .RESET_B(net249),
    .Q(\line_cache[193][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25021_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00830_),
    .RESET_B(net250),
    .Q(\line_cache[193][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25022_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00831_),
    .RESET_B(net250),
    .Q(\line_cache[193][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25023_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00832_),
    .RESET_B(net247),
    .Q(\line_cache[194][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25024_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00833_),
    .RESET_B(net250),
    .Q(\line_cache[194][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25025_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00834_),
    .RESET_B(net250),
    .Q(\line_cache[194][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25026_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00835_),
    .RESET_B(net250),
    .Q(\line_cache[194][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25027_ (.CLK(clknet_leaf_98_clk_i),
    .D(_00836_),
    .RESET_B(net250),
    .Q(\line_cache[194][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25028_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00837_),
    .RESET_B(net248),
    .Q(\line_cache[194][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25029_ (.CLK(clknet_leaf_100_clk_i),
    .D(_00838_),
    .RESET_B(net248),
    .Q(\line_cache[194][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25030_ (.CLK(clknet_leaf_97_clk_i),
    .D(_00839_),
    .RESET_B(net250),
    .Q(\line_cache[194][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25031_ (.CLK(clknet_leaf_136_clk_i),
    .D(_00840_),
    .RESET_B(net332),
    .Q(\line_cache[195][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25032_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00841_),
    .RESET_B(net335),
    .Q(\line_cache[195][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25033_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00842_),
    .RESET_B(net335),
    .Q(\line_cache[195][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25034_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00843_),
    .RESET_B(net250),
    .Q(\line_cache[195][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25035_ (.CLK(clknet_leaf_136_clk_i),
    .D(_00844_),
    .RESET_B(net332),
    .Q(\line_cache[195][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25036_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00845_),
    .RESET_B(net250),
    .Q(\line_cache[195][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25037_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00846_),
    .RESET_B(net335),
    .Q(\line_cache[195][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25038_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00847_),
    .RESET_B(net250),
    .Q(\line_cache[195][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25039_ (.CLK(clknet_leaf_136_clk_i),
    .D(net1472),
    .RESET_B(net332),
    .Q(\line_cache[196][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25040_ (.CLK(clknet_leaf_96_clk_i),
    .D(_00849_),
    .RESET_B(net335),
    .Q(\line_cache[196][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25041_ (.CLK(clknet_leaf_136_clk_i),
    .D(net2587),
    .RESET_B(net332),
    .Q(\line_cache[196][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25042_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00851_),
    .RESET_B(net335),
    .Q(\line_cache[196][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25043_ (.CLK(clknet_leaf_135_clk_i),
    .D(net1540),
    .RESET_B(net332),
    .Q(\line_cache[196][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25044_ (.CLK(clknet_leaf_137_clk_i),
    .D(net2708),
    .RESET_B(net333),
    .Q(\line_cache[196][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25045_ (.CLK(clknet_leaf_139_clk_i),
    .D(net3552),
    .RESET_B(net335),
    .Q(\line_cache[196][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25046_ (.CLK(clknet_leaf_139_clk_i),
    .D(net3695),
    .RESET_B(net335),
    .Q(\line_cache[196][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25047_ (.CLK(clknet_leaf_136_clk_i),
    .D(net432),
    .RESET_B(net332),
    .Q(\line_cache[197][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25048_ (.CLK(clknet_leaf_138_clk_i),
    .D(net2460),
    .RESET_B(net335),
    .Q(\line_cache[197][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25049_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00858_),
    .RESET_B(net335),
    .Q(\line_cache[197][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25050_ (.CLK(clknet_leaf_138_clk_i),
    .D(net2259),
    .RESET_B(net335),
    .Q(\line_cache[197][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25051_ (.CLK(clknet_leaf_137_clk_i),
    .D(_00860_),
    .RESET_B(net333),
    .Q(\line_cache[197][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25052_ (.CLK(clknet_leaf_139_clk_i),
    .D(_00861_),
    .RESET_B(net335),
    .Q(\line_cache[197][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25053_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00862_),
    .RESET_B(net335),
    .Q(\line_cache[197][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25054_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00863_),
    .RESET_B(net335),
    .Q(\line_cache[197][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25055_ (.CLK(clknet_leaf_136_clk_i),
    .D(_00864_),
    .RESET_B(net334),
    .Q(\line_cache[198][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25056_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00865_),
    .RESET_B(net343),
    .Q(\line_cache[198][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25057_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00866_),
    .RESET_B(net343),
    .Q(\line_cache[198][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25058_ (.CLK(clknet_leaf_138_clk_i),
    .D(net1244),
    .RESET_B(net336),
    .Q(\line_cache[198][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25059_ (.CLK(clknet_leaf_136_clk_i),
    .D(net872),
    .RESET_B(net334),
    .Q(\line_cache[198][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25060_ (.CLK(clknet_leaf_138_clk_i),
    .D(net1760),
    .RESET_B(net335),
    .Q(\line_cache[198][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25061_ (.CLK(clknet_leaf_138_clk_i),
    .D(net2242),
    .RESET_B(net335),
    .Q(\line_cache[198][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25062_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00871_),
    .RESET_B(net335),
    .Q(\line_cache[198][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25063_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00872_),
    .RESET_B(net336),
    .Q(\line_cache[199][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25064_ (.CLK(clknet_leaf_138_clk_i),
    .D(_00873_),
    .RESET_B(net336),
    .Q(\line_cache[199][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25065_ (.CLK(clknet_leaf_137_clk_i),
    .D(net1664),
    .RESET_B(net333),
    .Q(\line_cache[199][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25066_ (.CLK(clknet_leaf_132_clk_i),
    .D(net2664),
    .RESET_B(net333),
    .Q(\line_cache[199][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25067_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00876_),
    .RESET_B(net336),
    .Q(\line_cache[199][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25068_ (.CLK(clknet_leaf_141_clk_i),
    .D(_00877_),
    .RESET_B(net336),
    .Q(\line_cache[199][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25069_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00878_),
    .RESET_B(net336),
    .Q(\line_cache[199][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25070_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00879_),
    .RESET_B(net336),
    .Q(\line_cache[199][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25071_ (.CLK(clknet_leaf_137_clk_i),
    .D(net1286),
    .RESET_B(net333),
    .Q(\line_cache[200][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25072_ (.CLK(clknet_leaf_140_clk_i),
    .D(_00897_),
    .RESET_B(net336),
    .Q(\line_cache[200][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25073_ (.CLK(clknet_leaf_137_clk_i),
    .D(net1779),
    .RESET_B(net333),
    .Q(\line_cache[200][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25074_ (.CLK(clknet_leaf_141_clk_i),
    .D(_00899_),
    .RESET_B(net336),
    .Q(\line_cache[200][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25075_ (.CLK(clknet_leaf_141_clk_i),
    .D(_00900_),
    .RESET_B(net336),
    .Q(\line_cache[200][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25076_ (.CLK(clknet_leaf_137_clk_i),
    .D(net2647),
    .RESET_B(net333),
    .Q(\line_cache[200][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25077_ (.CLK(clknet_leaf_138_clk_i),
    .D(net3761),
    .RESET_B(net336),
    .Q(\line_cache[200][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25078_ (.CLK(clknet_leaf_138_clk_i),
    .D(net3771),
    .RESET_B(net336),
    .Q(\line_cache[200][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25079_ (.CLK(clknet_leaf_132_clk_i),
    .D(_00904_),
    .RESET_B(net334),
    .Q(\line_cache[201][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25080_ (.CLK(clknet_leaf_138_clk_i),
    .D(net2376),
    .RESET_B(net336),
    .Q(\line_cache[201][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25081_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00906_),
    .RESET_B(net336),
    .Q(\line_cache[201][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25082_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00907_),
    .RESET_B(net341),
    .Q(\line_cache[201][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25083_ (.CLK(clknet_leaf_132_clk_i),
    .D(net1036),
    .RESET_B(net334),
    .Q(\line_cache[201][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25084_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00909_),
    .RESET_B(net336),
    .Q(\line_cache[201][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25085_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00910_),
    .RESET_B(net341),
    .Q(\line_cache[201][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25086_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00911_),
    .RESET_B(net343),
    .Q(\line_cache[201][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25087_ (.CLK(clknet_leaf_137_clk_i),
    .D(net1112),
    .RESET_B(net334),
    .Q(\line_cache[202][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25088_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00913_),
    .RESET_B(net341),
    .Q(\line_cache[202][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25089_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00914_),
    .RESET_B(net341),
    .Q(\line_cache[202][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25090_ (.CLK(clknet_leaf_141_clk_i),
    .D(net1336),
    .RESET_B(net341),
    .Q(\line_cache[202][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25091_ (.CLK(clknet_leaf_132_clk_i),
    .D(net1950),
    .RESET_B(net334),
    .Q(\line_cache[202][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25092_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00917_),
    .RESET_B(net336),
    .Q(\line_cache[202][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25093_ (.CLK(clknet_leaf_137_clk_i),
    .D(net2381),
    .RESET_B(net334),
    .Q(\line_cache[202][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25094_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00919_),
    .RESET_B(net341),
    .Q(\line_cache[202][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25095_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00920_),
    .RESET_B(net342),
    .Q(\line_cache[203][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25096_ (.CLK(clknet_leaf_142_clk_i),
    .D(net704),
    .RESET_B(net341),
    .Q(\line_cache[203][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25097_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00922_),
    .RESET_B(net341),
    .Q(\line_cache[203][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25098_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00923_),
    .RESET_B(net342),
    .Q(\line_cache[203][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25099_ (.CLK(clknet_leaf_132_clk_i),
    .D(net1294),
    .RESET_B(net334),
    .Q(\line_cache[203][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25100_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00925_),
    .RESET_B(net341),
    .Q(\line_cache[203][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25101_ (.CLK(clknet_leaf_131_clk_i),
    .D(net438),
    .RESET_B(net337),
    .Q(\line_cache[203][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25102_ (.CLK(clknet_leaf_142_clk_i),
    .D(_00927_),
    .RESET_B(net341),
    .Q(\line_cache[203][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25103_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00928_),
    .RESET_B(net337),
    .Q(\line_cache[204][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25104_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00929_),
    .RESET_B(net341),
    .Q(\line_cache[204][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25105_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00930_),
    .RESET_B(net341),
    .Q(\line_cache[204][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25106_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00931_),
    .RESET_B(net337),
    .Q(\line_cache[204][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25107_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00932_),
    .RESET_B(net338),
    .Q(\line_cache[204][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25108_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00933_),
    .RESET_B(net338),
    .Q(\line_cache[204][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25109_ (.CLK(clknet_leaf_133_clk_i),
    .D(_00934_),
    .RESET_B(net337),
    .Q(\line_cache[204][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25110_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00935_),
    .RESET_B(net338),
    .Q(\line_cache[204][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25111_ (.CLK(clknet_leaf_144_clk_i),
    .D(_00936_),
    .RESET_B(net339),
    .Q(\line_cache[205][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25112_ (.CLK(clknet_leaf_142_clk_i),
    .D(net2114),
    .RESET_B(net341),
    .Q(\line_cache[205][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25113_ (.CLK(clknet_leaf_144_clk_i),
    .D(net1456),
    .RESET_B(net342),
    .Q(\line_cache[205][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25114_ (.CLK(clknet_leaf_144_clk_i),
    .D(net1058),
    .RESET_B(net341),
    .Q(\line_cache[205][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25115_ (.CLK(clknet_leaf_132_clk_i),
    .D(net2147),
    .RESET_B(net338),
    .Q(\line_cache[205][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25116_ (.CLK(clknet_leaf_130_clk_i),
    .D(_00941_),
    .RESET_B(net337),
    .Q(\line_cache[205][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25117_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00942_),
    .RESET_B(net338),
    .Q(\line_cache[205][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25118_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00943_),
    .RESET_B(net338),
    .Q(\line_cache[205][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25119_ (.CLK(clknet_leaf_145_clk_i),
    .D(net496),
    .RESET_B(net339),
    .Q(\line_cache[206][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25120_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00945_),
    .RESET_B(net338),
    .Q(\line_cache[206][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25121_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00946_),
    .RESET_B(net338),
    .Q(\line_cache[206][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25122_ (.CLK(clknet_leaf_143_clk_i),
    .D(net824),
    .RESET_B(net342),
    .Q(\line_cache[206][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25123_ (.CLK(clknet_leaf_132_clk_i),
    .D(net530),
    .RESET_B(net338),
    .Q(\line_cache[206][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25124_ (.CLK(clknet_leaf_142_clk_i),
    .D(net982),
    .RESET_B(net341),
    .Q(\line_cache[206][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25125_ (.CLK(clknet_leaf_130_clk_i),
    .D(_00950_),
    .RESET_B(net337),
    .Q(\line_cache[206][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25126_ (.CLK(clknet_leaf_142_clk_i),
    .D(net998),
    .RESET_B(net341),
    .Q(\line_cache[206][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25127_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00952_),
    .RESET_B(net339),
    .Q(\line_cache[207][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25128_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00953_),
    .RESET_B(net342),
    .Q(\line_cache[207][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25129_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00954_),
    .RESET_B(net342),
    .Q(\line_cache[207][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25130_ (.CLK(clknet_leaf_143_clk_i),
    .D(net2336),
    .RESET_B(net342),
    .Q(\line_cache[207][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25131_ (.CLK(clknet_leaf_145_clk_i),
    .D(net2002),
    .RESET_B(net340),
    .Q(\line_cache[207][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25132_ (.CLK(clknet_leaf_129_clk_i),
    .D(_00957_),
    .RESET_B(net339),
    .Q(\line_cache[207][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25133_ (.CLK(clknet_leaf_131_clk_i),
    .D(_00958_),
    .RESET_B(net339),
    .Q(\line_cache[207][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25134_ (.CLK(clknet_leaf_145_clk_i),
    .D(net2080),
    .RESET_B(net340),
    .Q(\line_cache[207][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25135_ (.CLK(clknet_leaf_145_clk_i),
    .D(net1944),
    .RESET_B(net340),
    .Q(\line_cache[208][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25136_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00961_),
    .RESET_B(net342),
    .Q(\line_cache[208][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25137_ (.CLK(clknet_leaf_143_clk_i),
    .D(net2324),
    .RESET_B(net342),
    .Q(\line_cache[208][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25138_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00963_),
    .RESET_B(net342),
    .Q(\line_cache[208][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25139_ (.CLK(clknet_leaf_146_clk_i),
    .D(net1683),
    .RESET_B(net340),
    .Q(\line_cache[208][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25140_ (.CLK(clknet_leaf_146_clk_i),
    .D(net1426),
    .RESET_B(net339),
    .Q(\line_cache[208][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25141_ (.CLK(clknet_leaf_145_clk_i),
    .D(_00966_),
    .RESET_B(net340),
    .Q(\line_cache[208][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25142_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00967_),
    .RESET_B(net342),
    .Q(\line_cache[208][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25143_ (.CLK(clknet_leaf_145_clk_i),
    .D(net1440),
    .RESET_B(net340),
    .Q(\line_cache[209][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25144_ (.CLK(clknet_leaf_143_clk_i),
    .D(net2452),
    .RESET_B(net366),
    .Q(\line_cache[209][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25145_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00970_),
    .RESET_B(net366),
    .Q(\line_cache[209][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25146_ (.CLK(clknet_leaf_151_clk_i),
    .D(net2488),
    .RESET_B(net366),
    .Q(\line_cache[209][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25147_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00972_),
    .RESET_B(net366),
    .Q(\line_cache[209][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25148_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00973_),
    .RESET_B(net342),
    .Q(\line_cache[209][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25149_ (.CLK(clknet_leaf_146_clk_i),
    .D(net1818),
    .RESET_B(net339),
    .Q(\line_cache[209][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25150_ (.CLK(clknet_leaf_143_clk_i),
    .D(_00975_),
    .RESET_B(net342),
    .Q(\line_cache[209][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25151_ (.CLK(clknet_leaf_145_clk_i),
    .D(net1978),
    .RESET_B(net340),
    .Q(\line_cache[210][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25152_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00985_),
    .RESET_B(net366),
    .Q(\line_cache[210][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25153_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00986_),
    .RESET_B(net366),
    .Q(\line_cache[210][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25154_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00987_),
    .RESET_B(net366),
    .Q(\line_cache[210][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25155_ (.CLK(clknet_leaf_149_clk_i),
    .D(net1076),
    .RESET_B(net362),
    .Q(\line_cache[210][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25156_ (.CLK(clknet_leaf_143_clk_i),
    .D(net1963),
    .RESET_B(net342),
    .Q(\line_cache[210][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25157_ (.CLK(clknet_leaf_149_clk_i),
    .D(_00990_),
    .RESET_B(net340),
    .Q(\line_cache[210][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25158_ (.CLK(clknet_leaf_143_clk_i),
    .D(net1960),
    .RESET_B(net342),
    .Q(\line_cache[210][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25159_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00992_),
    .RESET_B(net366),
    .Q(\line_cache[211][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25160_ (.CLK(clknet_leaf_148_clk_i),
    .D(net446),
    .RESET_B(net362),
    .Q(\line_cache[211][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25161_ (.CLK(clknet_leaf_151_clk_i),
    .D(net1234),
    .RESET_B(net366),
    .Q(\line_cache[211][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25162_ (.CLK(clknet_leaf_151_clk_i),
    .D(net1054),
    .RESET_B(net366),
    .Q(\line_cache[211][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25163_ (.CLK(clknet_leaf_147_clk_i),
    .D(net720),
    .RESET_B(net362),
    .Q(\line_cache[211][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25164_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00997_),
    .RESET_B(net366),
    .Q(\line_cache[211][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25165_ (.CLK(clknet_leaf_145_clk_i),
    .D(net466),
    .RESET_B(net362),
    .Q(\line_cache[211][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25166_ (.CLK(clknet_leaf_147_clk_i),
    .D(net560),
    .RESET_B(net362),
    .Q(\line_cache[211][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25167_ (.CLK(clknet_leaf_149_clk_i),
    .D(net548),
    .RESET_B(net362),
    .Q(\line_cache[212][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25168_ (.CLK(clknet_leaf_159_clk_i),
    .D(net1156),
    .RESET_B(net363),
    .Q(\line_cache[212][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25169_ (.CLK(clknet_leaf_149_clk_i),
    .D(net534),
    .RESET_B(net365),
    .Q(\line_cache[212][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25170_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01003_),
    .RESET_B(net366),
    .Q(\line_cache[212][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25171_ (.CLK(clknet_leaf_159_clk_i),
    .D(net580),
    .RESET_B(net362),
    .Q(\line_cache[212][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25172_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01005_),
    .RESET_B(net364),
    .Q(\line_cache[212][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25173_ (.CLK(clknet_leaf_145_clk_i),
    .D(_01006_),
    .RESET_B(net365),
    .Q(\line_cache[212][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25174_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01007_),
    .RESET_B(net365),
    .Q(\line_cache[212][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25175_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01008_),
    .RESET_B(net364),
    .Q(\line_cache[213][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25176_ (.CLK(clknet_leaf_148_clk_i),
    .D(net556),
    .RESET_B(net362),
    .Q(\line_cache[213][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25177_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01010_),
    .RESET_B(net366),
    .Q(\line_cache[213][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25178_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01011_),
    .RESET_B(net366),
    .Q(\line_cache[213][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25179_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01012_),
    .RESET_B(net364),
    .Q(\line_cache[213][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25180_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01013_),
    .RESET_B(net366),
    .Q(\line_cache[213][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25181_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01014_),
    .RESET_B(net365),
    .Q(\line_cache[213][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25182_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01015_),
    .RESET_B(net365),
    .Q(\line_cache[213][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25183_ (.CLK(clknet_leaf_149_clk_i),
    .D(net760),
    .RESET_B(net364),
    .Q(\line_cache[214][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25184_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01017_),
    .RESET_B(net364),
    .Q(\line_cache[214][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25185_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01018_),
    .RESET_B(net364),
    .Q(\line_cache[214][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25186_ (.CLK(clknet_leaf_149_clk_i),
    .D(net456),
    .RESET_B(net365),
    .Q(\line_cache[214][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25187_ (.CLK(clknet_leaf_157_clk_i),
    .D(net602),
    .RESET_B(net363),
    .Q(\line_cache[214][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25188_ (.CLK(clknet_leaf_150_clk_i),
    .D(net450),
    .RESET_B(net364),
    .Q(\line_cache[214][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25189_ (.CLK(clknet_leaf_146_clk_i),
    .D(net1838),
    .RESET_B(net340),
    .Q(\line_cache[214][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25190_ (.CLK(clknet_leaf_148_clk_i),
    .D(net422),
    .RESET_B(net365),
    .Q(\line_cache[214][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25191_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01024_),
    .RESET_B(net362),
    .Q(\line_cache[215][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25192_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01025_),
    .RESET_B(net350),
    .Q(\line_cache[215][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25193_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01026_),
    .RESET_B(net363),
    .Q(\line_cache[215][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25194_ (.CLK(clknet_leaf_147_clk_i),
    .D(net2553),
    .RESET_B(net362),
    .Q(\line_cache[215][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25195_ (.CLK(clknet_leaf_146_clk_i),
    .D(net1940),
    .RESET_B(net362),
    .Q(\line_cache[215][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25196_ (.CLK(clknet_leaf_129_clk_i),
    .D(net2505),
    .RESET_B(net339),
    .Q(\line_cache[215][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25197_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01030_),
    .RESET_B(net363),
    .Q(\line_cache[215][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25198_ (.CLK(clknet_leaf_129_clk_i),
    .D(net1526),
    .RESET_B(net339),
    .Q(\line_cache[215][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25199_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01032_),
    .RESET_B(net362),
    .Q(\line_cache[216][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25200_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01033_),
    .RESET_B(net350),
    .Q(\line_cache[216][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25201_ (.CLK(clknet_leaf_128_clk_i),
    .D(net2061),
    .RESET_B(net331),
    .Q(\line_cache[216][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25202_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01035_),
    .RESET_B(net350),
    .Q(\line_cache[216][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25203_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01036_),
    .RESET_B(net362),
    .Q(\line_cache[216][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25204_ (.CLK(clknet_leaf_128_clk_i),
    .D(net2163),
    .RESET_B(net339),
    .Q(\line_cache[216][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25205_ (.CLK(clknet_leaf_146_clk_i),
    .D(net3659),
    .RESET_B(net362),
    .Q(\line_cache[216][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25206_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01039_),
    .RESET_B(net339),
    .Q(\line_cache[216][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25207_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01040_),
    .RESET_B(net362),
    .Q(\line_cache[217][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25208_ (.CLK(clknet_leaf_128_clk_i),
    .D(net1982),
    .RESET_B(net331),
    .Q(\line_cache[217][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25209_ (.CLK(clknet_leaf_182_clk_i),
    .D(_01042_),
    .RESET_B(net350),
    .Q(\line_cache[217][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25210_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01043_),
    .RESET_B(net350),
    .Q(\line_cache[217][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25211_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01044_),
    .RESET_B(net337),
    .Q(\line_cache[217][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25212_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01045_),
    .RESET_B(net339),
    .Q(\line_cache[217][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25213_ (.CLK(clknet_leaf_129_clk_i),
    .D(net2198),
    .RESET_B(net339),
    .Q(\line_cache[217][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25214_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01047_),
    .RESET_B(net339),
    .Q(\line_cache[217][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25215_ (.CLK(clknet_leaf_147_clk_i),
    .D(net714),
    .RESET_B(net362),
    .Q(\line_cache[218][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25216_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01049_),
    .RESET_B(net331),
    .Q(\line_cache[218][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25217_ (.CLK(clknet_leaf_183_clk_i),
    .D(_01050_),
    .RESET_B(net331),
    .Q(\line_cache[218][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25218_ (.CLK(clknet_leaf_183_clk_i),
    .D(net852),
    .RESET_B(net350),
    .Q(\line_cache[218][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25219_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01052_),
    .RESET_B(net337),
    .Q(\line_cache[218][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25220_ (.CLK(clknet_leaf_128_clk_i),
    .D(net1814),
    .RESET_B(net339),
    .Q(\line_cache[218][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25221_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01054_),
    .RESET_B(net337),
    .Q(\line_cache[218][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25222_ (.CLK(clknet_leaf_146_clk_i),
    .D(net964),
    .RESET_B(net339),
    .Q(\line_cache[218][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25223_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01056_),
    .RESET_B(net337),
    .Q(\line_cache[219][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25224_ (.CLK(clknet_leaf_126_clk_i),
    .D(net762),
    .RESET_B(net328),
    .Q(\line_cache[219][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25225_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01058_),
    .RESET_B(net337),
    .Q(\line_cache[219][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25226_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01059_),
    .RESET_B(net331),
    .Q(\line_cache[219][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25227_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01060_),
    .RESET_B(net337),
    .Q(\line_cache[219][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25228_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01061_),
    .RESET_B(net337),
    .Q(\line_cache[219][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25229_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01062_),
    .RESET_B(net328),
    .Q(\line_cache[219][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25230_ (.CLK(clknet_leaf_128_clk_i),
    .D(net2521),
    .RESET_B(net331),
    .Q(\line_cache[219][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25231_ (.CLK(clknet_leaf_127_clk_i),
    .D(net1026),
    .RESET_B(net328),
    .Q(\line_cache[220][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25232_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01073_),
    .RESET_B(net328),
    .Q(\line_cache[220][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25233_ (.CLK(clknet_leaf_127_clk_i),
    .D(net926),
    .RESET_B(net328),
    .Q(\line_cache[220][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25234_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01075_),
    .RESET_B(net328),
    .Q(\line_cache[220][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25235_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01076_),
    .RESET_B(net321),
    .Q(\line_cache[220][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25236_ (.CLK(clknet_leaf_127_clk_i),
    .D(net1805),
    .RESET_B(net328),
    .Q(\line_cache[220][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25237_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01078_),
    .RESET_B(net329),
    .Q(\line_cache[220][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25238_ (.CLK(clknet_leaf_128_clk_i),
    .D(net2047),
    .RESET_B(net331),
    .Q(\line_cache[220][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25239_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01080_),
    .RESET_B(net328),
    .Q(\line_cache[221][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25240_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01081_),
    .RESET_B(net328),
    .Q(\line_cache[221][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25241_ (.CLK(clknet_leaf_127_clk_i),
    .D(net1825),
    .RESET_B(net329),
    .Q(\line_cache[221][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25242_ (.CLK(clknet_leaf_127_clk_i),
    .D(net2227),
    .RESET_B(net329),
    .Q(\line_cache[221][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25243_ (.CLK(clknet_leaf_126_clk_i),
    .D(net1382),
    .RESET_B(net329),
    .Q(\line_cache[221][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25244_ (.CLK(clknet_leaf_184_clk_i),
    .D(_01085_),
    .RESET_B(net328),
    .Q(\line_cache[221][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25245_ (.CLK(clknet_leaf_124_clk_i),
    .D(net1679),
    .RESET_B(net329),
    .Q(\line_cache[221][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25246_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01087_),
    .RESET_B(net328),
    .Q(\line_cache[221][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25247_ (.CLK(clknet_leaf_125_clk_i),
    .D(net2760),
    .RESET_B(net321),
    .Q(\line_cache[222][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25248_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01089_),
    .RESET_B(net328),
    .Q(\line_cache[222][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25249_ (.CLK(clknet_leaf_185_clk_i),
    .D(_01090_),
    .RESET_B(net328),
    .Q(\line_cache[222][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25250_ (.CLK(clknet_leaf_128_clk_i),
    .D(net2051),
    .RESET_B(net329),
    .Q(\line_cache[222][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25251_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01092_),
    .RESET_B(net321),
    .Q(\line_cache[222][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25252_ (.CLK(clknet_leaf_129_clk_i),
    .D(net1728),
    .RESET_B(net337),
    .Q(\line_cache[222][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25253_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01094_),
    .RESET_B(net328),
    .Q(\line_cache[222][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25254_ (.CLK(clknet_leaf_128_clk_i),
    .D(net2043),
    .RESET_B(net329),
    .Q(\line_cache[222][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25255_ (.CLK(clknet_leaf_124_clk_i),
    .D(net2141),
    .RESET_B(net321),
    .Q(\line_cache[223][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25256_ (.CLK(clknet_leaf_124_clk_i),
    .D(net1574),
    .RESET_B(net321),
    .Q(\line_cache[223][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25257_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01098_),
    .RESET_B(net321),
    .Q(\line_cache[223][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25258_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01099_),
    .RESET_B(net321),
    .Q(\line_cache[223][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25259_ (.CLK(clknet_leaf_124_clk_i),
    .D(net2622),
    .RESET_B(net322),
    .Q(\line_cache[223][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25260_ (.CLK(clknet_leaf_127_clk_i),
    .D(net2122),
    .RESET_B(net322),
    .Q(\line_cache[223][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25261_ (.CLK(clknet_leaf_130_clk_i),
    .D(net1366),
    .RESET_B(net337),
    .Q(\line_cache[223][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25262_ (.CLK(clknet_leaf_124_clk_i),
    .D(net2478),
    .RESET_B(net329),
    .Q(\line_cache[223][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25263_ (.CLK(clknet_leaf_134_clk_i),
    .D(net594),
    .RESET_B(net333),
    .Q(\line_cache[224][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25264_ (.CLK(clknet_leaf_122_clk_i),
    .D(net522),
    .RESET_B(net321),
    .Q(\line_cache[224][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25265_ (.CLK(clknet_leaf_123_clk_i),
    .D(net962),
    .RESET_B(net320),
    .Q(\line_cache[224][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25266_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01107_),
    .RESET_B(net322),
    .Q(\line_cache[224][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25267_ (.CLK(clknet_leaf_123_clk_i),
    .D(net552),
    .RESET_B(net320),
    .Q(\line_cache[224][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25268_ (.CLK(clknet_leaf_124_clk_i),
    .D(net638),
    .RESET_B(net322),
    .Q(\line_cache[224][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25269_ (.CLK(clknet_leaf_130_clk_i),
    .D(net3247),
    .RESET_B(net333),
    .Q(\line_cache[224][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25270_ (.CLK(clknet_leaf_133_clk_i),
    .D(net3302),
    .RESET_B(net333),
    .Q(\line_cache[224][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25271_ (.CLK(clknet_leaf_133_clk_i),
    .D(_01112_),
    .RESET_B(net333),
    .Q(\line_cache[225][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25272_ (.CLK(clknet_leaf_123_clk_i),
    .D(net2394),
    .RESET_B(net322),
    .Q(\line_cache[225][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25273_ (.CLK(clknet_leaf_122_clk_i),
    .D(net546),
    .RESET_B(net320),
    .Q(\line_cache[225][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25274_ (.CLK(clknet_leaf_124_clk_i),
    .D(net1604),
    .RESET_B(net322),
    .Q(\line_cache[225][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25275_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01116_),
    .RESET_B(net320),
    .Q(\line_cache[225][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25276_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01117_),
    .RESET_B(net322),
    .Q(\line_cache[225][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25277_ (.CLK(clknet_leaf_134_clk_i),
    .D(net568),
    .RESET_B(net333),
    .Q(\line_cache[225][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25278_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01119_),
    .RESET_B(net322),
    .Q(\line_cache[225][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25279_ (.CLK(clknet_leaf_134_clk_i),
    .D(net512),
    .RESET_B(net333),
    .Q(\line_cache[226][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25280_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01121_),
    .RESET_B(net322),
    .Q(\line_cache[226][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25281_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01122_),
    .RESET_B(net322),
    .Q(\line_cache[226][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25282_ (.CLK(clknet_leaf_125_clk_i),
    .D(net430),
    .RESET_B(net321),
    .Q(\line_cache[226][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25283_ (.CLK(clknet_leaf_123_clk_i),
    .D(net700),
    .RESET_B(net320),
    .Q(\line_cache[226][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25284_ (.CLK(clknet_leaf_125_clk_i),
    .D(net488),
    .RESET_B(net321),
    .Q(\line_cache[226][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25285_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01126_),
    .RESET_B(net337),
    .Q(\line_cache[226][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25286_ (.CLK(clknet_leaf_133_clk_i),
    .D(net424),
    .RESET_B(net333),
    .Q(\line_cache[226][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25287_ (.CLK(clknet_leaf_134_clk_i),
    .D(net566),
    .RESET_B(net333),
    .Q(\line_cache[227][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25288_ (.CLK(clknet_leaf_132_clk_i),
    .D(_01129_),
    .RESET_B(net333),
    .Q(\line_cache[227][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25289_ (.CLK(clknet_leaf_137_clk_i),
    .D(_01130_),
    .RESET_B(net334),
    .Q(\line_cache[227][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25290_ (.CLK(clknet_leaf_134_clk_i),
    .D(net604),
    .RESET_B(net332),
    .Q(\line_cache[227][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25291_ (.CLK(clknet_leaf_134_clk_i),
    .D(net738),
    .RESET_B(net332),
    .Q(\line_cache[227][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25292_ (.CLK(clknet_leaf_134_clk_i),
    .D(net674),
    .RESET_B(net332),
    .Q(\line_cache[227][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25293_ (.CLK(clknet_leaf_134_clk_i),
    .D(net1559),
    .RESET_B(net323),
    .Q(\line_cache[227][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25294_ (.CLK(clknet_leaf_135_clk_i),
    .D(net686),
    .RESET_B(net332),
    .Q(\line_cache[227][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25295_ (.CLK(clknet_leaf_134_clk_i),
    .D(net1246),
    .RESET_B(net332),
    .Q(\line_cache[228][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25296_ (.CLK(clknet_leaf_135_clk_i),
    .D(net440),
    .RESET_B(net334),
    .Q(\line_cache[228][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25297_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01138_),
    .RESET_B(net248),
    .Q(\line_cache[228][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25298_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01139_),
    .RESET_B(net248),
    .Q(\line_cache[228][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25299_ (.CLK(clknet_leaf_102_clk_i),
    .D(net588),
    .RESET_B(net332),
    .Q(\line_cache[228][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25300_ (.CLK(clknet_leaf_101_clk_i),
    .D(net596),
    .RESET_B(net247),
    .Q(\line_cache[228][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25301_ (.CLK(clknet_leaf_101_clk_i),
    .D(net3664),
    .RESET_B(net247),
    .Q(\line_cache[228][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25302_ (.CLK(clknet_leaf_101_clk_i),
    .D(net3393),
    .RESET_B(net247),
    .Q(\line_cache[228][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25303_ (.CLK(clknet_leaf_134_clk_i),
    .D(net482),
    .RESET_B(net332),
    .Q(\line_cache[229][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25304_ (.CLK(clknet_leaf_135_clk_i),
    .D(net708),
    .RESET_B(net332),
    .Q(\line_cache[229][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25305_ (.CLK(clknet_leaf_135_clk_i),
    .D(net426),
    .RESET_B(net334),
    .Q(\line_cache[229][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25306_ (.CLK(clknet_leaf_135_clk_i),
    .D(net620),
    .RESET_B(net334),
    .Q(\line_cache[229][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25307_ (.CLK(clknet_leaf_135_clk_i),
    .D(net520),
    .RESET_B(net332),
    .Q(\line_cache[229][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25308_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01149_),
    .RESET_B(net248),
    .Q(\line_cache[229][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25309_ (.CLK(clknet_leaf_101_clk_i),
    .D(net646),
    .RESET_B(net247),
    .Q(\line_cache[229][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25310_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01151_),
    .RESET_B(net248),
    .Q(\line_cache[229][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25311_ (.CLK(clknet_leaf_134_clk_i),
    .D(net494),
    .RESET_B(net332),
    .Q(\line_cache[230][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25312_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01161_),
    .RESET_B(net248),
    .Q(\line_cache[230][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25313_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01162_),
    .RESET_B(net248),
    .Q(\line_cache[230][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25314_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01163_),
    .RESET_B(net248),
    .Q(\line_cache[230][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25315_ (.CLK(clknet_leaf_102_clk_i),
    .D(net1084),
    .RESET_B(net247),
    .Q(\line_cache[230][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25316_ (.CLK(clknet_leaf_101_clk_i),
    .D(net776),
    .RESET_B(net247),
    .Q(\line_cache[230][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25317_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01166_),
    .RESET_B(net247),
    .Q(\line_cache[230][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25318_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01167_),
    .RESET_B(net246),
    .Q(\line_cache[230][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25319_ (.CLK(clknet_leaf_102_clk_i),
    .D(net670),
    .RESET_B(net247),
    .Q(\line_cache[231][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25320_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01169_),
    .RESET_B(net247),
    .Q(\line_cache[231][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25321_ (.CLK(clknet_leaf_102_clk_i),
    .D(net668),
    .RESET_B(net247),
    .Q(\line_cache[231][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25322_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01171_),
    .RESET_B(net245),
    .Q(\line_cache[231][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25323_ (.CLK(clknet_leaf_123_clk_i),
    .D(net1549),
    .RESET_B(net323),
    .Q(\line_cache[231][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25324_ (.CLK(clknet_leaf_102_clk_i),
    .D(net1596),
    .RESET_B(net247),
    .Q(\line_cache[231][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25325_ (.CLK(clknet_leaf_113_clk_i),
    .D(net1218),
    .RESET_B(net237),
    .Q(\line_cache[231][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25326_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01175_),
    .RESET_B(net246),
    .Q(\line_cache[231][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25327_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01176_),
    .RESET_B(net245),
    .Q(\line_cache[232][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25328_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01177_),
    .RESET_B(net245),
    .Q(\line_cache[232][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25329_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01178_),
    .RESET_B(net245),
    .Q(\line_cache[232][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25330_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01179_),
    .RESET_B(net245),
    .Q(\line_cache[232][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25331_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01180_),
    .RESET_B(net247),
    .Q(\line_cache[232][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25332_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01181_),
    .RESET_B(net245),
    .Q(\line_cache[232][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25333_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01182_),
    .RESET_B(net237),
    .Q(\line_cache[232][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25334_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01183_),
    .RESET_B(net235),
    .Q(\line_cache[232][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25335_ (.CLK(clknet_leaf_112_clk_i),
    .D(net636),
    .RESET_B(net238),
    .Q(\line_cache[233][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25336_ (.CLK(clknet_leaf_115_clk_i),
    .D(net2072),
    .RESET_B(net237),
    .Q(\line_cache[233][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25337_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01186_),
    .RESET_B(net235),
    .Q(\line_cache[233][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25338_ (.CLK(clknet_leaf_113_clk_i),
    .D(net2442),
    .RESET_B(net237),
    .Q(\line_cache[233][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25339_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01188_),
    .RESET_B(net238),
    .Q(\line_cache[233][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25340_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01189_),
    .RESET_B(net235),
    .Q(\line_cache[233][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25341_ (.CLK(clknet_leaf_113_clk_i),
    .D(net2273),
    .RESET_B(net238),
    .Q(\line_cache[233][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25342_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01191_),
    .RESET_B(net247),
    .Q(\line_cache[233][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25343_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01192_),
    .RESET_B(net238),
    .Q(\line_cache[234][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25344_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01193_),
    .RESET_B(net238),
    .Q(\line_cache[234][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25345_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01194_),
    .RESET_B(net238),
    .Q(\line_cache[234][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25346_ (.CLK(clknet_leaf_113_clk_i),
    .D(net1692),
    .RESET_B(net238),
    .Q(\line_cache[234][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25347_ (.CLK(clknet_leaf_123_clk_i),
    .D(net1030),
    .RESET_B(net323),
    .Q(\line_cache[234][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25348_ (.CLK(clknet_leaf_112_clk_i),
    .D(net956),
    .RESET_B(net238),
    .Q(\line_cache[234][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25349_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01198_),
    .RESET_B(net238),
    .Q(\line_cache[234][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25350_ (.CLK(clknet_leaf_111_clk_i),
    .D(net2126),
    .RESET_B(net238),
    .Q(\line_cache[234][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25351_ (.CLK(clknet_leaf_114_clk_i),
    .D(net910),
    .RESET_B(net237),
    .Q(\line_cache[235][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25352_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01201_),
    .RESET_B(net237),
    .Q(\line_cache[235][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25353_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01202_),
    .RESET_B(net237),
    .Q(\line_cache[235][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25354_ (.CLK(clknet_leaf_113_clk_i),
    .D(net2579),
    .RESET_B(net237),
    .Q(\line_cache[235][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25355_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01204_),
    .RESET_B(net237),
    .Q(\line_cache[235][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25356_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01205_),
    .RESET_B(net237),
    .Q(\line_cache[235][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25357_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01206_),
    .RESET_B(net237),
    .Q(\line_cache[235][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25358_ (.CLK(clknet_leaf_113_clk_i),
    .D(net2457),
    .RESET_B(net323),
    .Q(\line_cache[235][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25359_ (.CLK(clknet_leaf_116_clk_i),
    .D(net2155),
    .RESET_B(net233),
    .Q(\line_cache[236][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25360_ (.CLK(clknet_leaf_122_clk_i),
    .D(net1629),
    .RESET_B(net320),
    .Q(\line_cache[236][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25361_ (.CLK(clknet_leaf_114_clk_i),
    .D(net1414),
    .RESET_B(net237),
    .Q(\line_cache[236][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25362_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01211_),
    .RESET_B(net321),
    .Q(\line_cache[236][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25363_ (.CLK(clknet_leaf_116_clk_i),
    .D(net2374),
    .RESET_B(net233),
    .Q(\line_cache[236][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25364_ (.CLK(clknet_leaf_113_clk_i),
    .D(net1820),
    .RESET_B(net237),
    .Q(\line_cache[236][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25365_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01214_),
    .RESET_B(net320),
    .Q(\line_cache[236][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25366_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01215_),
    .RESET_B(net320),
    .Q(\line_cache[236][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25367_ (.CLK(clknet_leaf_114_clk_i),
    .D(net1504),
    .RESET_B(net320),
    .Q(\line_cache[237][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25368_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01217_),
    .RESET_B(net321),
    .Q(\line_cache[237][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25369_ (.CLK(clknet_leaf_122_clk_i),
    .D(net1718),
    .RESET_B(net320),
    .Q(\line_cache[237][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25370_ (.CLK(clknet_leaf_122_clk_i),
    .D(net1976),
    .RESET_B(net320),
    .Q(\line_cache[237][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25371_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01220_),
    .RESET_B(net234),
    .Q(\line_cache[237][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25372_ (.CLK(clknet_leaf_121_clk_i),
    .D(net3751),
    .RESET_B(net321),
    .Q(\line_cache[237][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25373_ (.CLK(clknet_leaf_123_clk_i),
    .D(net2225),
    .RESET_B(net323),
    .Q(\line_cache[237][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25374_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01223_),
    .RESET_B(net321),
    .Q(\line_cache[237][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25375_ (.CLK(clknet_leaf_117_clk_i),
    .D(net1312),
    .RESET_B(net316),
    .Q(\line_cache[238][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25376_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01225_),
    .RESET_B(net321),
    .Q(\line_cache[238][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25377_ (.CLK(clknet_leaf_122_clk_i),
    .D(net3722),
    .RESET_B(net320),
    .Q(\line_cache[238][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25378_ (.CLK(clknet_leaf_122_clk_i),
    .D(net1580),
    .RESET_B(net320),
    .Q(\line_cache[238][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25379_ (.CLK(clknet_leaf_120_clk_i),
    .D(net2107),
    .RESET_B(net316),
    .Q(\line_cache[238][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25380_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01229_),
    .RESET_B(net320),
    .Q(\line_cache[238][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25381_ (.CLK(clknet_leaf_122_clk_i),
    .D(net1452),
    .RESET_B(net320),
    .Q(\line_cache[238][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25382_ (.CLK(clknet_leaf_125_clk_i),
    .D(net1014),
    .RESET_B(net320),
    .Q(\line_cache[238][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25383_ (.CLK(clknet_leaf_117_clk_i),
    .D(net3657),
    .RESET_B(net234),
    .Q(\line_cache[239][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25384_ (.CLK(clknet_leaf_121_clk_i),
    .D(net3619),
    .RESET_B(net318),
    .Q(\line_cache[239][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25385_ (.CLK(clknet_leaf_120_clk_i),
    .D(net570),
    .RESET_B(net316),
    .Q(\line_cache[239][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25386_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01235_),
    .RESET_B(net318),
    .Q(\line_cache[239][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25387_ (.CLK(clknet_leaf_117_clk_i),
    .D(net544),
    .RESET_B(net316),
    .Q(\line_cache[239][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25388_ (.CLK(clknet_leaf_117_clk_i),
    .D(net3215),
    .RESET_B(net234),
    .Q(\line_cache[239][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25389_ (.CLK(clknet_leaf_120_clk_i),
    .D(net538),
    .RESET_B(net316),
    .Q(\line_cache[239][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25390_ (.CLK(clknet_leaf_120_clk_i),
    .D(net988),
    .RESET_B(net316),
    .Q(\line_cache[239][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25391_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01248_),
    .RESET_B(net319),
    .Q(\line_cache[240][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25392_ (.CLK(clknet_leaf_120_clk_i),
    .D(net1946),
    .RESET_B(net318),
    .Q(\line_cache[240][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25393_ (.CLK(clknet_leaf_120_clk_i),
    .D(net1524),
    .RESET_B(net319),
    .Q(\line_cache[240][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25394_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01251_),
    .RESET_B(net318),
    .Q(\line_cache[240][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25395_ (.CLK(clknet_leaf_119_clk_i),
    .D(net660),
    .RESET_B(net316),
    .Q(\line_cache[240][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25396_ (.CLK(clknet_leaf_119_clk_i),
    .D(net838),
    .RESET_B(net316),
    .Q(\line_cache[240][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25397_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01254_),
    .RESET_B(net316),
    .Q(\line_cache[240][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25398_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01255_),
    .RESET_B(net317),
    .Q(\line_cache[240][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25399_ (.CLK(clknet_leaf_117_clk_i),
    .D(net524),
    .RESET_B(net234),
    .Q(\line_cache[241][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25400_ (.CLK(clknet_leaf_120_clk_i),
    .D(net542),
    .RESET_B(net319),
    .Q(\line_cache[241][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25401_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01258_),
    .RESET_B(net318),
    .Q(\line_cache[241][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25402_ (.CLK(clknet_leaf_120_clk_i),
    .D(net592),
    .RESET_B(net318),
    .Q(\line_cache[241][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25403_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01260_),
    .RESET_B(net317),
    .Q(\line_cache[241][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25404_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01261_),
    .RESET_B(net317),
    .Q(\line_cache[241][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25405_ (.CLK(clknet_leaf_120_clk_i),
    .D(net480),
    .RESET_B(net319),
    .Q(\line_cache[241][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25406_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01263_),
    .RESET_B(net317),
    .Q(\line_cache[241][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25407_ (.CLK(clknet_leaf_118_clk_i),
    .D(net550),
    .RESET_B(net316),
    .Q(\line_cache[242][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25408_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01265_),
    .RESET_B(net318),
    .Q(\line_cache[242][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25409_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01266_),
    .RESET_B(net319),
    .Q(\line_cache[242][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25410_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01267_),
    .RESET_B(net318),
    .Q(\line_cache[242][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25411_ (.CLK(clknet_leaf_118_clk_i),
    .D(net454),
    .RESET_B(net233),
    .Q(\line_cache[242][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25412_ (.CLK(clknet_leaf_118_clk_i),
    .D(net536),
    .RESET_B(net233),
    .Q(\line_cache[242][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25413_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01270_),
    .RESET_B(net316),
    .Q(\line_cache[242][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25414_ (.CLK(clknet_leaf_193_clk_i),
    .D(net448),
    .RESET_B(net317),
    .Q(\line_cache[242][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25415_ (.CLK(clknet_leaf_191_clk_i),
    .D(_01272_),
    .RESET_B(net317),
    .Q(\line_cache[243][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25416_ (.CLK(clknet_leaf_192_clk_i),
    .D(net470),
    .RESET_B(net317),
    .Q(\line_cache[243][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25417_ (.CLK(clknet_leaf_119_clk_i),
    .D(net418),
    .RESET_B(net316),
    .Q(\line_cache[243][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25418_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01275_),
    .RESET_B(net317),
    .Q(\line_cache[243][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25419_ (.CLK(clknet_leaf_119_clk_i),
    .D(net502),
    .RESET_B(net316),
    .Q(\line_cache[243][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25420_ (.CLK(clknet_leaf_192_clk_i),
    .D(net428),
    .RESET_B(net317),
    .Q(\line_cache[243][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25421_ (.CLK(clknet_leaf_193_clk_i),
    .D(net458),
    .RESET_B(net316),
    .Q(\line_cache[243][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25422_ (.CLK(clknet_leaf_193_clk_i),
    .D(net528),
    .RESET_B(net316),
    .Q(\line_cache[243][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25423_ (.CLK(clknet_leaf_194_clk_i),
    .D(net706),
    .RESET_B(net274),
    .Q(\line_cache[244][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25424_ (.CLK(clknet_leaf_199_clk_i),
    .D(_01281_),
    .RESET_B(net274),
    .Q(\line_cache[244][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25425_ (.CLK(clknet_leaf_193_clk_i),
    .D(net1052),
    .RESET_B(net273),
    .Q(\line_cache[244][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25426_ (.CLK(clknet_leaf_199_clk_i),
    .D(_01283_),
    .RESET_B(net283),
    .Q(\line_cache[244][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25427_ (.CLK(clknet_leaf_193_clk_i),
    .D(net734),
    .RESET_B(net316),
    .Q(\line_cache[244][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25428_ (.CLK(clknet_leaf_192_clk_i),
    .D(net682),
    .RESET_B(net317),
    .Q(\line_cache[244][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25429_ (.CLK(clknet_leaf_192_clk_i),
    .D(_01286_),
    .RESET_B(net317),
    .Q(\line_cache[244][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25430_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01287_),
    .RESET_B(net274),
    .Q(\line_cache[244][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25431_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01288_),
    .RESET_B(net274),
    .Q(\line_cache[245][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25432_ (.CLK(clknet_leaf_194_clk_i),
    .D(_01289_),
    .RESET_B(net274),
    .Q(\line_cache[245][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25433_ (.CLK(clknet_leaf_194_clk_i),
    .D(net1114),
    .RESET_B(net273),
    .Q(\line_cache[245][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25434_ (.CLK(clknet_leaf_194_clk_i),
    .D(net826),
    .RESET_B(net275),
    .Q(\line_cache[245][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25435_ (.CLK(clknet_leaf_39_clk_i),
    .D(net1146),
    .RESET_B(net273),
    .Q(\line_cache[245][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25436_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01293_),
    .RESET_B(net275),
    .Q(\line_cache[245][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25437_ (.CLK(clknet_leaf_193_clk_i),
    .D(net1354),
    .RESET_B(net273),
    .Q(\line_cache[245][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25438_ (.CLK(clknet_leaf_198_clk_i),
    .D(_01295_),
    .RESET_B(net283),
    .Q(\line_cache[245][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25439_ (.CLK(clknet_leaf_195_clk_i),
    .D(net936),
    .RESET_B(net275),
    .Q(\line_cache[246][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25440_ (.CLK(clknet_leaf_195_clk_i),
    .D(_01297_),
    .RESET_B(net275),
    .Q(\line_cache[246][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25441_ (.CLK(clknet_leaf_198_clk_i),
    .D(_01298_),
    .RESET_B(net283),
    .Q(\line_cache[246][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25442_ (.CLK(clknet_leaf_198_clk_i),
    .D(_01299_),
    .RESET_B(net283),
    .Q(\line_cache[246][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25443_ (.CLK(clknet_leaf_285_clk_i),
    .D(net1240),
    .RESET_B(net275),
    .Q(\line_cache[246][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25444_ (.CLK(clknet_leaf_193_clk_i),
    .D(net1012),
    .RESET_B(net275),
    .Q(\line_cache[246][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25445_ (.CLK(clknet_leaf_193_clk_i),
    .D(net1196),
    .RESET_B(net275),
    .Q(\line_cache[246][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25446_ (.CLK(clknet_leaf_194_clk_i),
    .D(net886),
    .RESET_B(net275),
    .Q(\line_cache[246][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25447_ (.CLK(clknet_leaf_196_clk_i),
    .D(net1402),
    .RESET_B(net274),
    .Q(\line_cache[247][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25448_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1450),
    .RESET_B(net273),
    .Q(\line_cache[247][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25449_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1927),
    .RESET_B(net273),
    .Q(\line_cache[247][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25450_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1701),
    .RESET_B(net273),
    .Q(\line_cache[247][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25451_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01308_),
    .RESET_B(net273),
    .Q(\line_cache[247][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25452_ (.CLK(clknet_leaf_196_clk_i),
    .D(_01309_),
    .RESET_B(net274),
    .Q(\line_cache[247][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25453_ (.CLK(clknet_leaf_196_clk_i),
    .D(net798),
    .RESET_B(net274),
    .Q(\line_cache[247][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25454_ (.CLK(clknet_leaf_196_clk_i),
    .D(_01311_),
    .RESET_B(net274),
    .Q(\line_cache[247][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25455_ (.CLK(clknet_leaf_283_clk_i),
    .D(_01312_),
    .RESET_B(net271),
    .Q(\line_cache[248][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25456_ (.CLK(clknet_leaf_284_clk_i),
    .D(net2102),
    .RESET_B(net273),
    .Q(\line_cache[248][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25457_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01314_),
    .RESET_B(net273),
    .Q(\line_cache[248][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25458_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01315_),
    .RESET_B(net273),
    .Q(\line_cache[248][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25459_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01316_),
    .RESET_B(net273),
    .Q(\line_cache[248][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25460_ (.CLK(clknet_leaf_283_clk_i),
    .D(_01317_),
    .RESET_B(net274),
    .Q(\line_cache[248][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25461_ (.CLK(clknet_leaf_196_clk_i),
    .D(_01318_),
    .RESET_B(net274),
    .Q(\line_cache[248][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25462_ (.CLK(clknet_leaf_283_clk_i),
    .D(_01319_),
    .RESET_B(net274),
    .Q(\line_cache[248][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25463_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01320_),
    .RESET_B(net200),
    .Q(\line_cache[249][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25464_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1699),
    .RESET_B(net273),
    .Q(\line_cache[249][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25465_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1899),
    .RESET_B(net273),
    .Q(\line_cache[249][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25466_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1662),
    .RESET_B(net275),
    .Q(\line_cache[249][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25467_ (.CLK(clknet_leaf_287_clk_i),
    .D(net1056),
    .RESET_B(net273),
    .Q(\line_cache[249][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25468_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01325_),
    .RESET_B(net271),
    .Q(\line_cache[249][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25469_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1442),
    .RESET_B(net275),
    .Q(\line_cache[249][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25470_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01327_),
    .RESET_B(net271),
    .Q(\line_cache[249][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25471_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01336_),
    .RESET_B(net200),
    .Q(\line_cache[250][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25472_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01337_),
    .RESET_B(net271),
    .Q(\line_cache[250][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25473_ (.CLK(clknet_leaf_282_clk_i),
    .D(_01338_),
    .RESET_B(net272),
    .Q(\line_cache[250][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25474_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01339_),
    .RESET_B(net275),
    .Q(\line_cache[250][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25475_ (.CLK(clknet_leaf_287_clk_i),
    .D(net1867),
    .RESET_B(net200),
    .Q(\line_cache[250][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25476_ (.CLK(clknet_leaf_283_clk_i),
    .D(net2023),
    .RESET_B(net274),
    .Q(\line_cache[250][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25477_ (.CLK(clknet_leaf_284_clk_i),
    .D(_01342_),
    .RESET_B(net273),
    .Q(\line_cache[250][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25478_ (.CLK(clknet_leaf_284_clk_i),
    .D(net1528),
    .RESET_B(net274),
    .Q(\line_cache[250][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25479_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01344_),
    .RESET_B(net200),
    .Q(\line_cache[251][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25480_ (.CLK(clknet_leaf_285_clk_i),
    .D(net1376),
    .RESET_B(net200),
    .Q(\line_cache[251][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25481_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01346_),
    .RESET_B(net200),
    .Q(\line_cache[251][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25482_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01347_),
    .RESET_B(net200),
    .Q(\line_cache[251][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25483_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01348_),
    .RESET_B(net201),
    .Q(\line_cache[251][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25484_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01349_),
    .RESET_B(net200),
    .Q(\line_cache[251][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25485_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01350_),
    .RESET_B(net201),
    .Q(\line_cache[251][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25486_ (.CLK(clknet_leaf_38_clk_i),
    .D(net1799),
    .RESET_B(net201),
    .Q(\line_cache[251][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25487_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01352_),
    .RESET_B(net233),
    .Q(\line_cache[252][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25488_ (.CLK(clknet_leaf_39_clk_i),
    .D(net606),
    .RESET_B(net233),
    .Q(\line_cache[252][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25489_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01354_),
    .RESET_B(net200),
    .Q(\line_cache[252][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25490_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01355_),
    .RESET_B(net201),
    .Q(\line_cache[252][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25491_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01356_),
    .RESET_B(net234),
    .Q(\line_cache[252][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25492_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01357_),
    .RESET_B(net233),
    .Q(\line_cache[252][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25493_ (.CLK(clknet_leaf_40_clk_i),
    .D(net3958),
    .RESET_B(net231),
    .Q(\line_cache[252][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25494_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01359_),
    .RESET_B(net201),
    .Q(\line_cache[252][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25495_ (.CLK(clknet_leaf_40_clk_i),
    .D(net1226),
    .RESET_B(net233),
    .Q(\line_cache[253][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25496_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01361_),
    .RESET_B(net233),
    .Q(\line_cache[253][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25497_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01362_),
    .RESET_B(net200),
    .Q(\line_cache[253][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25498_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01363_),
    .RESET_B(net201),
    .Q(\line_cache[253][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25499_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01364_),
    .RESET_B(net231),
    .Q(\line_cache[253][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25500_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01365_),
    .RESET_B(net233),
    .Q(\line_cache[253][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25501_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01366_),
    .RESET_B(net233),
    .Q(\line_cache[253][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25502_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01367_),
    .RESET_B(net201),
    .Q(\line_cache[253][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25503_ (.CLK(clknet_leaf_40_clk_i),
    .D(net666),
    .RESET_B(net233),
    .Q(\line_cache[254][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25504_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01369_),
    .RESET_B(net233),
    .Q(\line_cache[254][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25505_ (.CLK(clknet_leaf_285_clk_i),
    .D(_01370_),
    .RESET_B(net201),
    .Q(\line_cache[254][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25506_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01371_),
    .RESET_B(net201),
    .Q(\line_cache[254][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25507_ (.CLK(clknet_leaf_39_clk_i),
    .D(net1756),
    .RESET_B(net233),
    .Q(\line_cache[254][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25508_ (.CLK(clknet_leaf_39_clk_i),
    .D(net1024),
    .RESET_B(net233),
    .Q(\line_cache[254][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25509_ (.CLK(clknet_leaf_39_clk_i),
    .D(net2135),
    .RESET_B(net233),
    .Q(\line_cache[254][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25510_ (.CLK(clknet_leaf_38_clk_i),
    .D(net1994),
    .RESET_B(net201),
    .Q(\line_cache[254][7] ));
 sky130_fd_sc_hd__dfrtp_2 _25511_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01376_),
    .RESET_B(net231),
    .Q(\line_cache[255][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25512_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01377_),
    .RESET_B(net231),
    .Q(\line_cache[255][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25513_ (.CLK(clknet_leaf_43_clk_i),
    .D(_01378_),
    .RESET_B(net225),
    .Q(\line_cache[255][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25514_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01379_),
    .RESET_B(net231),
    .Q(\line_cache[255][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25515_ (.CLK(clknet_leaf_41_clk_i),
    .D(_01380_),
    .RESET_B(net231),
    .Q(\line_cache[255][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25516_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01381_),
    .RESET_B(net231),
    .Q(\line_cache[255][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25517_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01382_),
    .RESET_B(net225),
    .Q(\line_cache[255][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25518_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01383_),
    .RESET_B(net231),
    .Q(\line_cache[255][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25519_ (.CLK(clknet_leaf_43_clk_i),
    .D(net1712),
    .RESET_B(net225),
    .Q(\line_cache[256][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25520_ (.CLK(clknet_leaf_41_clk_i),
    .D(_01385_),
    .RESET_B(net231),
    .Q(\line_cache[256][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25521_ (.CLK(clknet_leaf_41_clk_i),
    .D(net2421),
    .RESET_B(net225),
    .Q(\line_cache[256][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25522_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01387_),
    .RESET_B(net234),
    .Q(\line_cache[256][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25523_ (.CLK(clknet_leaf_42_clk_i),
    .D(net1654),
    .RESET_B(net225),
    .Q(\line_cache[256][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25524_ (.CLK(clknet_leaf_41_clk_i),
    .D(net3855),
    .RESET_B(net231),
    .Q(\line_cache[256][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25525_ (.CLK(clknet_leaf_41_clk_i),
    .D(net4120),
    .RESET_B(net232),
    .Q(\line_cache[256][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25526_ (.CLK(clknet_leaf_41_clk_i),
    .D(net4113),
    .RESET_B(net232),
    .Q(\line_cache[256][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25527_ (.CLK(clknet_leaf_41_clk_i),
    .D(net1954),
    .RESET_B(net231),
    .Q(\line_cache[257][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25528_ (.CLK(clknet_leaf_115_clk_i),
    .D(net1268),
    .RESET_B(net232),
    .Q(\line_cache[257][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25529_ (.CLK(clknet_leaf_116_clk_i),
    .D(net1831),
    .RESET_B(net232),
    .Q(\line_cache[257][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25530_ (.CLK(clknet_leaf_47_clk_i),
    .D(net2391),
    .RESET_B(net232),
    .Q(\line_cache[257][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25531_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01396_),
    .RESET_B(net237),
    .Q(\line_cache[257][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25532_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01397_),
    .RESET_B(net235),
    .Q(\line_cache[257][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25533_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01398_),
    .RESET_B(net237),
    .Q(\line_cache[257][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25534_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01399_),
    .RESET_B(net234),
    .Q(\line_cache[257][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25535_ (.CLK(clknet_leaf_41_clk_i),
    .D(net514),
    .RESET_B(net231),
    .Q(\line_cache[258][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25536_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01401_),
    .RESET_B(net232),
    .Q(\line_cache[258][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25537_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01402_),
    .RESET_B(net234),
    .Q(\line_cache[258][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25538_ (.CLK(clknet_leaf_42_clk_i),
    .D(net442),
    .RESET_B(net232),
    .Q(\line_cache[258][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25539_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01404_),
    .RESET_B(net234),
    .Q(\line_cache[258][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25540_ (.CLK(clknet_leaf_40_clk_i),
    .D(net916),
    .RESET_B(net231),
    .Q(\line_cache[258][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25541_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01406_),
    .RESET_B(net234),
    .Q(\line_cache[258][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25542_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01407_),
    .RESET_B(net234),
    .Q(\line_cache[258][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25543_ (.CLK(clknet_leaf_42_clk_i),
    .D(net902),
    .RESET_B(net225),
    .Q(\line_cache[259][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25544_ (.CLK(clknet_leaf_41_clk_i),
    .D(net812),
    .RESET_B(net232),
    .Q(\line_cache[259][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25545_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01410_),
    .RESET_B(net234),
    .Q(\line_cache[259][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25546_ (.CLK(clknet_leaf_47_clk_i),
    .D(net772),
    .RESET_B(net229),
    .Q(\line_cache[259][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25547_ (.CLK(clknet_leaf_115_clk_i),
    .D(net816),
    .RESET_B(net235),
    .Q(\line_cache[259][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25548_ (.CLK(clknet_leaf_110_clk_i),
    .D(net692),
    .RESET_B(net235),
    .Q(\line_cache[259][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25549_ (.CLK(clknet_leaf_41_clk_i),
    .D(net526),
    .RESET_B(net232),
    .Q(\line_cache[259][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25550_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01415_),
    .RESET_B(net234),
    .Q(\line_cache[259][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25551_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01424_),
    .RESET_B(net235),
    .Q(\line_cache[260][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25552_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01425_),
    .RESET_B(net235),
    .Q(\line_cache[260][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25553_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01426_),
    .RESET_B(net235),
    .Q(\line_cache[260][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25554_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01427_),
    .RESET_B(net237),
    .Q(\line_cache[260][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25555_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01428_),
    .RESET_B(net235),
    .Q(\line_cache[260][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25556_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01429_),
    .RESET_B(net235),
    .Q(\line_cache[260][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25557_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01430_),
    .RESET_B(net235),
    .Q(\line_cache[260][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25558_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01431_),
    .RESET_B(net235),
    .Q(\line_cache[260][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25559_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01432_),
    .RESET_B(net235),
    .Q(\line_cache[261][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25560_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01433_),
    .RESET_B(net229),
    .Q(\line_cache[261][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25561_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01434_),
    .RESET_B(net235),
    .Q(\line_cache[261][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25562_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01435_),
    .RESET_B(net245),
    .Q(\line_cache[261][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25563_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01436_),
    .RESET_B(net245),
    .Q(\line_cache[261][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25564_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01437_),
    .RESET_B(net236),
    .Q(\line_cache[261][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25565_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01438_),
    .RESET_B(net236),
    .Q(\line_cache[261][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25566_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01439_),
    .RESET_B(net236),
    .Q(\line_cache[261][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25567_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01440_),
    .RESET_B(net236),
    .Q(\line_cache[262][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25568_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01441_),
    .RESET_B(net245),
    .Q(\line_cache[262][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25569_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01442_),
    .RESET_B(net236),
    .Q(\line_cache[262][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25570_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01443_),
    .RESET_B(net245),
    .Q(\line_cache[262][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25571_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01444_),
    .RESET_B(net245),
    .Q(\line_cache[262][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25572_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01445_),
    .RESET_B(net236),
    .Q(\line_cache[262][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25573_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01446_),
    .RESET_B(net236),
    .Q(\line_cache[262][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25574_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01447_),
    .RESET_B(net236),
    .Q(\line_cache[262][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25575_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01448_),
    .RESET_B(net235),
    .Q(\line_cache[263][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25576_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01449_),
    .RESET_B(net241),
    .Q(\line_cache[263][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25577_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01450_),
    .RESET_B(net229),
    .Q(\line_cache[263][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25578_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01451_),
    .RESET_B(net241),
    .Q(\line_cache[263][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25579_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01452_),
    .RESET_B(net241),
    .Q(\line_cache[263][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25580_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01453_),
    .RESET_B(net229),
    .Q(\line_cache[263][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25581_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01454_),
    .RESET_B(net229),
    .Q(\line_cache[263][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25582_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01455_),
    .RESET_B(net229),
    .Q(\line_cache[263][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25583_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01456_),
    .RESET_B(net229),
    .Q(\line_cache[264][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25584_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01457_),
    .RESET_B(net241),
    .Q(\line_cache[264][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25585_ (.CLK(clknet_leaf_109_clk_i),
    .D(net1288),
    .RESET_B(net229),
    .Q(\line_cache[264][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25586_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01459_),
    .RESET_B(net229),
    .Q(\line_cache[264][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25587_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01460_),
    .RESET_B(net241),
    .Q(\line_cache[264][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25588_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01461_),
    .RESET_B(net229),
    .Q(\line_cache[264][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25589_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01462_),
    .RESET_B(net229),
    .Q(\line_cache[264][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25590_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01463_),
    .RESET_B(net230),
    .Q(\line_cache[264][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25591_ (.CLK(clknet_leaf_109_clk_i),
    .D(net912),
    .RESET_B(net229),
    .Q(\line_cache[265][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25592_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01465_),
    .RESET_B(net227),
    .Q(\line_cache[265][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25593_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01466_),
    .RESET_B(net228),
    .Q(\line_cache[265][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25594_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01467_),
    .RESET_B(net227),
    .Q(\line_cache[265][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25595_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01468_),
    .RESET_B(net228),
    .Q(\line_cache[265][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25596_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01469_),
    .RESET_B(net241),
    .Q(\line_cache[265][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25597_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01470_),
    .RESET_B(net228),
    .Q(\line_cache[265][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25598_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01471_),
    .RESET_B(net230),
    .Q(\line_cache[265][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25599_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01472_),
    .RESET_B(net230),
    .Q(\line_cache[266][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25600_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01473_),
    .RESET_B(net228),
    .Q(\line_cache[266][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25601_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01474_),
    .RESET_B(net240),
    .Q(\line_cache[266][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25602_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01475_),
    .RESET_B(net227),
    .Q(\line_cache[266][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25603_ (.CLK(clknet_leaf_49_clk_i),
    .D(net1418),
    .RESET_B(net227),
    .Q(\line_cache[266][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25604_ (.CLK(clknet_leaf_107_clk_i),
    .D(net1130),
    .RESET_B(net230),
    .Q(\line_cache[266][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25605_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01478_),
    .RESET_B(net228),
    .Q(\line_cache[266][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25606_ (.CLK(clknet_leaf_107_clk_i),
    .D(net1332),
    .RESET_B(net230),
    .Q(\line_cache[266][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25607_ (.CLK(clknet_leaf_48_clk_i),
    .D(net510),
    .RESET_B(net227),
    .Q(\line_cache[267][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25608_ (.CLK(clknet_leaf_49_clk_i),
    .D(net932),
    .RESET_B(net228),
    .Q(\line_cache[267][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25609_ (.CLK(clknet_leaf_49_clk_i),
    .D(net644),
    .RESET_B(net227),
    .Q(\line_cache[267][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25610_ (.CLK(clknet_leaf_51_clk_i),
    .D(net584),
    .RESET_B(net227),
    .Q(\line_cache[267][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25611_ (.CLK(clknet_leaf_48_clk_i),
    .D(net1180),
    .RESET_B(net227),
    .Q(\line_cache[267][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25612_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01485_),
    .RESET_B(net228),
    .Q(\line_cache[267][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25613_ (.CLK(clknet_leaf_49_clk_i),
    .D(net558),
    .RESET_B(net227),
    .Q(\line_cache[267][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25614_ (.CLK(clknet_leaf_48_clk_i),
    .D(net1448),
    .RESET_B(net227),
    .Q(\line_cache[267][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25615_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01488_),
    .RESET_B(net212),
    .Q(\line_cache[268][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25616_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01489_),
    .RESET_B(net212),
    .Q(\line_cache[268][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25617_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01490_),
    .RESET_B(net227),
    .Q(\line_cache[268][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25618_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01491_),
    .RESET_B(net228),
    .Q(\line_cache[268][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25619_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01492_),
    .RESET_B(net227),
    .Q(\line_cache[268][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25620_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01493_),
    .RESET_B(net228),
    .Q(\line_cache[268][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25621_ (.CLK(clknet_leaf_107_clk_i),
    .D(net4009),
    .RESET_B(net228),
    .Q(\line_cache[268][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25622_ (.CLK(clknet_leaf_48_clk_i),
    .D(net1608),
    .RESET_B(net227),
    .Q(\line_cache[268][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25623_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01496_),
    .RESET_B(net212),
    .Q(\line_cache[269][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25624_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01497_),
    .RESET_B(net212),
    .Q(\line_cache[269][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25625_ (.CLK(clknet_leaf_88_clk_i),
    .D(net2004),
    .RESET_B(net220),
    .Q(\line_cache[269][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25626_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01499_),
    .RESET_B(net220),
    .Q(\line_cache[269][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25627_ (.CLK(clknet_leaf_88_clk_i),
    .D(net1350),
    .RESET_B(net240),
    .Q(\line_cache[269][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25628_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01501_),
    .RESET_B(net240),
    .Q(\line_cache[269][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25629_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01502_),
    .RESET_B(net220),
    .Q(\line_cache[269][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25630_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01503_),
    .RESET_B(net240),
    .Q(\line_cache[269][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25631_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01512_),
    .RESET_B(net220),
    .Q(\line_cache[270][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25632_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01513_),
    .RESET_B(net240),
    .Q(\line_cache[270][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25633_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01514_),
    .RESET_B(net240),
    .Q(\line_cache[270][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25634_ (.CLK(clknet_leaf_87_clk_i),
    .D(net1736),
    .RESET_B(net220),
    .Q(\line_cache[270][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25635_ (.CLK(clknet_leaf_88_clk_i),
    .D(net1154),
    .RESET_B(net240),
    .Q(\line_cache[270][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25636_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01517_),
    .RESET_B(net240),
    .Q(\line_cache[270][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25637_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01518_),
    .RESET_B(net212),
    .Q(\line_cache[270][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25638_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01519_),
    .RESET_B(net240),
    .Q(\line_cache[270][7] ));
 sky130_fd_sc_hd__dfrtp_4 _25639_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01520_),
    .RESET_B(net240),
    .Q(\line_cache[271][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25640_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01521_),
    .RESET_B(net224),
    .Q(\line_cache[271][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25641_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01522_),
    .RESET_B(net227),
    .Q(\line_cache[271][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25642_ (.CLK(clknet_leaf_46_clk_i),
    .D(_01523_),
    .RESET_B(net224),
    .Q(\line_cache[271][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25643_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01524_),
    .RESET_B(net224),
    .Q(\line_cache[271][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25644_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01525_),
    .RESET_B(net227),
    .Q(\line_cache[271][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25645_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01526_),
    .RESET_B(net240),
    .Q(\line_cache[271][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25646_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01527_),
    .RESET_B(net240),
    .Q(\line_cache[271][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25647_ (.CLK(clknet_leaf_87_clk_i),
    .D(net2614),
    .RESET_B(net220),
    .Q(\line_cache[272][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25648_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01529_),
    .RESET_B(net222),
    .Q(\line_cache[272][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25649_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01530_),
    .RESET_B(net222),
    .Q(\line_cache[272][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25650_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01531_),
    .RESET_B(net218),
    .Q(\line_cache[272][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25651_ (.CLK(clknet_leaf_86_clk_i),
    .D(net2625),
    .RESET_B(net220),
    .Q(\line_cache[272][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25652_ (.CLK(clknet_leaf_87_clk_i),
    .D(net1987),
    .RESET_B(net220),
    .Q(\line_cache[272][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25653_ (.CLK(clknet_leaf_86_clk_i),
    .D(net3821),
    .RESET_B(net220),
    .Q(\line_cache[272][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25654_ (.CLK(clknet_leaf_86_clk_i),
    .D(net3679),
    .RESET_B(net221),
    .Q(\line_cache[272][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25655_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01536_),
    .RESET_B(net218),
    .Q(\line_cache[273][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25656_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01537_),
    .RESET_B(net222),
    .Q(\line_cache[273][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25657_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01538_),
    .RESET_B(net219),
    .Q(\line_cache[273][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25658_ (.CLK(clknet_leaf_85_clk_i),
    .D(net2581),
    .RESET_B(net219),
    .Q(\line_cache[273][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25659_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01540_),
    .RESET_B(net221),
    .Q(\line_cache[273][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25660_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01541_),
    .RESET_B(net221),
    .Q(\line_cache[273][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25661_ (.CLK(clknet_leaf_71_clk_i),
    .D(net2637),
    .RESET_B(net218),
    .Q(\line_cache[273][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25662_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01543_),
    .RESET_B(net221),
    .Q(\line_cache[273][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25663_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01544_),
    .RESET_B(net219),
    .Q(\line_cache[274][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25664_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01545_),
    .RESET_B(net219),
    .Q(\line_cache[274][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25665_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01546_),
    .RESET_B(net222),
    .Q(\line_cache[274][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25666_ (.CLK(clknet_leaf_85_clk_i),
    .D(net1933),
    .RESET_B(net219),
    .Q(\line_cache[274][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25667_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01548_),
    .RESET_B(net222),
    .Q(\line_cache[274][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25668_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01549_),
    .RESET_B(net219),
    .Q(\line_cache[274][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25669_ (.CLK(clknet_leaf_72_clk_i),
    .D(net1911),
    .RESET_B(net219),
    .Q(\line_cache[274][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25670_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01551_),
    .RESET_B(net219),
    .Q(\line_cache[274][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25671_ (.CLK(clknet_leaf_86_clk_i),
    .D(net860),
    .RESET_B(net221),
    .Q(\line_cache[275][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25672_ (.CLK(clknet_leaf_85_clk_i),
    .D(net1627),
    .RESET_B(net219),
    .Q(\line_cache[275][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25673_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01554_),
    .RESET_B(net219),
    .Q(\line_cache[275][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25674_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01555_),
    .RESET_B(net222),
    .Q(\line_cache[275][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25675_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01556_),
    .RESET_B(net222),
    .Q(\line_cache[275][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25676_ (.CLK(clknet_leaf_72_clk_i),
    .D(net2018),
    .RESET_B(net219),
    .Q(\line_cache[275][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25677_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01558_),
    .RESET_B(net219),
    .Q(\line_cache[275][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25678_ (.CLK(clknet_5_11__leaf_clk_i),
    .D(_01559_),
    .RESET_B(net222),
    .Q(\line_cache[275][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25679_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01560_),
    .RESET_B(net222),
    .Q(\line_cache[276][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25680_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01561_),
    .RESET_B(net222),
    .Q(\line_cache[276][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25681_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01562_),
    .RESET_B(net222),
    .Q(\line_cache[276][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25682_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01563_),
    .RESET_B(net222),
    .Q(\line_cache[276][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25683_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01564_),
    .RESET_B(net222),
    .Q(\line_cache[276][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25684_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01565_),
    .RESET_B(net221),
    .Q(\line_cache[276][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25685_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01566_),
    .RESET_B(net240),
    .Q(\line_cache[276][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25686_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01567_),
    .RESET_B(net221),
    .Q(\line_cache[276][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25687_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01568_),
    .RESET_B(net243),
    .Q(\line_cache[277][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25688_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01569_),
    .RESET_B(net222),
    .Q(\line_cache[277][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25689_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01570_),
    .RESET_B(net222),
    .Q(\line_cache[277][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25690_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01571_),
    .RESET_B(net222),
    .Q(\line_cache[277][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25691_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01572_),
    .RESET_B(net223),
    .Q(\line_cache[277][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25692_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01573_),
    .RESET_B(net223),
    .Q(\line_cache[277][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25693_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01574_),
    .RESET_B(net243),
    .Q(\line_cache[277][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25694_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01575_),
    .RESET_B(net243),
    .Q(\line_cache[277][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25695_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01576_),
    .RESET_B(net243),
    .Q(\line_cache[278][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25696_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01577_),
    .RESET_B(net243),
    .Q(\line_cache[278][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25697_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01578_),
    .RESET_B(net243),
    .Q(\line_cache[278][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25698_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01579_),
    .RESET_B(net244),
    .Q(\line_cache[278][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25699_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01580_),
    .RESET_B(net244),
    .Q(\line_cache[278][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25700_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01581_),
    .RESET_B(net243),
    .Q(\line_cache[278][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25701_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01582_),
    .RESET_B(net243),
    .Q(\line_cache[278][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25702_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01583_),
    .RESET_B(net243),
    .Q(\line_cache[278][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25703_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01584_),
    .RESET_B(net240),
    .Q(\line_cache[279][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25704_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01585_),
    .RESET_B(net243),
    .Q(\line_cache[279][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25705_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01586_),
    .RESET_B(net243),
    .Q(\line_cache[279][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25706_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01587_),
    .RESET_B(net243),
    .Q(\line_cache[279][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25707_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01588_),
    .RESET_B(net244),
    .Q(\line_cache[279][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25708_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01589_),
    .RESET_B(net243),
    .Q(\line_cache[279][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25709_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01590_),
    .RESET_B(net243),
    .Q(\line_cache[279][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25710_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01591_),
    .RESET_B(net243),
    .Q(\line_cache[279][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25711_ (.CLK(clknet_leaf_89_clk_i),
    .D(net2196),
    .RESET_B(net240),
    .Q(\line_cache[280][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25712_ (.CLK(clknet_leaf_89_clk_i),
    .D(net1410),
    .RESET_B(net242),
    .Q(\line_cache[280][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25713_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01602_),
    .RESET_B(net243),
    .Q(\line_cache[280][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25714_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01603_),
    .RESET_B(net242),
    .Q(\line_cache[280][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25715_ (.CLK(clknet_leaf_90_clk_i),
    .D(net2598),
    .RESET_B(net241),
    .Q(\line_cache[280][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25716_ (.CLK(clknet_leaf_90_clk_i),
    .D(net3428),
    .RESET_B(net242),
    .Q(\line_cache[280][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25717_ (.CLK(clknet_leaf_89_clk_i),
    .D(net3717),
    .RESET_B(net242),
    .Q(\line_cache[280][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25718_ (.CLK(clknet_leaf_90_clk_i),
    .D(net874),
    .RESET_B(net241),
    .Q(\line_cache[280][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25719_ (.CLK(clknet_leaf_90_clk_i),
    .D(net710),
    .RESET_B(net241),
    .Q(\line_cache[281][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25720_ (.CLK(clknet_leaf_88_clk_i),
    .D(net2571),
    .RESET_B(net240),
    .Q(\line_cache[281][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25721_ (.CLK(clknet_leaf_89_clk_i),
    .D(net1476),
    .RESET_B(net242),
    .Q(\line_cache[281][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25722_ (.CLK(clknet_leaf_89_clk_i),
    .D(net2576),
    .RESET_B(net242),
    .Q(\line_cache[281][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25723_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01612_),
    .RESET_B(net244),
    .Q(\line_cache[281][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25724_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01613_),
    .RESET_B(net242),
    .Q(\line_cache[281][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25725_ (.CLK(clknet_leaf_89_clk_i),
    .D(net1816),
    .RESET_B(net242),
    .Q(\line_cache[281][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25726_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01615_),
    .RESET_B(net244),
    .Q(\line_cache[281][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25727_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01616_),
    .RESET_B(net244),
    .Q(\line_cache[282][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25728_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01617_),
    .RESET_B(net249),
    .Q(\line_cache[282][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25729_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01618_),
    .RESET_B(net244),
    .Q(\line_cache[282][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25730_ (.CLK(clknet_leaf_90_clk_i),
    .D(net1262),
    .RESET_B(net242),
    .Q(\line_cache[282][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25731_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01620_),
    .RESET_B(net244),
    .Q(\line_cache[282][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25732_ (.CLK(clknet_leaf_104_clk_i),
    .D(net878),
    .RESET_B(net242),
    .Q(\line_cache[282][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25733_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01622_),
    .RESET_B(net244),
    .Q(\line_cache[282][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25734_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01623_),
    .RESET_B(net244),
    .Q(\line_cache[282][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25735_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01624_),
    .RESET_B(net242),
    .Q(\line_cache[283][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25736_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01625_),
    .RESET_B(net249),
    .Q(\line_cache[283][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25737_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01626_),
    .RESET_B(net244),
    .Q(\line_cache[283][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25738_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01627_),
    .RESET_B(net244),
    .Q(\line_cache[283][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25739_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01628_),
    .RESET_B(net244),
    .Q(\line_cache[283][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25740_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01629_),
    .RESET_B(net249),
    .Q(\line_cache[283][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25741_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01630_),
    .RESET_B(net244),
    .Q(\line_cache[283][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25742_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01631_),
    .RESET_B(net249),
    .Q(\line_cache[283][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25743_ (.CLK(clknet_leaf_104_clk_i),
    .D(net2302),
    .RESET_B(net242),
    .Q(\line_cache[284][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25744_ (.CLK(clknet_leaf_99_clk_i),
    .D(net2120),
    .RESET_B(net246),
    .Q(\line_cache[284][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25745_ (.CLK(clknet_leaf_105_clk_i),
    .D(net2620),
    .RESET_B(net241),
    .Q(\line_cache[284][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25746_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01635_),
    .RESET_B(net246),
    .Q(\line_cache[284][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25747_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01636_),
    .RESET_B(net245),
    .Q(\line_cache[284][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25748_ (.CLK(clknet_leaf_104_clk_i),
    .D(net1619),
    .RESET_B(net246),
    .Q(\line_cache[284][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25749_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01638_),
    .RESET_B(net241),
    .Q(\line_cache[284][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25750_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01639_),
    .RESET_B(net246),
    .Q(\line_cache[284][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25751_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01640_),
    .RESET_B(net241),
    .Q(\line_cache[285][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25752_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01641_),
    .RESET_B(net249),
    .Q(\line_cache[285][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25753_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01642_),
    .RESET_B(net241),
    .Q(\line_cache[285][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25754_ (.CLK(clknet_leaf_104_clk_i),
    .D(net2172),
    .RESET_B(net242),
    .Q(\line_cache[285][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25755_ (.CLK(clknet_leaf_103_clk_i),
    .D(net2223),
    .RESET_B(net245),
    .Q(\line_cache[285][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25756_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01645_),
    .RESET_B(net246),
    .Q(\line_cache[285][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25757_ (.CLK(clknet_leaf_105_clk_i),
    .D(net1458),
    .RESET_B(net241),
    .Q(\line_cache[285][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25758_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01647_),
    .RESET_B(net246),
    .Q(\line_cache[285][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25759_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01648_),
    .RESET_B(net241),
    .Q(\line_cache[286][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25760_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01649_),
    .RESET_B(net249),
    .Q(\line_cache[286][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25761_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01650_),
    .RESET_B(net249),
    .Q(\line_cache[286][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25762_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01651_),
    .RESET_B(net246),
    .Q(\line_cache[286][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25763_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01652_),
    .RESET_B(net246),
    .Q(\line_cache[286][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25764_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01653_),
    .RESET_B(net246),
    .Q(\line_cache[286][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25765_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01654_),
    .RESET_B(net249),
    .Q(\line_cache[286][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25766_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01655_),
    .RESET_B(net249),
    .Q(\line_cache[286][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25767_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01656_),
    .RESET_B(net229),
    .Q(\line_cache[287][0] ));
 sky130_fd_sc_hd__dfrtp_4 _25768_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01657_),
    .RESET_B(net245),
    .Q(\line_cache[287][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25769_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01658_),
    .RESET_B(net229),
    .Q(\line_cache[287][2] ));
 sky130_fd_sc_hd__dfrtp_2 _25770_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01659_),
    .RESET_B(net229),
    .Q(\line_cache[287][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25771_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01660_),
    .RESET_B(net227),
    .Q(\line_cache[287][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25772_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01661_),
    .RESET_B(net229),
    .Q(\line_cache[287][5] ));
 sky130_fd_sc_hd__dfrtp_4 _25773_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01662_),
    .RESET_B(net241),
    .Q(\line_cache[287][6] ));
 sky130_fd_sc_hd__dfrtp_4 _25774_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01663_),
    .RESET_B(net245),
    .Q(\line_cache[287][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25775_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01664_),
    .RESET_B(net220),
    .Q(\line_cache[288][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25776_ (.CLK(clknet_leaf_71_clk_i),
    .D(net862),
    .RESET_B(net218),
    .Q(\line_cache[288][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25777_ (.CLK(clknet_leaf_74_clk_i),
    .D(net2475),
    .RESET_B(net218),
    .Q(\line_cache[288][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25778_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01667_),
    .RESET_B(net220),
    .Q(\line_cache[288][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25779_ (.CLK(clknet_leaf_69_clk_i),
    .D(net2295),
    .RESET_B(net220),
    .Q(\line_cache[288][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25780_ (.CLK(clknet_leaf_68_clk_i),
    .D(net1770),
    .RESET_B(net211),
    .Q(\line_cache[288][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25781_ (.CLK(clknet_leaf_68_clk_i),
    .D(net3550),
    .RESET_B(net211),
    .Q(\line_cache[288][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25782_ (.CLK(clknet_leaf_70_clk_i),
    .D(net3581),
    .RESET_B(net218),
    .Q(\line_cache[288][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25783_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01672_),
    .RESET_B(net220),
    .Q(\line_cache[289][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25784_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01673_),
    .RESET_B(net218),
    .Q(\line_cache[289][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25785_ (.CLK(clknet_leaf_74_clk_i),
    .D(net1795),
    .RESET_B(net218),
    .Q(\line_cache[289][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25786_ (.CLK(clknet_leaf_68_clk_i),
    .D(net1909),
    .RESET_B(net213),
    .Q(\line_cache[289][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25787_ (.CLK(clknet_leaf_69_clk_i),
    .D(net1474),
    .RESET_B(net220),
    .Q(\line_cache[289][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25788_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01677_),
    .RESET_B(net218),
    .Q(\line_cache[289][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25789_ (.CLK(clknet_leaf_68_clk_i),
    .D(net1508),
    .RESET_B(net211),
    .Q(\line_cache[289][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25790_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01679_),
    .RESET_B(net218),
    .Q(\line_cache[289][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25791_ (.CLK(clknet_leaf_69_clk_i),
    .D(net1484),
    .RESET_B(net213),
    .Q(\line_cache[290][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25792_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01689_),
    .RESET_B(net216),
    .Q(\line_cache[290][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25793_ (.CLK(clknet_leaf_74_clk_i),
    .D(_01690_),
    .RESET_B(net216),
    .Q(\line_cache[290][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25794_ (.CLK(clknet_leaf_69_clk_i),
    .D(net1212),
    .RESET_B(net213),
    .Q(\line_cache[290][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25795_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01692_),
    .RESET_B(net220),
    .Q(\line_cache[290][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25796_ (.CLK(clknet_leaf_67_clk_i),
    .D(net1004),
    .RESET_B(net211),
    .Q(\line_cache[290][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25797_ (.CLK(clknet_leaf_68_clk_i),
    .D(net1697),
    .RESET_B(net214),
    .Q(\line_cache[290][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25798_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01695_),
    .RESET_B(net218),
    .Q(\line_cache[290][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25799_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01696_),
    .RESET_B(net213),
    .Q(\line_cache[291][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25800_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01697_),
    .RESET_B(net218),
    .Q(\line_cache[291][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25801_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01698_),
    .RESET_B(net218),
    .Q(\line_cache[291][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25802_ (.CLK(clknet_leaf_69_clk_i),
    .D(net2160),
    .RESET_B(net213),
    .Q(\line_cache[291][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25803_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01700_),
    .RESET_B(net220),
    .Q(\line_cache[291][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25804_ (.CLK(clknet_leaf_67_clk_i),
    .D(net2041),
    .RESET_B(net214),
    .Q(\line_cache[291][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25805_ (.CLK(clknet_leaf_68_clk_i),
    .D(net2340),
    .RESET_B(net214),
    .Q(\line_cache[291][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25806_ (.CLK(clknet_leaf_70_clk_i),
    .D(net1827),
    .RESET_B(net218),
    .Q(\line_cache[291][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25807_ (.CLK(clknet_leaf_50_clk_i),
    .D(net2316),
    .RESET_B(net212),
    .Q(\line_cache[292][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25808_ (.CLK(clknet_leaf_52_clk_i),
    .D(net572),
    .RESET_B(net211),
    .Q(\line_cache[292][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25809_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01706_),
    .RESET_B(net213),
    .Q(\line_cache[292][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25810_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01707_),
    .RESET_B(net212),
    .Q(\line_cache[292][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25811_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01708_),
    .RESET_B(net213),
    .Q(\line_cache[292][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25812_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01709_),
    .RESET_B(net214),
    .Q(\line_cache[292][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25813_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01710_),
    .RESET_B(net211),
    .Q(\line_cache[292][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25814_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01711_),
    .RESET_B(net214),
    .Q(\line_cache[292][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25815_ (.CLK(clknet_leaf_50_clk_i),
    .D(net1420),
    .RESET_B(net212),
    .Q(\line_cache[293][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25816_ (.CLK(clknet_leaf_51_clk_i),
    .D(net2232),
    .RESET_B(net211),
    .Q(\line_cache[293][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25817_ (.CLK(clknet_leaf_67_clk_i),
    .D(net978),
    .RESET_B(net214),
    .Q(\line_cache[293][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25818_ (.CLK(clknet_leaf_51_clk_i),
    .D(net1656),
    .RESET_B(net212),
    .Q(\line_cache[293][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25819_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01716_),
    .RESET_B(net213),
    .Q(\line_cache[293][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25820_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01717_),
    .RESET_B(net206),
    .Q(\line_cache[293][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25821_ (.CLK(clknet_leaf_51_clk_i),
    .D(net2157),
    .RESET_B(net212),
    .Q(\line_cache[293][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25822_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01719_),
    .RESET_B(net206),
    .Q(\line_cache[293][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25823_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01720_),
    .RESET_B(net212),
    .Q(\line_cache[294][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25824_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01721_),
    .RESET_B(net211),
    .Q(\line_cache[294][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25825_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01722_),
    .RESET_B(net211),
    .Q(\line_cache[294][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25826_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01723_),
    .RESET_B(net213),
    .Q(\line_cache[294][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25827_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01724_),
    .RESET_B(net212),
    .Q(\line_cache[294][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25828_ (.CLK(clknet_leaf_67_clk_i),
    .D(net1000),
    .RESET_B(net214),
    .Q(\line_cache[294][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25829_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01726_),
    .RESET_B(net223),
    .Q(\line_cache[294][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25830_ (.CLK(clknet_leaf_66_clk_i),
    .D(net1060),
    .RESET_B(net211),
    .Q(\line_cache[294][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25831_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01728_),
    .RESET_B(net212),
    .Q(\line_cache[295][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25832_ (.CLK(clknet_leaf_66_clk_i),
    .D(net848),
    .RESET_B(net211),
    .Q(\line_cache[295][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25833_ (.CLK(clknet_leaf_66_clk_i),
    .D(net1675),
    .RESET_B(net211),
    .Q(\line_cache[295][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25834_ (.CLK(clknet_leaf_51_clk_i),
    .D(net1726),
    .RESET_B(net212),
    .Q(\line_cache[295][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25835_ (.CLK(clknet_leaf_50_clk_i),
    .D(net2269),
    .RESET_B(net212),
    .Q(\line_cache[295][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25836_ (.CLK(clknet_leaf_52_clk_i),
    .D(net2143),
    .RESET_B(net211),
    .Q(\line_cache[295][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25837_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01734_),
    .RESET_B(net211),
    .Q(\line_cache[295][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25838_ (.CLK(clknet_leaf_52_clk_i),
    .D(net2290),
    .RESET_B(net211),
    .Q(\line_cache[295][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25839_ (.CLK(clknet_leaf_54_clk_i),
    .D(net2211),
    .RESET_B(net209),
    .Q(\line_cache[296][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25840_ (.CLK(clknet_leaf_52_clk_i),
    .D(net1650),
    .RESET_B(net211),
    .Q(\line_cache[296][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25841_ (.CLK(clknet_leaf_54_clk_i),
    .D(net2288),
    .RESET_B(net207),
    .Q(\line_cache[296][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25842_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01739_),
    .RESET_B(net209),
    .Q(\line_cache[296][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25843_ (.CLK(clknet_leaf_55_clk_i),
    .D(net2235),
    .RESET_B(net209),
    .Q(\line_cache[296][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25844_ (.CLK(clknet_leaf_57_clk_i),
    .D(net3710),
    .RESET_B(net207),
    .Q(\line_cache[296][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25845_ (.CLK(clknet_leaf_57_clk_i),
    .D(net3809),
    .RESET_B(net207),
    .Q(\line_cache[296][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25846_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01743_),
    .RESET_B(net212),
    .Q(\line_cache[296][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25847_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01744_),
    .RESET_B(net209),
    .Q(\line_cache[297][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25848_ (.CLK(clknet_leaf_53_clk_i),
    .D(net1849),
    .RESET_B(net207),
    .Q(\line_cache[297][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25849_ (.CLK(clknet_leaf_58_clk_i),
    .D(net1176),
    .RESET_B(net208),
    .Q(\line_cache[297][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25850_ (.CLK(clknet_leaf_56_clk_i),
    .D(net1740),
    .RESET_B(net209),
    .Q(\line_cache[297][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25851_ (.CLK(clknet_leaf_55_clk_i),
    .D(net790),
    .RESET_B(net209),
    .Q(\line_cache[297][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25852_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01749_),
    .RESET_B(net205),
    .Q(\line_cache[297][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25853_ (.CLK(clknet_leaf_56_clk_i),
    .D(net1738),
    .RESET_B(net207),
    .Q(\line_cache[297][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25854_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01751_),
    .RESET_B(net208),
    .Q(\line_cache[297][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25855_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01752_),
    .RESET_B(net209),
    .Q(\line_cache[298][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25856_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01753_),
    .RESET_B(net208),
    .Q(\line_cache[298][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25857_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01754_),
    .RESET_B(net208),
    .Q(\line_cache[298][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25858_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01755_),
    .RESET_B(net210),
    .Q(\line_cache[298][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25859_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01756_),
    .RESET_B(net210),
    .Q(\line_cache[298][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25860_ (.CLK(clknet_leaf_58_clk_i),
    .D(net1777),
    .RESET_B(net208),
    .Q(\line_cache[298][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25861_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01758_),
    .RESET_B(net205),
    .Q(\line_cache[298][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25862_ (.CLK(clknet_leaf_53_clk_i),
    .D(net658),
    .RESET_B(net208),
    .Q(\line_cache[298][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25863_ (.CLK(clknet_leaf_51_clk_i),
    .D(net788),
    .RESET_B(net210),
    .Q(\line_cache[299][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25864_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01761_),
    .RESET_B(net208),
    .Q(\line_cache[299][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25865_ (.CLK(clknet_leaf_58_clk_i),
    .D(net1208),
    .RESET_B(net208),
    .Q(\line_cache[299][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25866_ (.CLK(clknet_leaf_55_clk_i),
    .D(net1703),
    .RESET_B(net209),
    .Q(\line_cache[299][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25867_ (.CLK(clknet_leaf_54_clk_i),
    .D(net1920),
    .RESET_B(net210),
    .Q(\line_cache[299][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25868_ (.CLK(clknet_leaf_54_clk_i),
    .D(net2300),
    .RESET_B(net208),
    .Q(\line_cache[299][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25869_ (.CLK(clknet_leaf_54_clk_i),
    .D(net1274),
    .RESET_B(net208),
    .Q(\line_cache[299][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25870_ (.CLK(clknet_leaf_54_clk_i),
    .D(net2192),
    .RESET_B(net210),
    .Q(\line_cache[299][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25871_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01784_),
    .RESET_B(net224),
    .Q(\line_cache[300][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25872_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01785_),
    .RESET_B(net224),
    .Q(\line_cache[300][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25873_ (.CLK(clknet_leaf_46_clk_i),
    .D(_01786_),
    .RESET_B(net224),
    .Q(\line_cache[300][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25874_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01787_),
    .RESET_B(net224),
    .Q(\line_cache[300][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25875_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01788_),
    .RESET_B(net210),
    .Q(\line_cache[300][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25876_ (.CLK(clknet_leaf_46_clk_i),
    .D(_01789_),
    .RESET_B(net225),
    .Q(\line_cache[300][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25877_ (.CLK(clknet_leaf_46_clk_i),
    .D(_01790_),
    .RESET_B(net224),
    .Q(\line_cache[300][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25878_ (.CLK(clknet_leaf_46_clk_i),
    .D(_01791_),
    .RESET_B(net224),
    .Q(\line_cache[300][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25879_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01792_),
    .RESET_B(net224),
    .Q(\line_cache[301][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25880_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01793_),
    .RESET_B(net224),
    .Q(\line_cache[301][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25881_ (.CLK(clknet_leaf_46_clk_i),
    .D(net1260),
    .RESET_B(net224),
    .Q(\line_cache[301][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25882_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01795_),
    .RESET_B(net226),
    .Q(\line_cache[301][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25883_ (.CLK(clknet_leaf_46_clk_i),
    .D(_01796_),
    .RESET_B(net226),
    .Q(\line_cache[301][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25884_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01797_),
    .RESET_B(net225),
    .Q(\line_cache[301][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25885_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01798_),
    .RESET_B(net226),
    .Q(\line_cache[301][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25886_ (.CLK(clknet_leaf_46_clk_i),
    .D(_01799_),
    .RESET_B(net226),
    .Q(\line_cache[301][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25887_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01800_),
    .RESET_B(net224),
    .Q(\line_cache[302][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25888_ (.CLK(clknet_leaf_43_clk_i),
    .D(_01801_),
    .RESET_B(net225),
    .Q(\line_cache[302][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25889_ (.CLK(clknet_leaf_47_clk_i),
    .D(_01802_),
    .RESET_B(net225),
    .Q(\line_cache[302][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25890_ (.CLK(clknet_leaf_47_clk_i),
    .D(net1969),
    .RESET_B(net225),
    .Q(\line_cache[302][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25891_ (.CLK(clknet_leaf_47_clk_i),
    .D(net554),
    .RESET_B(net226),
    .Q(\line_cache[302][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25892_ (.CLK(clknet_leaf_42_clk_i),
    .D(_01805_),
    .RESET_B(net226),
    .Q(\line_cache[302][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25893_ (.CLK(clknet_leaf_42_clk_i),
    .D(net1022),
    .RESET_B(net226),
    .Q(\line_cache[302][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25894_ (.CLK(clknet_leaf_47_clk_i),
    .D(net564),
    .RESET_B(net226),
    .Q(\line_cache[302][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25895_ (.CLK(clknet_leaf_44_clk_i),
    .D(net866),
    .RESET_B(net225),
    .Q(\line_cache[303][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25896_ (.CLK(clknet_leaf_44_clk_i),
    .D(net728),
    .RESET_B(net224),
    .Q(\line_cache[303][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25897_ (.CLK(clknet_leaf_44_clk_i),
    .D(net1144),
    .RESET_B(net225),
    .Q(\line_cache[303][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25898_ (.CLK(clknet_leaf_43_clk_i),
    .D(_01811_),
    .RESET_B(net225),
    .Q(\line_cache[303][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25899_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01812_),
    .RESET_B(net224),
    .Q(\line_cache[303][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25900_ (.CLK(clknet_leaf_44_clk_i),
    .D(net1948),
    .RESET_B(net224),
    .Q(\line_cache[303][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25901_ (.CLK(clknet_leaf_43_clk_i),
    .D(net986),
    .RESET_B(net225),
    .Q(\line_cache[303][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25902_ (.CLK(clknet_leaf_44_clk_i),
    .D(net1388),
    .RESET_B(net225),
    .Q(\line_cache[303][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25903_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01816_),
    .RESET_B(net194),
    .Q(\line_cache[304][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25904_ (.CLK(clknet_leaf_35_clk_i),
    .D(net1338),
    .RESET_B(net193),
    .Q(\line_cache[304][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25905_ (.CLK(clknet_leaf_35_clk_i),
    .D(net1972),
    .RESET_B(net193),
    .Q(\line_cache[304][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25906_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01819_),
    .RESET_B(net199),
    .Q(\line_cache[304][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25907_ (.CLK(clknet_leaf_37_clk_i),
    .D(_01820_),
    .RESET_B(net199),
    .Q(\line_cache[304][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25908_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01821_),
    .RESET_B(net199),
    .Q(\line_cache[304][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25909_ (.CLK(clknet_leaf_37_clk_i),
    .D(net3671),
    .RESET_B(net199),
    .Q(\line_cache[304][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25910_ (.CLK(clknet_leaf_40_clk_i),
    .D(net3816),
    .RESET_B(net231),
    .Q(\line_cache[304][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25911_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01824_),
    .RESET_B(net194),
    .Q(\line_cache[305][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25912_ (.CLK(clknet_leaf_35_clk_i),
    .D(net2419),
    .RESET_B(net193),
    .Q(\line_cache[305][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25913_ (.CLK(clknet_leaf_37_clk_i),
    .D(_01826_),
    .RESET_B(net202),
    .Q(\line_cache[305][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25914_ (.CLK(clknet_leaf_43_clk_i),
    .D(net2535),
    .RESET_B(net193),
    .Q(\line_cache[305][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25915_ (.CLK(clknet_leaf_35_clk_i),
    .D(_01828_),
    .RESET_B(net203),
    .Q(\line_cache[305][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25916_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01829_),
    .RESET_B(net202),
    .Q(\line_cache[305][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25917_ (.CLK(clknet_leaf_43_clk_i),
    .D(net2187),
    .RESET_B(net231),
    .Q(\line_cache[305][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25918_ (.CLK(clknet_leaf_40_clk_i),
    .D(_01831_),
    .RESET_B(net231),
    .Q(\line_cache[305][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25919_ (.CLK(clknet_leaf_44_clk_i),
    .D(net972),
    .RESET_B(net203),
    .Q(\line_cache[306][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25920_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01833_),
    .RESET_B(net194),
    .Q(\line_cache[306][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25921_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01834_),
    .RESET_B(net194),
    .Q(\line_cache[306][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25922_ (.CLK(clknet_leaf_35_clk_i),
    .D(net1576),
    .RESET_B(net193),
    .Q(\line_cache[306][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25923_ (.CLK(clknet_leaf_32_clk_i),
    .D(net740),
    .RESET_B(net193),
    .Q(\line_cache[306][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25924_ (.CLK(clknet_leaf_35_clk_i),
    .D(net1547),
    .RESET_B(net203),
    .Q(\line_cache[306][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25925_ (.CLK(clknet_leaf_35_clk_i),
    .D(net1875),
    .RESET_B(net193),
    .Q(\line_cache[306][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25926_ (.CLK(clknet_leaf_33_clk_i),
    .D(net1404),
    .RESET_B(net194),
    .Q(\line_cache[306][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25927_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01840_),
    .RESET_B(net194),
    .Q(\line_cache[307][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25928_ (.CLK(clknet_leaf_34_clk_i),
    .D(net1006),
    .RESET_B(net203),
    .Q(\line_cache[307][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25929_ (.CLK(clknet_leaf_34_clk_i),
    .D(_01842_),
    .RESET_B(net194),
    .Q(\line_cache[307][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25930_ (.CLK(clknet_leaf_31_clk_i),
    .D(net1038),
    .RESET_B(net193),
    .Q(\line_cache[307][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25931_ (.CLK(clknet_leaf_32_clk_i),
    .D(net730),
    .RESET_B(net193),
    .Q(\line_cache[307][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25932_ (.CLK(clknet_leaf_37_clk_i),
    .D(net1742),
    .RESET_B(net203),
    .Q(\line_cache[307][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25933_ (.CLK(clknet_leaf_35_clk_i),
    .D(_01846_),
    .RESET_B(net193),
    .Q(\line_cache[307][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25934_ (.CLK(clknet_leaf_33_clk_i),
    .D(_01847_),
    .RESET_B(net194),
    .Q(\line_cache[307][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25935_ (.CLK(clknet_leaf_34_clk_i),
    .D(net2343),
    .RESET_B(net194),
    .Q(\line_cache[308][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25936_ (.CLK(clknet_leaf_56_clk_i),
    .D(net1306),
    .RESET_B(net207),
    .Q(\line_cache[308][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25937_ (.CLK(clknet_leaf_55_clk_i),
    .D(net2352),
    .RESET_B(net209),
    .Q(\line_cache[308][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25938_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01851_),
    .RESET_B(net209),
    .Q(\line_cache[308][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25939_ (.CLK(clknet_leaf_55_clk_i),
    .D(net1606),
    .RESET_B(net209),
    .Q(\line_cache[308][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25940_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01853_),
    .RESET_B(net172),
    .Q(\line_cache[308][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25941_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01854_),
    .RESET_B(net207),
    .Q(\line_cache[308][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25942_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01855_),
    .RESET_B(net207),
    .Q(\line_cache[308][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25943_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01856_),
    .RESET_B(net173),
    .Q(\line_cache[309][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25944_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01857_),
    .RESET_B(net172),
    .Q(\line_cache[309][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25945_ (.CLK(clknet_leaf_56_clk_i),
    .D(net1020),
    .RESET_B(net207),
    .Q(\line_cache[309][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25946_ (.CLK(clknet_leaf_56_clk_i),
    .D(net2384),
    .RESET_B(net209),
    .Q(\line_cache[309][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25947_ (.CLK(clknet_leaf_55_clk_i),
    .D(net1314),
    .RESET_B(net209),
    .Q(\line_cache[309][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25948_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01861_),
    .RESET_B(net172),
    .Q(\line_cache[309][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25949_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01862_),
    .RESET_B(net207),
    .Q(\line_cache[309][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25950_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01863_),
    .RESET_B(net207),
    .Q(\line_cache[309][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25951_ (.CLK(clknet_leaf_45_clk_i),
    .D(_01872_),
    .RESET_B(net194),
    .Q(\line_cache[310][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25952_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01873_),
    .RESET_B(net207),
    .Q(\line_cache[310][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25953_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01874_),
    .RESET_B(net205),
    .Q(\line_cache[310][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25954_ (.CLK(clknet_leaf_56_clk_i),
    .D(net1358),
    .RESET_B(net209),
    .Q(\line_cache[310][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25955_ (.CLK(clknet_leaf_45_clk_i),
    .D(net1625),
    .RESET_B(net209),
    .Q(\line_cache[310][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25956_ (.CLK(clknet_leaf_22_clk_i),
    .D(net1470),
    .RESET_B(net172),
    .Q(\line_cache[310][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25957_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01878_),
    .RESET_B(net207),
    .Q(\line_cache[310][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25958_ (.CLK(clknet_leaf_56_clk_i),
    .D(net1048),
    .RESET_B(net207),
    .Q(\line_cache[310][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25959_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01880_),
    .RESET_B(net194),
    .Q(\line_cache[311][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25960_ (.CLK(clknet_leaf_57_clk_i),
    .D(net1090),
    .RESET_B(net207),
    .Q(\line_cache[311][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25961_ (.CLK(clknet_leaf_56_clk_i),
    .D(net1210),
    .RESET_B(net207),
    .Q(\line_cache[311][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25962_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01883_),
    .RESET_B(net209),
    .Q(\line_cache[311][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25963_ (.CLK(clknet_leaf_23_clk_i),
    .D(net1416),
    .RESET_B(net173),
    .Q(\line_cache[311][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25964_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01885_),
    .RESET_B(net172),
    .Q(\line_cache[311][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25965_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01886_),
    .RESET_B(net205),
    .Q(\line_cache[311][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25966_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01887_),
    .RESET_B(net173),
    .Q(\line_cache[311][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25967_ (.CLK(clknet_leaf_34_clk_i),
    .D(net1974),
    .RESET_B(net194),
    .Q(\line_cache[312][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25968_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01889_),
    .RESET_B(net201),
    .Q(\line_cache[312][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25969_ (.CLK(clknet_leaf_35_clk_i),
    .D(net1642),
    .RESET_B(net202),
    .Q(\line_cache[312][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25970_ (.CLK(clknet_leaf_288_clk_i),
    .D(_01891_),
    .RESET_B(net199),
    .Q(\line_cache[312][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25971_ (.CLK(clknet_leaf_36_clk_i),
    .D(net1174),
    .RESET_B(net199),
    .Q(\line_cache[312][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25972_ (.CLK(clknet_leaf_36_clk_i),
    .D(net3669),
    .RESET_B(net199),
    .Q(\line_cache[312][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25973_ (.CLK(clknet_leaf_37_clk_i),
    .D(net3757),
    .RESET_B(net199),
    .Q(\line_cache[312][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25974_ (.CLK(clknet_leaf_36_clk_i),
    .D(net818),
    .RESET_B(net199),
    .Q(\line_cache[312][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25975_ (.CLK(clknet_leaf_31_clk_i),
    .D(net746),
    .RESET_B(net193),
    .Q(\line_cache[313][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25976_ (.CLK(clknet_leaf_37_clk_i),
    .D(net2185),
    .RESET_B(net202),
    .Q(\line_cache[313][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25977_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01898_),
    .RESET_B(net202),
    .Q(\line_cache[313][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25978_ (.CLK(clknet_leaf_36_clk_i),
    .D(net2086),
    .RESET_B(net199),
    .Q(\line_cache[313][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25979_ (.CLK(clknet_leaf_288_clk_i),
    .D(_01900_),
    .RESET_B(net199),
    .Q(\line_cache[313][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25980_ (.CLK(clknet_leaf_38_clk_i),
    .D(_01901_),
    .RESET_B(net202),
    .Q(\line_cache[313][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25981_ (.CLK(clknet_leaf_36_clk_i),
    .D(net1378),
    .RESET_B(net199),
    .Q(\line_cache[313][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25982_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01903_),
    .RESET_B(net200),
    .Q(\line_cache[313][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25983_ (.CLK(clknet_leaf_31_clk_i),
    .D(net576),
    .RESET_B(net193),
    .Q(\line_cache[314][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25984_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01905_),
    .RESET_B(net200),
    .Q(\line_cache[314][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25985_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01906_),
    .RESET_B(net201),
    .Q(\line_cache[314][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25986_ (.CLK(clknet_leaf_288_clk_i),
    .D(net1797),
    .RESET_B(net199),
    .Q(\line_cache[314][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25987_ (.CLK(clknet_leaf_31_clk_i),
    .D(net2059),
    .RESET_B(net193),
    .Q(\line_cache[314][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25988_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01909_),
    .RESET_B(net200),
    .Q(\line_cache[314][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25989_ (.CLK(clknet_leaf_36_clk_i),
    .D(net1142),
    .RESET_B(net193),
    .Q(\line_cache[314][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25990_ (.CLK(clknet_leaf_288_clk_i),
    .D(net1615),
    .RESET_B(net199),
    .Q(\line_cache[314][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25991_ (.CLK(clknet_leaf_288_clk_i),
    .D(_01912_),
    .RESET_B(net195),
    .Q(\line_cache[315][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25992_ (.CLK(clknet_leaf_286_clk_i),
    .D(_01913_),
    .RESET_B(net200),
    .Q(\line_cache[315][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25993_ (.CLK(clknet_leaf_37_clk_i),
    .D(net698),
    .RESET_B(net199),
    .Q(\line_cache[315][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25994_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01915_),
    .RESET_B(net200),
    .Q(\line_cache[315][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25995_ (.CLK(clknet_leaf_31_clk_i),
    .D(net1436),
    .RESET_B(net193),
    .Q(\line_cache[315][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25996_ (.CLK(clknet_leaf_287_clk_i),
    .D(_01917_),
    .RESET_B(net200),
    .Q(\line_cache[315][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25997_ (.CLK(clknet_leaf_31_clk_i),
    .D(net830),
    .RESET_B(net193),
    .Q(\line_cache[315][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25998_ (.CLK(clknet_leaf_288_clk_i),
    .D(net2088),
    .RESET_B(net199),
    .Q(\line_cache[315][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25999_ (.CLK(clknet_leaf_288_clk_i),
    .D(net2701),
    .RESET_B(net195),
    .Q(\line_cache[316][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26000_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01921_),
    .RESET_B(net195),
    .Q(\line_cache[316][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26001_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01922_),
    .RESET_B(net191),
    .Q(\line_cache[316][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26002_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01923_),
    .RESET_B(net195),
    .Q(\line_cache[316][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26003_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01924_),
    .RESET_B(net197),
    .Q(\line_cache[316][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26004_ (.CLK(clknet_leaf_294_clk_i),
    .D(net3627),
    .RESET_B(net198),
    .Q(\line_cache[316][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26005_ (.CLK(clknet_leaf_288_clk_i),
    .D(net3724),
    .RESET_B(net198),
    .Q(\line_cache[316][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26006_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01927_),
    .RESET_B(net198),
    .Q(\line_cache[316][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26007_ (.CLK(clknet_leaf_289_clk_i),
    .D(net672),
    .RESET_B(net197),
    .Q(\line_cache[317][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26008_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01929_),
    .RESET_B(net195),
    .Q(\line_cache[317][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26009_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01930_),
    .RESET_B(net198),
    .Q(\line_cache[317][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26010_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01931_),
    .RESET_B(net195),
    .Q(\line_cache[317][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26011_ (.CLK(clknet_leaf_289_clk_i),
    .D(net1132),
    .RESET_B(net197),
    .Q(\line_cache[317][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26012_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01933_),
    .RESET_B(net197),
    .Q(\line_cache[317][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26013_ (.CLK(clknet_leaf_294_clk_i),
    .D(net2517),
    .RESET_B(net198),
    .Q(\line_cache[317][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26014_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01935_),
    .RESET_B(net198),
    .Q(\line_cache[317][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26015_ (.CLK(clknet_leaf_288_clk_i),
    .D(net476),
    .RESET_B(net198),
    .Q(\line_cache[318][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26016_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01937_),
    .RESET_B(net195),
    .Q(\line_cache[318][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26017_ (.CLK(clknet_leaf_294_clk_i),
    .D(net1040),
    .RESET_B(net191),
    .Q(\line_cache[318][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26018_ (.CLK(clknet_leaf_288_clk_i),
    .D(_01939_),
    .RESET_B(net197),
    .Q(\line_cache[318][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26019_ (.CLK(clknet_leaf_290_clk_i),
    .D(net780),
    .RESET_B(net196),
    .Q(\line_cache[318][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26020_ (.CLK(clknet_leaf_289_clk_i),
    .D(_01941_),
    .RESET_B(net197),
    .Q(\line_cache[318][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26021_ (.CLK(clknet_leaf_292_clk_i),
    .D(_01942_),
    .RESET_B(net196),
    .Q(\line_cache[318][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26022_ (.CLK(clknet_leaf_290_clk_i),
    .D(net1694),
    .RESET_B(net197),
    .Q(\line_cache[318][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26023_ (.CLK(clknet_leaf_30_clk_i),
    .D(net484),
    .RESET_B(net192),
    .Q(\line_cache[319][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26024_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01945_),
    .RESET_B(net192),
    .Q(\line_cache[319][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26025_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01946_),
    .RESET_B(net192),
    .Q(\line_cache[319][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26026_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01947_),
    .RESET_B(net195),
    .Q(\line_cache[319][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26027_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01948_),
    .RESET_B(net191),
    .Q(\line_cache[319][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26028_ (.CLK(clknet_leaf_295_clk_i),
    .D(_01949_),
    .RESET_B(net191),
    .Q(\line_cache[319][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26029_ (.CLK(clknet_leaf_294_clk_i),
    .D(_01950_),
    .RESET_B(net192),
    .Q(\line_cache[319][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26030_ (.CLK(clknet_leaf_293_clk_i),
    .D(_01951_),
    .RESET_B(net195),
    .Q(\line_cache[319][7] ));
 sky130_fd_sc_hd__buf_1 _26067_ (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_108_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_109_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_110_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_111_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_112_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_113_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_114_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_115_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_116_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_117_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_118_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_119_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_120_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_121_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_122_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_123_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_124_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_125_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_126_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_127_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_128_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_129_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_130_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_131_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_132_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_133_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_134_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_135_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_136_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_137_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_138_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_139_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_140_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_141_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_142_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_143_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_144_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_145_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_146_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_147_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_148_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_149_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_150_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_151_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_152_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_153_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_154_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_155_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_156_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_157_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_158_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_159_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_160_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_161_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_162_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_163_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_164_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_165_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_166_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_167_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_168_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_169_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_170_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_171_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_172_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_173_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_174_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_175_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_176_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_177_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_178_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_179_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_180_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_181_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_182_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_183_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_184_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_185_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_186_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_187_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_188_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_189_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_190_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_191_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_192_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_193_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_194_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_195_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_196_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_197_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_198_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_199_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_200_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_201_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_202_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_203_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_204_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_205_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_206_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_207_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_208_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_209_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_210_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_211_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_212_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_213_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_214_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_215_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_216_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_217_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_218_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_219_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_220_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_221_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_222_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_223_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_224_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_225_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_226_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_227_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_228_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_229_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_230_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_231_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_232_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_233_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_234_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_235_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_236_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_237_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_238_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_239_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_240_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_241_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_242_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_243_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_244_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_245_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_246_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_247_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_248_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_249_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_250_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_251_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_252_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_253_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_254_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_255_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_256_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_257_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_258_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_259_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_260_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_261_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_262_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_263_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_264_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_265_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_266_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_267_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_268_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_269_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_270_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_271_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_272_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_273_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_274_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_275_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_276_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_277_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_278_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_279_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_280_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_281_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_282_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_283_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_284_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_285_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_286_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_287_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_288_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_289_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_290_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_291_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_292_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_293_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_294_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_295_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_296_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_297_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_298_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_299_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_300_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_301_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_301_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_302_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_303_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_303_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_304_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_304_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_305_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_305_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_306_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_306_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_307_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_307_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_308_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_308_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_309_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_309_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_310_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_310_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_311_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_311_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_312_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_312_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_313_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_313_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_314_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_314_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_315_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_315_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_316_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_316_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_317_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_317_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_318_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_318_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_319_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_319_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_320_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_320_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_321_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_321_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_322_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_322_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_323_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_323_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_324_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_324_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_325_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_325_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_326_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_326_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_327_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_327_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_328_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_328_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_329_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_329_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_330_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_330_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_331_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_331_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_332_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_332_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout147 (.A(net154),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_8 fanout148 (.A(net154),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net154),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_8 fanout150 (.A(net154),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net154),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_8 fanout152 (.A(net154),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(net174),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_8 fanout155 (.A(net158),
    .X(net155));
 sky130_fd_sc_hd__buf_4 fanout156 (.A(net158),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(net174),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_8 fanout159 (.A(net161),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_8 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(net174),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(net165),
    .X(net162));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(net165),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net174),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_6 fanout168 (.A(net174),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net171),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_8 fanout171 (.A(net174),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net252),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_8 fanout175 (.A(net189),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net189),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net189),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(net189),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(net189),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_8 fanout182 (.A(net189),
    .X(net182));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net189),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout184 (.A(net189),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net189),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_8 fanout186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_8 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(net252),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout190 (.A(net192),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(net203),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_8 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 fanout194 (.A(net203),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(net198),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_8 fanout196 (.A(net198),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 fanout198 (.A(net203),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 fanout199 (.A(net202),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout200 (.A(net202),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net252),
    .X(net203));
 sky130_fd_sc_hd__buf_6 fanout204 (.A(net223),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net223),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(net223),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_8 fanout207 (.A(net210),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net210),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(net223),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net214),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(net214),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(net223),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_8 fanout215 (.A(net217),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net223),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(net221),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_8 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_8 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_6 fanout223 (.A(net252),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_8 fanout224 (.A(net226),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net252),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_8 fanout227 (.A(net230),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(net230),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net252),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 fanout231 (.A(net239),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net239),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 fanout233 (.A(net239),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net239),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_8 fanout235 (.A(net239),
    .X(net235));
 sky130_fd_sc_hd__buf_2 fanout236 (.A(net239),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_8 fanout237 (.A(net239),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net252),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_8 fanout240 (.A(net242),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_8 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_8 fanout242 (.A(net251),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_8 fanout243 (.A(net251),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net251),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_8 fanout245 (.A(net251),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net251),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_8 fanout247 (.A(net251),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 fanout248 (.A(net251),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_8 fanout249 (.A(net251),
    .X(net249));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_8 fanout252 (.A(net83),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 fanout253 (.A(net261),
    .X(net253));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net261),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_8 fanout255 (.A(net261),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(net261),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_8 fanout257 (.A(net261),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 fanout258 (.A(net261),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_8 fanout259 (.A(net261),
    .X(net259));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(net284),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 fanout262 (.A(net284),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_4 fanout263 (.A(net284),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_8 fanout264 (.A(net284),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(net284),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_8 fanout266 (.A(net269),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 fanout267 (.A(net269),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_8 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net284),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(net284),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_8 fanout272 (.A(net284),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_8 fanout273 (.A(net275),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_8 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(net284),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_8 fanout276 (.A(net279),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_8 fanout277 (.A(net279),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(net284),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_8 fanout280 (.A(net283),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_8 fanout281 (.A(net283),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__buf_4 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_6 fanout284 (.A(net370),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(net299),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 fanout286 (.A(net299),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_8 fanout287 (.A(net299),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(net299),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_8 fanout289 (.A(net292),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_4 fanout290 (.A(net292),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_8 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(net299),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_8 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_4 fanout294 (.A(net299),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_8 fanout295 (.A(net299),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net299),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_8 fanout297 (.A(net299),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_4 fanout299 (.A(net370),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_8 fanout300 (.A(net307),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_8 fanout301 (.A(net307),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 fanout302 (.A(net307),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_8 fanout303 (.A(net307),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net307),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_8 fanout305 (.A(net307),
    .X(net305));
 sky130_fd_sc_hd__buf_4 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__buf_4 fanout307 (.A(net370),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_8 fanout308 (.A(net315),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_8 fanout309 (.A(net315),
    .X(net309));
 sky130_fd_sc_hd__buf_4 fanout310 (.A(net315),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_8 fanout311 (.A(net315),
    .X(net311));
 sky130_fd_sc_hd__buf_2 fanout312 (.A(net315),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_8 fanout313 (.A(net315),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_4 fanout315 (.A(net370),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_8 fanout316 (.A(net319),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_8 fanout317 (.A(net319),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 fanout319 (.A(net344),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_8 fanout320 (.A(net323),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_8 fanout321 (.A(net323),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(net344),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_8 fanout324 (.A(net327),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_8 fanout325 (.A(net327),
    .X(net325));
 sky130_fd_sc_hd__buf_4 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 fanout327 (.A(net344),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_8 fanout328 (.A(net344),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_4 fanout329 (.A(net344),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_8 fanout330 (.A(net344),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_4 fanout331 (.A(net344),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_8 fanout332 (.A(net334),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_8 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_8 fanout334 (.A(net343),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_8 fanout335 (.A(net343),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_8 fanout336 (.A(net343),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_8 fanout337 (.A(net343),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_4 fanout338 (.A(net343),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_8 fanout339 (.A(net343),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 fanout340 (.A(net343),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_8 fanout341 (.A(net343),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_8 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_8 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__buf_4 fanout344 (.A(net370),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_8 fanout345 (.A(net348),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 fanout346 (.A(net348),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_8 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_4 fanout348 (.A(net361),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_8 fanout349 (.A(net361),
    .X(net349));
 sky130_fd_sc_hd__buf_2 fanout350 (.A(net361),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_8 fanout351 (.A(net361),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_4 fanout352 (.A(net361),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_8 fanout353 (.A(net361),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 fanout354 (.A(net361),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_8 fanout355 (.A(net361),
    .X(net355));
 sky130_fd_sc_hd__buf_4 fanout356 (.A(net361),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_8 fanout357 (.A(net360),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_8 fanout358 (.A(net360),
    .X(net358));
 sky130_fd_sc_hd__buf_4 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_4 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_4 fanout361 (.A(net370),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_8 fanout362 (.A(net365),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_8 fanout363 (.A(net365),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_4 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_8 fanout366 (.A(net370),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_8 fanout367 (.A(net369),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_8 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_4 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_8 fanout370 (.A(net83),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\line_cache[126][4] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00194_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_01779_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_00433_),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\line_cache[36][0] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_01992_),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\line_cache[280][1] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_01601_),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\line_cache[124][2] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_00218_),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\line_cache[236][2] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_01210_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\line_cache[311][4] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\line_cache[106][0] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_01884_),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\line_cache[266][4] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_01476_),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\line_cache[293][0] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_01712_),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\line_cache[167][2] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_00594_),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\line_cache[79][3] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_02371_),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\line_cache[208][5] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_00056_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_00965_),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\line_cache[164][0] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_00568_),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\line_cache[29][0] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_01768_),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\line_cache[71][6] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_02310_),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\line_cache[61][6] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_02222_),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\line_cache[315][4] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\line_cache[267][0] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_01916_),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\line_cache[135][2] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_00314_),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\line_cache[209][0] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_00968_),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\line_cache[249][6] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_01326_),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\line_cache[107][1] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_00065_),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\line_cache[121][6] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_01480_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_00198_),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\line_cache[267][7] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_01487_),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\line_cache[247][1] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_01305_),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\line_cache[238][6] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_01230_),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\line_cache[180][5] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_00717_),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\line_cache[205][2] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\line_cache[226][0] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_00938_),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\line_cache[285][6] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_01646_),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\line_cache[142][7] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_00383_),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\line_cache[155][2] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_00490_),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\line_cache[28][4] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_01684_),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\line_cache[127][6] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_01120_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_00246_),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\line_cache[126][0] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_00232_),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\line_cache[310][5] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_01877_),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\line_cache[196][0] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_00848_),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\line_cache[289][4] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_01676_),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\line_cache[281][2] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\line_cache[258][0] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_01610_),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\line_cache[40][4] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_02036_),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\line_cache[155][3] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_00491_),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\line_cache[173][4] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_00652_),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\line_cache[290][0] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_01688_),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\line_cache[155][6] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_01400_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_00494_),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\line_cache[13][4] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_00356_),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\line_cache[16][1] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_00617_),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\line_cache[36][2] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_01994_),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\line_cache[178][7] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_00695_),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\line_cache[62][6] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\line_cache[133][3] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_02230_),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\line_cache[187][0] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_00768_),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\line_cache[43][6] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_02062_),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\line_cache[72][7] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_02319_),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\line_cache[237][0] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_01216_),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\line_cache[172][7] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\line_cache[243][2] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_00299_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_00647_),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\line_cache[289][6] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_01678_),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\line_cache[140][1] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_00361_),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\line_cache[83][5] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_02413_),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\line_cache[173][0] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_00648_),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\line_cache[137][4] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\line_cache[12][7] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_00332_),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\line_cache[138][3] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_00339_),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\line_cache[24][4] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_01332_),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\line_cache[78][5] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_02365_),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\line_cache[240][2] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_01250_),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\line_cache[215][7] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_00271_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_01031_),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\line_cache[250][7] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_01343_),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\line_cache[157][0] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_00504_),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\line_cache[146][4] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_00412_),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\line_cache[39][0] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_02016_),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\line_cache[59][6] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\line_cache[229][4] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_02198_),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\line_cache[14][7] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_00447_),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\line_cache[196][4] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_00852_),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\line_cache[55][0] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_02160_),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\line_cache[103][6] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\line_cache[11][2] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(_00178_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_01148_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\line_cache[306][5] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(_01837_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(\line_cache[231][4] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(_01172_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\line_cache[67][6] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(_02270_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\line_cache[85][0] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(_02424_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\line_cache[81][6] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(_02398_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\line_cache[224][1] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\line_cache[111][3] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(_00107_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\line_cache[227][6] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(_01134_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\line_cache[86][7] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(_02439_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\line_cache[55][7] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(_02167_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\line_cache[73][6] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(_02326_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_01105_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\line_cache[124][4] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(_00220_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\line_cache[136][1] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(_00321_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\line_cache[102][3] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\line_cache[174][5] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_00661_),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\line_cache[223][1] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_01097_),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\line_cache[306][3] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\line_cache[241][0] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_01835_),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\line_cache[71][7] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_02311_),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\line_cache[238][3] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_01227_),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\line_cache[155][1] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(_00489_),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\line_cache[100][4] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_00012_),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\line_cache[132][5] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_01256_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_00293_),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\line_cache[12][0] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_00264_),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\line_cache[32][5] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_01965_),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\line_cache[188][5] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_00781_),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\line_cache[162][3] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_00555_),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\line_cache[231][5] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\line_cache[259][6] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_01173_),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\line_cache[23][1] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_01241_),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\line_cache[174][4] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_00660_),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\line_cache[104][7] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_00047_),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\line_cache[225][3] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_01115_),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\line_cache[308][4] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_01274_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_01414_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_01852_),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\line_cache[268][7] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_01495_),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\line_cache[11][1] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(\line_cache[106][3] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(_00059_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\line_cache[180][4] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(_00716_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\line_cache[314][7] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(_01911_),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\line_cache[243][7] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\line_cache[94][4] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(_02508_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\line_cache[284][5] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(_01637_),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\line_cache[152][7] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(_00471_),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\line_cache[155][4] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(_00492_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\line_cache[310][4] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(_01876_),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_01279_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\line_cache[275][1] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(_01553_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\line_cache[236][1] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(_01209_),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\line_cache[188][0] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\line_cache[18][0] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_00792_),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\line_cache[123][4] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_00212_),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\line_cache[139][4] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\line_cache[206][4] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_00348_),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\line_cache[172][5] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_00645_),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\line_cache[97][0] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_02528_),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\line_cache[312][2] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_01890_),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\line_cache[55][1] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_02161_),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\line_cache[28][7] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_00948_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_01687_),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\line_cache[35][2] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_01986_),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\line_cache[296][1] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_01737_),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\line_cache[96][1] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_02521_),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\line_cache[256][4] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_01388_),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\line_cache[293][3] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\line_cache[3][6] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_01715_),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\line_cache[123][5] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_00213_),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\line_cache[154][4] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_00484_),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\line_cache[249][3] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_01323_),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\line_cache[199][2] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_00874_),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\line_cache[3][4] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_02030_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_02028_),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\line_cache[117][6] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_00158_),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\line_cache[110][6] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_00102_),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\line_cache[28][5] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_01685_),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\line_cache[284][4] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\line_cache[295][2] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(_01730_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\line_cache[212][2] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\line_cache[8][7] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(_02471_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(\line_cache[221][6] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(_01086_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(\line_cache[27][6] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(_01598_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\line_cache[208][4] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(_00964_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\line_cache[64][4] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(_02244_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_01002_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\line_cache[95][1] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(_02513_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\line_cache[88][1] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\line_cache[108][5] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_00077_),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\line_cache[234][3] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_01195_),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\line_cache[318][7] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(_01943_),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\line_cache[310][0] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\line_cache[242][5] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\line_cache[290][6] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(_01694_),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\line_cache[249][1] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(_01321_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\line_cache[247][3] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(_01307_),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\line_cache[299][3] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(_01763_),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\line_cache[119][6] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(_00174_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\line_cache[189][2] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_01269_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\line_cache[240][0] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\line_cache[152][4] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_00468_),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\line_cache[116][1] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(_00145_),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\line_cache[256][0] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(_01384_),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\line_cache[99][2] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(_02546_),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\line_cache[175][5] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\line_cache[239][6] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(_00669_),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\line_cache[237][2] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(_01218_),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\line_cache[151][0] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(_00456_),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\line_cache[152][1] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(_00465_),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\line_cache[139][3] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(_00347_),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\line_cache[295][3] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_01238_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(_01731_),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\line_cache[222][5] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(_01093_),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\line_cache[26][6] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(_01510_),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\line_cache[11][4] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(_00180_),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\line_cache[55][5] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_02165_),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\line_cache[270][3] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\line_cache[104][4] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(_01515_),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\line_cache[297][6] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(_01750_),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\line_cache[297][3] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_01747_),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\line_cache[307][5] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_01845_),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\line_cache[83][1] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(_02409_),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\line_cache[0][2] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_00044_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(_00002_),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\line_cache[17][0] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(_00704_),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\line_cache[94][6] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(_02510_),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\line_cache[174][6] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(_00662_),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\line_cache[37][3] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(_02003_),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\line_cache[254][4] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\line_cache[241][1] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(_01372_),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\line_cache[103][7] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(_00039_),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\line_cache[198][5] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(_00869_),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\line_cache[54][6] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(_02158_),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\line_cache[76][5] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(_02349_),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\line_cache[116][4] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_01257_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_00148_),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\line_cache[95][0] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_02512_),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\line_cache[288][5] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_01669_),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\line_cache[119][5] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_00173_),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\line_cache[179][0] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_00696_),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\line_cache[201][0] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\line_cache[239][4] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(\line_cache[298][5] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(_01757_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\line_cache[200][2] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(_00898_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(\line_cache[28][2] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(_01682_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(\line_cache[92][4] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(_02492_),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\line_cache[13][6] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(_00358_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_01236_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\line_cache[185][6] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\line_cache[129][0] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(_00256_),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\line_cache[185][4] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(_00756_),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\line_cache[117][0] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(_00152_),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\line_cache[123][2] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\line_cache[289][2] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(_01674_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\line_cache[225][2] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\line_cache[314][3] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(_01907_),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\line_cache[251][7] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(_01351_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\line_cache[183][2] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\line_cache[88][2] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(_02450_),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\line_cache[233][4] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\line_cache[220][5] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(_01077_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00786_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_01114_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(\line_cache[121][0] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(_00192_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(\line_cache[57][0] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(_02176_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(\line_cache[185][1] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(_00753_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\line_cache[318][5] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\line_cache[218][5] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(_01053_),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\line_cache[281][6] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\line_cache[212][0] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_01614_),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\line_cache[209][6] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_00974_),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\line_cache[236][5] ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(_01213_),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\line_cache[162][5] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(\line_cache[34][3] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(_01979_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\line_cache[221][2] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(_01082_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_01000_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\line_cache[291][7] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(_01703_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\line_cache[110][0] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(_00096_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\line_cache[257][2] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(_01394_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\line_cache[13][0] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(_00352_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\line_cache[133][0] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(_00296_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\line_cache[242][0] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(\line_cache[199][1] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\line_cache[214][6] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(_01022_),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\line_cache[303][4] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(\line_cache[122][4] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(_00204_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(\line_cache[25][2] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(_01418_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\line_cache[197][4] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\line_cache[53][3] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_01264_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(_02147_),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\line_cache[145][2] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\line_cache[297][1] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(_01745_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\line_cache[130][5] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(_00277_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\line_cache[316][1] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\line_cache[118][3] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_00163_),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\line_cache[158][0] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\line_cache[224][4] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(\line_cache[266][6] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\line_cache[104][0] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(_00040_),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\res_h_counter[9] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(_02706_),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\line_cache[177][6] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(\line_cache[116][5] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(_00149_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\line_cache[14][5] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(_00445_),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_01108_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(\line_cache[250][4] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(_01340_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\line_cache[110][4] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(_00100_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(\line_cache[177][3] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\line_cache[10][6] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(\line_cache[9][1] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(_02553_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(\line_cache[306][6] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(_01838_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\line_cache[302][4] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(\pixel_double_counter[3] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(_08495_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(_02728_),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\line_cache[17][3] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(_00707_),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\line_cache[153][1] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(_00473_),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\line_cache[60][7] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(_02215_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\line_cache[172][4] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_01804_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(_00644_),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\line_cache[284][7] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\line_cache[89][6] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(_02462_),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\line_cache[39][3] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(_02019_),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\line_cache[23][0] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(_01240_),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(\line_cache[161][6] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(_00550_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\line_cache[213][1] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(\line_cache[122][5] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(_00205_),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\line_cache[249][2] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(_01322_),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\line_cache[99][5] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(_02549_),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\line_cache[103][0] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(_00032_),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\line_cache[142][6] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(_00382_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\line_cache[214][7] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_01009_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\line_cache[76][4] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(_02348_),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\line_cache[289][3] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(_01675_),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\line_cache[274][6] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(_01550_),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\pixel_double_counter[2] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(_08491_),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(_02727_),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\line_cache[153][2] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\line_cache[267][6] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(_00474_),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\line_cache[49][3] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(_02107_),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\line_cache[299][4] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(_01764_),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\line_cache[135][6] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\line_cache[20][1] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(_00977_),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\line_cache[89][4] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(_02460_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_01486_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\line_cache[247][2] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(_01306_),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\line_cache[100][1] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(_00009_),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\line_cache[190][4] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(_00804_),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\line_cache[274][3] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(_01547_),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\line_cache[67][7] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(_02271_),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\line_cache[211][7] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(\line_cache[93][2] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(_02498_),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(\line_cache[182][7] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\line_cache[215][4] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(_01028_),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(\line_cache[158][4] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(\line_cache[300][2] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\line_cache[208][0] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(_00960_),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(\line_cache[240][1] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_00999_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(_01249_),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(\line_cache[303][5] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(_01813_),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\line_cache[202][4] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_00916_),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\line_cache[158][3] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(_00515_),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\line_cache[257][0] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(_01392_),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(\line_cache[60][0] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\line_cache[125][3] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\line_cache[142][3] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\line_cache[8][1] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(_02465_),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\line_cache[210][7] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_00991_),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\line_cache[301][0] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(\line_cache[210][5] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(_00989_),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\line_cache[48][5] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(_02101_),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_00227_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\line_cache[173][1] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(_00649_),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\line_cache[302][3] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(_01803_),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(\line_cache[60][1] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\line_cache[304][2] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(_01818_),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\line_cache[312][0] ),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_01888_),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\line_cache[237][3] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\line_cache[302][7] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(_01219_),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\line_cache[210][0] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_00984_),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\line_cache[18][6] ),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(_00798_),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\line_cache[217][1] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(_01041_),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\line_cache[160][2] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_00538_),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\line_cache[53][0] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_01807_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(\line_cache[272][5] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(_01533_),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(\line_cache[124][5] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(_00221_),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\line_cache[66][7] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(\line_cache[23][3] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(_01243_),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\line_cache[254][7] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(_01375_),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\line_cache[142][4] ),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\line_cache[227][0] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(_00380_),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\line_cache[59][2] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(_02194_),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\line_cache[92][1] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(_02489_),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\line_cache[207][4] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(_00956_),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\line_cache[269][2] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(_01498_),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\line_cache[116][0] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_01023_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_01128_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_00144_),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\line_cache[120][4] ),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(_00188_),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\line_cache[78][4] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(_02364_),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\line_cache[122][7] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(_00207_),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(\line_cache[184][1] ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(_00745_),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\line_cache[144][2] ),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\line_cache[225][6] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(_00394_),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\line_cache[275][5] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_01557_),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\line_cache[53][1] ),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(_02145_),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(\line_cache[94][3] ),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(\line_cache[250][5] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(_01341_),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(\line_cache[178][3] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\line_cache[265][1] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_01118_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(\line_cache[319][2] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\line_cache[301][1] ),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\line_cache[135][7] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(_00319_),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(\line_cache[121][1] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(_00193_),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\line_cache[146][6] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(_00414_),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\line_cache[91][0] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(_02480_),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\line_cache[239][2] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(\line_cache[53][2] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\line_cache[54][4] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(\line_cache[144][0] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(_00392_),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\line_cache[291][5] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(_01701_),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(\line_cache[222][7] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(_01095_),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(\line_cache[191][7] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(_00815_),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_01234_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(\line_cache[220][7] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(_01079_),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\line_cache[128][0] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(_00248_),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\line_cache[222][3] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(_01091_),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\line_cache[305][4] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\line_cache[187][3] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(\line_cache[190][0] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(_00800_),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\line_cache[292][1] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\line_cache[293][4] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\line_cache[167][6] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\line_cache[314][4] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(_01908_),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\line_cache[216][2] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(_01034_),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\line_cache[22][3] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(_01155_),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(\line_cache[160][5] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(_00541_),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_01705_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\line_cache[184][4] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(_00748_),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\line_cache[89][1] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(_02457_),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\line_cache[317][2] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\line_cache[233][1] ),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(_01185_),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\line_cache[138][6] ),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(_00342_),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\line_cache[165][6] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\line_cache[129][6] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_00582_),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\line_cache[93][3] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(_02499_),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\line_cache[207][7] ),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_00959_),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\line_cache[301][3] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\line_cache[29][2] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\line_cache[51][5] ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(_02133_),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\line_cache[313][3] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_00262_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(_01899_),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\line_cache[315][7] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(_01919_),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\line_cache[232][7] ),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(\line_cache[59][4] ),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(_02196_),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(\line_cache[218][4] ),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\line_cache[249][0] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\line_cache[67][3] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(_02267_),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\line_cache[314][0] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\line_cache[140][0] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(_00360_),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\line_cache[79][2] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\line_cache[105][6] ),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(_00054_),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\line_cache[248][1] ),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(_01313_),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\line_cache[61][0] ),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(_02216_),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\line_cache[268][0] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\line_cache[226][7] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_01904_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\line_cache[238][4] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(_01228_),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\line_cache[62][0] ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\line_cache[130][4] ),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(_00276_),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\line_cache[186][6] ),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(_00766_),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\line_cache[205][1] ),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(_00937_),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\line_cache[27][0] ),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\line_cache[133][1] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\line_cache[128][2] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(_00250_),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(\line_cache[251][3] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\line_cache[284][1] ),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(_01633_),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\line_cache[223][5] ),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(_01101_),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\line_cache[73][1] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(_02321_),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\line_cache[234][7] ),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_00297_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(_01199_),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\line_cache[274][5] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(\line_cache[158][6] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(_00518_),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\line_cache[74][7] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(_02335_),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\line_cache[266][3] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\line_cache[163][1] ),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\line_cache[254][6] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(_01374_),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\line_cache[212][4] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\line_cache[143][0] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\line_cache[16][0] ),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(_00616_),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\line_cache[85][2] ),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\line_cache[223][0] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(_01096_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\line_cache[295][5] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(_01733_),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(\line_cache[127][7] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(_00247_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_01004_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\line_cache[205][4] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(_00940_),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\line_cache[39][5] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(_02021_),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(\line_cache[120][2] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(_00186_),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(\line_cache[18][5] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(_00797_),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\line_cache[236][0] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(_01208_),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\line_cache[126][7] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(\line_cache[293][6] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(_01718_),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(\line_cache[298][0] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\line_cache[291][3] ),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(_01699_),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\line_cache[319][6] ),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\line_cache[216][5] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(_01037_),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\line_cache[163][7] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(_00567_),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_00239_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\line_cache[77][1] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(_02353_),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(\line_cache[307][6] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(\line_cache[156][0] ),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(_00496_),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\line_cache[285][3] ),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(_01643_),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\line_cache[245][1] ),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(\line_cache[123][3] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(_00211_),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\line_cache[267][3] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(\line_cache[30][4] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(_01868_),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(\line_cache[55][3] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(_02163_),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\line_cache[90][5] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\line_cache[219][6] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(\line_cache[274][7] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\line_cache[289][0] ),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\line_cache[313][1] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(_01897_),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_01483_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(\line_cache[305][6] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(_01830_),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(\line_cache[235][2] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\line_cache[181][0] ),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(\line_cache[207][0] ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\line_cache[299][7] ),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(_01767_),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\line_cache[14][3] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(_00443_),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\line_cache[280][0] ),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\line_cache[156][1] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(_01600_),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\line_cache[217][6] ),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(_01046_),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\line_cache[75][4] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(_02340_),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(\line_cache[57][6] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(_02182_),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\line_cache[59][3] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(_02195_),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\line_cache[191][4] ),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_01127_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_00497_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(\line_cache[72][2] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(_02314_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(\line_cache[98][6] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(_02542_),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(\line_cache[296][0] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(_01736_),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(\line_cache[15][1] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\line_cache[187][4] ),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(_00772_),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\line_cache[48][2] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\line_cache[228][4] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(_02098_),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\line_cache[117][1] ),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(_00153_),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\line_cache[127][1] ),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(\line_cache[69][6] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(_02286_),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(\line_cache[285][4] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(_01644_),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(\line_cache[237][6] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(_01222_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_01140_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(\line_cache[221][3] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(_01083_),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(\line_cache[94][5] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\line_cache[111][7] ),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(_00111_),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\line_cache[293][1] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(_01713_),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(\line_cache[105][2] ),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(\line_cache[296][4] ),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(_01740_),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\line_cache[159][1] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(\line_cache[95][4] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(_02516_),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(\line_cache[48][4] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(_02100_),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(\line_cache[61][3] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(\line_cache[198][6] ),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(_00870_),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\line_cache[53][6] ),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(_02150_),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\line_cache[185][3] ),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_00521_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(_00755_),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\line_cache[77][3] ),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(_02355_),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\line_cache[99][0] ),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(\line_cache[83][3] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(_02411_),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(\line_cache[85][1] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(_02425_),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(\line_cache[60][4] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\line_cache[182][4] ),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\line_cache[241][3] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(\line_cache[37][1] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(_02001_),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(\line_cache[197][3] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(_00859_),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(\line_cache[80][5] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(_02389_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(\line_cache[264][0] ),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(\line_cache[149][4] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(\line_cache[92][0] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(_02488_),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_01259_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(\line_cache[161][1] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(_00545_),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(\line_cache[295][4] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(_01732_),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(\line_cache[49][1] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(_02105_),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(\line_cache[233][6] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(_01190_),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(\line_cache[157][6] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(_00510_),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\line_cache[224][0] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(\line_cache[120][5] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(_00189_),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(\line_cache[22][0] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(\line_cache[79][4] ),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(_02372_),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(\line_cache[13][1] ),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(\line_cache[15][5] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(\line_cache[184][2] ),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(_00746_),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(\line_cache[117][3] ),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_01104_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(_00155_),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\line_cache[296][2] ),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(_01738_),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(\line_cache[295][7] ),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(_01735_),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(\line_cache[60][5] ),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(\line_cache[270][6] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(\line_cache[11][3] ),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(\line_cache[288][4] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(_01668_),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\line_cache[228][5] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(\line_cache[201][2] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(\line_cache[179][3] ),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(\line_cache[147][1] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(\line_cache[299][5] ),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(_01765_),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(\line_cache[284][0] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(_01632_),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(\line_cache[183][6] ),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(\line_cache[49][6] ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(_02110_),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\line_cache[229][2] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_01141_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(\line_cache[64][5] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(_02245_),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(\line_cache[231][1] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(\line_cache[159][4] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(_00524_),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(\line_cache[22][5] ),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(\line_cache[274][0] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(\line_cache[120][0] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(_00184_),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(\line_cache[292][0] ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\line_cache[89][3] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(_01704_),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(\line_cache[21][1] ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(_01065_),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(\line_cache[90][7] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(\line_cache[156][4] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(_00500_),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(\line_cache[95][6] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(\line_cache[208][2] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(_00962_),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(\line_cache[36][4] ),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_02459_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(_01996_),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(\line_cache[316][7] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(\line_cache[102][0] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(\line_cache[57][2] ),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(_02178_),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(\line_cache[140][4] ),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(_00364_),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(\line_cache[186][7] ),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(\line_cache[118][5] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(\line_cache[207][3] ),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\line_cache[71][1] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(_00955_),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(\line_cache[34][6] ),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(_01982_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(\line_cache[291][6] ),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(_01702_),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(\line_cache[202][5] ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(\line_cache[308][0] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(_01848_),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(\line_cache[15][2] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(\line_cache[250][3] ),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_02305_),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(\line_cache[141][6] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(_00374_),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(\line_cache[39][7] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(_02023_),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(\line_cache[31][6] ),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(\line_cache[308][2] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(_01850_),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(\line_cache[159][3] ),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(_00523_),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(\line_cache[147][4] ),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\line_cache[214][4] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(_00420_),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(\line_cache[58][4] ),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(\line_cache[68][1] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(\line_cache[48][1] ),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(\line_cache[299][1] ),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(\line_cache[145][0] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(\line_cache[118][6] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(_00166_),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(\line_cache[58][0] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(\line_cache[78][6] ),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_01020_),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(_02366_),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(\line_cache[290][7] ),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(\line_cache[181][3] ),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(\line_cache[92][2] ),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(_02490_),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(\line_cache[154][6] ),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(_00486_),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(\line_cache[236][4] ),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(_01212_),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(\line_cache[201][1] ),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\line_cache[227][3] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(_00905_),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(\line_cache[247][4] ),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(\line_cache[0][5] ),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(\line_cache[103][2] ),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(\line_cache[202][6] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(_00918_),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(\line_cache[268][4] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(\line_cache[309][3] ),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(_01859_),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(\line_cache[65][2] ),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_01131_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(\line_cache[56][4] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(_02172_),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(\line_cache[233][2] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(\line_cache[311][7] ),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(\line_cache[257][3] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(_01395_),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(\line_cache[215][1] ),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(\line_cache[225][1] ),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(_01113_),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(\line_cache[14][0] ),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\line_cache[252][1] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(\line_cache[198][7] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(\line_cache[119][0] ),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(_00168_),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(\line_cache[99][3] ),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(_02547_),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(\line_cache[318][3] ),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(\line_cache[56][0] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(_02168_),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(\line_cache[51][6] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(\line_cache[216][7] ),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_00236_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_01146_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_01353_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(\line_cache[21][3] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(_01067_),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(\line_cache[296][7] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(\line_cache[82][4] ),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(\line_cache[85][6] ),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(_02430_),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(\line_cache[309][1] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(\line_cache[183][7] ),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(_00743_),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(\line_cache[72][1] ),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\line_cache[0][0] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(\line_cache[83][0] ),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(\line_cache[90][3] ),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(\line_cache[305][1] ),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(_01825_),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(\line_cache[256][2] ),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(_01386_),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(\line_cache[101][0] ),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(\line_cache[251][6] ),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(\line_cache[319][1] ),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(\line_cache[95][5] ),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_00000_),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(_02517_),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(\line_cache[84][4] ),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(_02420_),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(\line_cache[93][1] ),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(_02497_),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(\line_cache[53][4] ),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(\line_cache[43][4] ),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(_02060_),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(\line_cache[179][7] ),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(\line_cache[265][3] ),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\line_cache[82][5] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(\line_cache[300][1] ),
    .X(net2436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(\line_cache[105][1] ),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(_00049_),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(\line_cache[141][1] ),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(_00369_),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(\line_cache[233][3] ),
    .X(net2441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(_01187_),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(\line_cache[95][3] ),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(_02515_),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(\line_cache[159][0] ),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_02405_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(\line_cache[22][6] ),
    .X(net2446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(_01158_),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(\line_cache[301][6] ),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(\line_cache[183][4] ),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(_00740_),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(\line_cache[209][1] ),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(_00969_),
    .X(net2452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(\line_cache[147][6] ),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(\line_cache[128][5] ),
    .X(net2454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2049 (.A(_00253_),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\line_cache[132][1] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2050 (.A(\line_cache[235][7] ),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2051 (.A(_01207_),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2052 (.A(\line_cache[223][2] ),
    .X(net2458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2053 (.A(\line_cache[197][1] ),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2054 (.A(_00857_),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2055 (.A(\line_cache[28][1] ),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2056 (.A(\line_cache[146][5] ),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2057 (.A(\line_cache[111][0] ),
    .X(net2463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2058 (.A(\line_cache[38][0] ),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2059 (.A(\line_cache[256][1] ),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_00289_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2060 (.A(\line_cache[248][2] ),
    .X(net2466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2061 (.A(\line_cache[107][0] ),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2062 (.A(\line_cache[253][4] ),
    .X(net2468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2063 (.A(\line_cache[146][3] ),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2064 (.A(\line_cache[118][4] ),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2065 (.A(\line_cache[207][1] ),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2066 (.A(\line_cache[181][6] ),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2067 (.A(\line_cache[207][2] ),
    .X(net2473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2068 (.A(\line_cache[288][2] ),
    .X(net2474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2069 (.A(_01666_),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\line_cache[31][2] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2070 (.A(\line_cache[253][6] ),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2071 (.A(\line_cache[223][7] ),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2072 (.A(_01103_),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2073 (.A(\line_cache[31][0] ),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2074 (.A(\line_cache[268][1] ),
    .X(net2480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2075 (.A(\line_cache[20][0] ),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2076 (.A(_00976_),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2077 (.A(\line_cache[129][3] ),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2078 (.A(_00259_),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2079 (.A(\line_cache[95][7] ),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_01954_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2080 (.A(_02519_),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2081 (.A(\line_cache[209][3] ),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2082 (.A(_00971_),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2083 (.A(\line_cache[202][7] ),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2084 (.A(\line_cache[143][1] ),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2085 (.A(\line_cache[57][3] ),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2086 (.A(_02179_),
    .X(net2492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2087 (.A(\line_cache[129][1] ),
    .X(net2493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2088 (.A(_00257_),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2089 (.A(\line_cache[127][0] ),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\line_cache[28][0] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2090 (.A(\line_cache[128][4] ),
    .X(net2496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2091 (.A(_00252_),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2092 (.A(\line_cache[252][5] ),
    .X(net2498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2093 (.A(\line_cache[269][1] ),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2094 (.A(\line_cache[16][5] ),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2095 (.A(_00621_),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2096 (.A(\line_cache[177][1] ),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2097 (.A(\line_cache[217][4] ),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2098 (.A(\line_cache[215][5] ),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2099 (.A(_01029_),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\line_cache[243][5] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_01680_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2100 (.A(\line_cache[101][2] ),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2101 (.A(\line_cache[180][0] ),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2102 (.A(_00712_),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2103 (.A(\line_cache[97][1] ),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2104 (.A(_02529_),
    .X(net2510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2105 (.A(\line_cache[140][5] ),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2106 (.A(_00365_),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2107 (.A(\line_cache[311][5] ),
    .X(net2513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2108 (.A(\line_cache[252][7] ),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2109 (.A(\line_cache[146][7] ),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\line_cache[12][4] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2110 (.A(\line_cache[317][6] ),
    .X(net2516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2111 (.A(_01934_),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2112 (.A(\line_cache[16][4] ),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2113 (.A(_00620_),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2114 (.A(\line_cache[219][7] ),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2115 (.A(_01063_),
    .X(net2521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2116 (.A(\line_cache[57][1] ),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2117 (.A(_02177_),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2118 (.A(\line_cache[251][2] ),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2119 (.A(\line_cache[151][7] ),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_00268_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2120 (.A(_00463_),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2121 (.A(\line_cache[92][5] ),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2122 (.A(_02493_),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2123 (.A(\line_cache[210][3] ),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2124 (.A(\line_cache[182][6] ),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2125 (.A(\line_cache[65][1] ),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2126 (.A(_02249_),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2127 (.A(\line_cache[75][0] ),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2128 (.A(\line_cache[305][3] ),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2129 (.A(_01827_),
    .X(net2535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\line_cache[229][3] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2130 (.A(\line_cache[26][4] ),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2131 (.A(\line_cache[285][2] ),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2132 (.A(\line_cache[286][5] ),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2133 (.A(\line_cache[285][0] ),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2134 (.A(\line_cache[76][1] ),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2135 (.A(\line_cache[190][6] ),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2136 (.A(\line_cache[151][5] ),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2137 (.A(_00461_),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2138 (.A(\line_cache[65][3] ),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2139 (.A(_02251_),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_01147_),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2140 (.A(\line_cache[252][0] ),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2141 (.A(\line_cache[0][3] ),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2142 (.A(_00003_),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2143 (.A(\line_cache[150][5] ),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2144 (.A(\line_cache[254][3] ),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2145 (.A(\line_cache[151][1] ),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2146 (.A(\line_cache[215][3] ),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2147 (.A(_01027_),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2148 (.A(\line_cache[186][5] ),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2149 (.A(\line_cache[151][3] ),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\line_cache[139][6] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2150 (.A(_00459_),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2151 (.A(\line_cache[141][3] ),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2152 (.A(_00371_),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2153 (.A(\line_cache[51][4] ),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2154 (.A(_02132_),
    .X(net2560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2155 (.A(\line_cache[191][6] ),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2156 (.A(\line_cache[49][2] ),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2157 (.A(\line_cache[27][4] ),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2158 (.A(_01596_),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2159 (.A(\line_cache[15][3] ),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_00350_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2160 (.A(\line_cache[253][1] ),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2161 (.A(\line_cache[119][7] ),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2162 (.A(_00175_),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2163 (.A(\line_cache[189][3] ),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2164 (.A(\line_cache[281][1] ),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2165 (.A(_01609_),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2166 (.A(\line_cache[23][5] ),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2167 (.A(_01245_),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2168 (.A(\line_cache[188][4] ),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2169 (.A(\line_cache[281][3] ),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\line_cache[3][7] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2170 (.A(_01611_),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2171 (.A(\line_cache[31][7] ),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2172 (.A(\line_cache[235][3] ),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2173 (.A(_01203_),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2174 (.A(\line_cache[273][3] ),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2175 (.A(_01539_),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2176 (.A(\line_cache[286][0] ),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2177 (.A(\line_cache[15][4] ),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2178 (.A(\line_cache[143][2] ),
    .X(net2584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2179 (.A(\line_cache[251][4] ),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_02031_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2180 (.A(\line_cache[196][2] ),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2181 (.A(_00850_),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2182 (.A(\line_cache[119][3] ),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2183 (.A(_00171_),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2184 (.A(\line_cache[75][3] ),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2185 (.A(_02339_),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2186 (.A(\line_cache[26][5] ),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2187 (.A(\line_cache[145][4] ),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2188 (.A(\line_cache[275][2] ),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2189 (.A(\line_cache[2][6] ),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\line_cache[105][0] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2190 (.A(\line_cache[150][3] ),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2191 (.A(\line_cache[280][4] ),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2192 (.A(_01604_),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2193 (.A(\line_cache[145][1] ),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2194 (.A(_00401_),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2195 (.A(\line_cache[31][5] ),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2196 (.A(\line_cache[32][2] ),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2197 (.A(_01962_),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2198 (.A(\line_cache[286][3] ),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2199 (.A(\line_cache[27][5] ),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_01277_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_00048_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2200 (.A(_01597_),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2201 (.A(\line_cache[268][2] ),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2202 (.A(\line_cache[72][4] ),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2203 (.A(_02316_),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2204 (.A(\line_cache[186][3] ),
    .X(net2610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2205 (.A(\line_cache[151][2] ),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2206 (.A(\line_cache[182][3] ),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2207 (.A(\line_cache[272][0] ),
    .X(net2613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2208 (.A(_01528_),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2209 (.A(\line_cache[286][4] ),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\line_cache[133][2] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2210 (.A(\line_cache[144][5] ),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2211 (.A(_00397_),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2212 (.A(\line_cache[264][7] ),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2213 (.A(\line_cache[284][2] ),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2214 (.A(_01634_),
    .X(net2620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2215 (.A(\line_cache[223][4] ),
    .X(net2621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2216 (.A(_01100_),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2217 (.A(\line_cache[15][7] ),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2218 (.A(\line_cache[272][4] ),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2219 (.A(_01532_),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_00298_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2220 (.A(\line_cache[74][5] ),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2221 (.A(\line_cache[270][0] ),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2222 (.A(\line_cache[8][2] ),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2223 (.A(\line_cache[252][4] ),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2224 (.A(\line_cache[96][2] ),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2225 (.A(_02522_),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2226 (.A(\line_cache[190][5] ),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2227 (.A(\line_cache[90][0] ),
    .X(net2633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2228 (.A(\line_cache[215][2] ),
    .X(net2634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2229 (.A(\line_cache[32][1] ),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\line_cache[135][4] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2230 (.A(\line_cache[273][6] ),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2231 (.A(_01542_),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2232 (.A(\line_cache[311][0] ),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2233 (.A(\line_cache[74][0] ),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2234 (.A(\line_cache[23][7] ),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2235 (.A(_01247_),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2236 (.A(\line_cache[271][3] ),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2237 (.A(\line_cache[73][0] ),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2238 (.A(\line_cache[180][2] ),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2239 (.A(_00714_),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_00316_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2240 (.A(\line_cache[200][5] ),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2241 (.A(_00901_),
    .X(net2647));
 sky130_fd_sc_hd__buf_1 hold2242 (.A(\pixel_double_counter[0] ),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2243 (.A(_02725_),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2244 (.A(\line_cache[63][3] ),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2245 (.A(\line_cache[40][1] ),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2246 (.A(\line_cache[63][2] ),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2247 (.A(\line_cache[63][0] ),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2248 (.A(\line_cache[271][1] ),
    .X(net2654));
 sky130_fd_sc_hd__buf_1 hold2249 (.A(\pixel_double_counter[1] ),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\line_cache[82][3] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2250 (.A(_02726_),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2251 (.A(\line_cache[271][4] ),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2252 (.A(\line_cache[65][6] ),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2253 (.A(_02254_),
    .X(net2659));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2254 (.A(\line_double_counter[1] ),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2255 (.A(_08502_),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2256 (.A(_02730_),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2257 (.A(\line_cache[199][3] ),
    .X(net2663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2258 (.A(_00875_),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2259 (.A(\line_cache[251][5] ),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_02403_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2260 (.A(\line_cache[271][2] ),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2261 (.A(\line_cache[273][2] ),
    .X(net2667));
 sky130_fd_sc_hd__buf_1 hold2262 (.A(\res_v_counter[6] ),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2263 (.A(_08447_),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2264 (.A(_02713_),
    .X(net2670));
 sky130_fd_sc_hd__buf_1 hold2265 (.A(net110),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2266 (.A(_02599_),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2267 (.A(net120),
    .X(net2673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2268 (.A(_02609_),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2269 (.A(\line_cache[172][6] ),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\line_cache[20][2] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2270 (.A(_00646_),
    .X(net2676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2271 (.A(\line_double_counter[2] ),
    .X(net2677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2272 (.A(_08506_),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2273 (.A(_02731_),
    .X(net2679));
 sky130_fd_sc_hd__buf_1 hold2274 (.A(\line_double_counter[3] ),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2275 (.A(_08508_),
    .X(net2681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2276 (.A(_02732_),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2277 (.A(\line_cache[108][6] ),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2278 (.A(_00078_),
    .X(net2684));
 sky130_fd_sc_hd__buf_1 hold2279 (.A(\res_v_counter[8] ),
    .X(net2685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_00978_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2280 (.A(_02715_),
    .X(net2686));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2281 (.A(\res_v_counter[9] ),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2282 (.A(_08469_),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2283 (.A(_02716_),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2284 (.A(\line_cache[175][0] ),
    .X(net2690));
 sky130_fd_sc_hd__clkbuf_2 hold2285 (.A(\res_v_counter[2] ),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2286 (.A(_08423_),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2287 (.A(_02709_),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2288 (.A(\line_cache[271][5] ),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2289 (.A(\prescaler_counter[8] ),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\line_cache[233][0] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2290 (.A(_04998_),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2291 (.A(_02568_),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2292 (.A(\line_cache[287][0] ),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2293 (.A(\line_cache[315][0] ),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2294 (.A(\line_cache[316][0] ),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2295 (.A(_01920_),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2296 (.A(\fb_read_state[0] ),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2297 (.A(_02569_),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2298 (.A(\line_cache[287][3] ),
    .X(net2704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2299 (.A(\line_cache[0][1] ),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\line_cache[226][3] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_01184_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2300 (.A(\line_cache[287][4] ),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2301 (.A(\line_cache[196][5] ),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2302 (.A(_00853_),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2303 (.A(\line_cache[27][1] ),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2304 (.A(\line_cache[27][2] ),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2305 (.A(\line_cache[287][5] ),
    .X(net2711));
 sky130_fd_sc_hd__buf_1 hold2306 (.A(\res_h_active[8] ),
    .X(net2712));
 sky130_fd_sc_hd__buf_2 hold2307 (.A(_08770_),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2308 (.A(_08804_),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2309 (.A(_02571_),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\line_cache[224][5] ),
    .X(net637));
 sky130_fd_sc_hd__buf_1 hold2310 (.A(net93),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2311 (.A(_02582_),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2312 (.A(\line_cache[154][0] ),
    .X(net2718));
 sky130_fd_sc_hd__buf_1 hold2313 (.A(net111),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2314 (.A(_02600_),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2315 (.A(\line_cache[287][2] ),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2316 (.A(\line_cache[252][2] ),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2317 (.A(\line_cache[255][3] ),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2318 (.A(\line_cache[191][0] ),
    .X(net2724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2319 (.A(\line_cache[253][3] ),
    .X(net2725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_01109_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2320 (.A(net104),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2321 (.A(_02593_),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2322 (.A(\base_v_fporch[0] ),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2323 (.A(\res_v_counter[7] ),
    .X(net2729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2324 (.A(_02714_),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2325 (.A(\res_v_active[5] ),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2326 (.A(\base_v_bporch[0] ),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2327 (.A(\base_h_bporch[0] ),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2328 (.A(net106),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2329 (.A(_02595_),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\line_cache[10][4] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2330 (.A(\line_cache[255][7] ),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2331 (.A(\base_v_fporch[2] ),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2332 (.A(\res_v_active[3] ),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2333 (.A(\base_v_sync[0] ),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2334 (.A(\line_cache[253][2] ),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2335 (.A(net95),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2336 (.A(_02584_),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2337 (.A(net101),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2338 (.A(_02590_),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2339 (.A(\res_v_active[2] ),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_00092_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2340 (.A(\line_cache[255][1] ),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2341 (.A(\line_cache[255][4] ),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2342 (.A(net99),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2343 (.A(_02588_),
    .X(net2749));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2344 (.A(\res_h_counter[6] ),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2345 (.A(_02703_),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2346 (.A(\line_cache[92][7] ),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2347 (.A(_03669_),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2348 (.A(\line_cache[127][4] ),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2349 (.A(_03175_),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\line_cache[175][6] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2350 (.A(_00244_),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2351 (.A(\res_v_active[6] ),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2352 (.A(\line_cache[222][0] ),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2353 (.A(_10708_),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2354 (.A(_01088_),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2355 (.A(\prescaler[3] ),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2356 (.A(\prescaler_counter[7] ),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2357 (.A(_04995_),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2358 (.A(_04997_),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2359 (.A(net108),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_00670_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2360 (.A(_02597_),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2361 (.A(\line_cache[255][2] ),
    .X(net2767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2362 (.A(\line_cache[260][4] ),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2363 (.A(\line_cache[212][3] ),
    .X(net2769));
 sky130_fd_sc_hd__buf_2 hold2364 (.A(\res_h_counter[0] ),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2365 (.A(_02697_),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2366 (.A(\res_v_active[4] ),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2367 (.A(\line_cache[12][1] ),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2368 (.A(\line_cache[213][6] ),
    .X(net2774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2369 (.A(\resolution[2] ),
    .X(net2775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\line_cache[267][2] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2370 (.A(\line_cache[225][7] ),
    .X(net2776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2371 (.A(\line_cache[192][5] ),
    .X(net2777));
 sky130_fd_sc_hd__buf_1 hold2372 (.A(\res_v_counter[1] ),
    .X(net2778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2373 (.A(_02708_),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2374 (.A(\line_cache[225][0] ),
    .X(net2780));
 sky130_fd_sc_hd__buf_2 hold2375 (.A(\line_cache_idx[3] ),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2376 (.A(_02575_),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2377 (.A(\line_cache[318][1] ),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2378 (.A(\line_cache[258][1] ),
    .X(net2784));
 sky130_fd_sc_hd__buf_1 hold2379 (.A(\res_h_counter[3] ),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_01482_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2380 (.A(_02700_),
    .X(net2786));
 sky130_fd_sc_hd__buf_4 hold2381 (.A(\line_cache_idx[5] ),
    .X(net2787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2382 (.A(_02577_),
    .X(net2788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2383 (.A(\line_cache[2][4] ),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2384 (.A(\line_cache[98][0] ),
    .X(net2790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2385 (.A(\line_cache[234][1] ),
    .X(net2791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2386 (.A(\line_cache[214][1] ),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2387 (.A(net100),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2388 (.A(_02589_),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2389 (.A(\line_cache[194][7] ),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\line_cache[229][6] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2390 (.A(\line_cache[35][0] ),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2391 (.A(\line_cache[319][3] ),
    .X(net2797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2392 (.A(\line_cache[3][0] ),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2393 (.A(\line_cache[132][7] ),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2394 (.A(_03104_),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2395 (.A(\line_cache[259][2] ),
    .X(net2801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2396 (.A(\line_cache[302][1] ),
    .X(net2802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2397 (.A(\line_cache[227][1] ),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2398 (.A(\line_cache[44][0] ),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2399 (.A(\line_cache[192][4] ),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_01123_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_01150_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2400 (.A(\line_cache[192][2] ),
    .X(net2806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2401 (.A(\line_cache[97][6] ),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2402 (.A(\line_cache[194][3] ),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2403 (.A(net102),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2404 (.A(_02591_),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2405 (.A(\line_cache[114][6] ),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2406 (.A(\base_h_fporch[4] ),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2407 (.A(\line_cache[226][6] ),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2408 (.A(\line_cache[302][2] ),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2409 (.A(\line_cache[192][0] ),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\line_cache[1][1] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2410 (.A(\line_cache[258][4] ),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2411 (.A(\line_cache[304][0] ),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2412 (.A(\line_cache[319][5] ),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2413 (.A(\line_cache[226][1] ),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2414 (.A(\line_cache[2][1] ),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2415 (.A(\line_cache[221][0] ),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2416 (.A(\line_cache[194][6] ),
    .X(net2822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2417 (.A(\line_cache[37][6] ),
    .X(net2823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2418 (.A(\line_cache[318][6] ),
    .X(net2824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2419 (.A(\line_cache[225][4] ),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_00889_),
    .X(net648));
 sky130_fd_sc_hd__buf_1 hold2420 (.A(\res_v_counter[3] ),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2421 (.A(_02710_),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2422 (.A(\line_cache[1][7] ),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2423 (.A(\line_cache[2][2] ),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2424 (.A(\line_cache[192][1] ),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2425 (.A(\line_cache[198][0] ),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2426 (.A(\line_cache[129][7] ),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2427 (.A(\line_cache[12][3] ),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2428 (.A(\line_cache[222][6] ),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2429 (.A(\line_cache[213][7] ),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\line_cache[69][3] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2430 (.A(\line_cache[193][6] ),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2431 (.A(\line_cache[192][3] ),
    .X(net2837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2432 (.A(\line_cache[65][5] ),
    .X(net2838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2433 (.A(net122),
    .X(net2839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2434 (.A(_07779_),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2435 (.A(_02611_),
    .X(net2841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2436 (.A(\line_cache[142][2] ),
    .X(net2842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2437 (.A(\line_cache[97][7] ),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2438 (.A(\line_cache[115][0] ),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2439 (.A(\line_cache[278][3] ),
    .X(net2845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_02283_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2440 (.A(\line_cache[93][7] ),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2441 (.A(\line_cache[194][4] ),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2442 (.A(\line_cache[263][6] ),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2443 (.A(\line_cache[115][7] ),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2444 (.A(\line_cache[278][4] ),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2445 (.A(\line_cache[190][7] ),
    .X(net2851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2446 (.A(\line_cache[93][6] ),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2447 (.A(\line_cache[25][3] ),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2448 (.A(\line_cache[193][0] ),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2449 (.A(\line_cache[194][5] ),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\line_cache[139][5] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2450 (.A(\line_cache[41][4] ),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2451 (.A(\line_cache[113][7] ),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2452 (.A(\line_cache[194][0] ),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2453 (.A(\line_cache[204][7] ),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2454 (.A(_10970_),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2455 (.A(\line_cache[46][3] ),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2456 (.A(\line_cache[67][5] ),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2457 (.A(\line_cache[193][4] ),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2458 (.A(\line_cache[41][3] ),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2459 (.A(\line_cache[317][1] ),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_00349_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2460 (.A(\line_cache[267][5] ),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2461 (.A(\line_cache[5][7] ),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2462 (.A(\line_cache[204][6] ),
    .X(net2868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2463 (.A(_10968_),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2464 (.A(\line_cache[83][4] ),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2465 (.A(\line_cache[141][5] ),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2466 (.A(\line_cache[140][2] ),
    .X(net2872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2467 (.A(\line_cache[6][7] ),
    .X(net2873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2468 (.A(\line_cache[229][7] ),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2469 (.A(\line_cache[261][6] ),
    .X(net2875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\line_cache[82][7] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2470 (.A(\line_cache[269][5] ),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2471 (.A(\line_cache[302][5] ),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2472 (.A(\line_cache[40][7] ),
    .X(net2878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2473 (.A(_04408_),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2474 (.A(\line_cache[212][5] ),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2475 (.A(\line_cache[35][3] ),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2476 (.A(\line_cache[47][4] ),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2477 (.A(\line_cache[213][3] ),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2478 (.A(\line_cache[319][4] ),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2479 (.A(\line_cache[270][2] ),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_02407_),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2480 (.A(\line_cache[218][2] ),
    .X(net2886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2481 (.A(net107),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2482 (.A(_02596_),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2483 (.A(\line_cache[193][1] ),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2484 (.A(\line_cache[183][0] ),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2485 (.A(\line_cache[263][5] ),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2486 (.A(\line_cache[113][6] ),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2487 (.A(_03374_),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2488 (.A(\line_cache[186][2] ),
    .X(net2894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2489 (.A(\line_cache[42][3] ),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\line_cache[37][2] ),
    .X(net655));
 sky130_fd_sc_hd__buf_1 hold2490 (.A(\base_h_counter[9] ),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2491 (.A(_02686_),
    .X(net2897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2492 (.A(\line_cache[263][2] ),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2493 (.A(\line_cache[176][4] ),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2494 (.A(\line_cache[1][6] ),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2495 (.A(\line_cache[283][6] ),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2496 (.A(\line_cache[269][3] ),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2497 (.A(\line_cache[259][7] ),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2498 (.A(\line_cache[234][2] ),
    .X(net2904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2499 (.A(\prescaler_counter[5] ),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\line_cache[197][0] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_02002_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2500 (.A(_04988_),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2501 (.A(_04989_),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2502 (.A(\line_cache[295][6] ),
    .X(net2908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2503 (.A(\line_cache[114][2] ),
    .X(net2909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2504 (.A(\line_cache[7][1] ),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2505 (.A(\line_cache[183][1] ),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2506 (.A(\line_cache[226][2] ),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2507 (.A(\line_cache[118][2] ),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2508 (.A(\line_cache[265][6] ),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2509 (.A(\line_cache[98][7] ),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\line_cache[298][7] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2510 (.A(\line_cache[24][3] ),
    .X(net2916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2511 (.A(\line_cache[1][0] ),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2512 (.A(\line_cache[274][2] ),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2513 (.A(\line_cache[24][1] ),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2514 (.A(\line_cache[294][2] ),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2515 (.A(\line_cache[119][4] ),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2516 (.A(\line_cache[224][3] ),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2517 (.A(\line_cache[132][6] ),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2518 (.A(_03102_),
    .X(net2924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2519 (.A(\line_cache[217][7] ),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_01759_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2520 (.A(\line_cache[9][4] ),
    .X(net2926));
 sky130_fd_sc_hd__buf_2 hold2521 (.A(\line_cache_idx[7] ),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2522 (.A(_02579_),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2523 (.A(\line_cache[2][5] ),
    .X(net2929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2524 (.A(\line_cache[39][4] ),
    .X(net2930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2525 (.A(\line_cache[274][1] ),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2526 (.A(\line_cache[7][0] ),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2527 (.A(\line_cache[260][1] ),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2528 (.A(\line_cache[32][4] ),
    .X(net2934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2529 (.A(\line_cache[182][2] ),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\line_cache[240][4] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2530 (.A(\line_cache[157][2] ),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2531 (.A(\line_cache[141][7] ),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2532 (.A(\line_cache[10][2] ),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2533 (.A(\line_cache[203][3] ),
    .X(net2939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2534 (.A(\line_cache[29][5] ),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2535 (.A(\line_cache[240][6] ),
    .X(net2941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2536 (.A(\line_cache[294][1] ),
    .X(net2942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2537 (.A(\line_cache[177][5] ),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2538 (.A(\line_cache[261][1] ),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2539 (.A(\line_cache[122][0] ),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_01252_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2540 (.A(\line_cache[41][2] ),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2541 (.A(\line_cache[244][7] ),
    .X(net2947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2542 (.A(\line_cache[38][1] ),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2543 (.A(\line_cache[114][4] ),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2544 (.A(\line_cache[30][2] ),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2545 (.A(\line_cache[304][4] ),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2546 (.A(\line_cache[225][5] ),
    .X(net2952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2547 (.A(\line_cache[17][6] ),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2548 (.A(\line_cache[276][3] ),
    .X(net2954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2549 (.A(\line_cache[43][1] ),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\line_cache[54][7] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2550 (.A(net105),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2551 (.A(_02594_),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2552 (.A(\res_v_counter[0] ),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2553 (.A(_02707_),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2554 (.A(\line_cache[195][6] ),
    .X(net2960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2555 (.A(\line_cache[303][3] ),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2556 (.A(\line_cache[185][7] ),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2557 (.A(\line_cache[262][6] ),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2558 (.A(\line_cache[115][4] ),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2559 (.A(\line_cache[46][2] ),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_02159_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2560 (.A(\line_cache[34][1] ),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2561 (.A(\line_cache[77][7] ),
    .X(net2967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2562 (.A(\line_cache[213][0] ),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2563 (.A(\line_cache[114][1] ),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2564 (.A(\line_cache[21][6] ),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2565 (.A(\line_cache[315][3] ),
    .X(net2971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2566 (.A(\line_cache[113][0] ),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2567 (.A(\line_cache[36][1] ),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2568 (.A(\line_cache[41][1] ),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2569 (.A(\line_cache[280][3] ),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\line_cache[137][3] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2570 (.A(\line_cache[314][1] ),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2571 (.A(\line_cache[279][6] ),
    .X(net2977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2572 (.A(\line_cache[63][7] ),
    .X(net2978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2573 (.A(\line_cache[49][7] ),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2574 (.A(\line_cache[19][1] ),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2575 (.A(\line_cache[98][3] ),
    .X(net2981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2576 (.A(\line_cache[273][4] ),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2577 (.A(\line_cache[317][5] ),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2578 (.A(\line_cache[217][5] ),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2579 (.A(\line_cache[265][2] ),
    .X(net2985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_00331_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2580 (.A(\line_cache[193][7] ),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2581 (.A(\line_cache[41][7] ),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2582 (.A(\line_cache[38][3] ),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2583 (.A(\line_cache[10][1] ),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2584 (.A(\line_cache[164][7] ),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2585 (.A(_11560_),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2586 (.A(\line_cache[113][5] ),
    .X(net2992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2587 (.A(\line_cache[46][0] ),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2588 (.A(\line_cache[179][5] ),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2589 (.A(\line_cache[6][6] ),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\line_cache[254][0] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2590 (.A(\line_cache[8][0] ),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2591 (.A(\line_cache[45][7] ),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2592 (.A(\line_cache[112][0] ),
    .X(net2998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2593 (.A(\resolution[3] ),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2594 (.A(\line_cache[240][7] ),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2595 (.A(\line_cache[282][6] ),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2596 (.A(\line_cache[7][5] ),
    .X(net3002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2597 (.A(\line_cache[121][3] ),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2598 (.A(\line_cache[46][4] ),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2599 (.A(\line_cache[197][2] ),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_00856_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_01368_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2600 (.A(\line_cache[258][6] ),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2601 (.A(\line_cache[20][5] ),
    .X(net3007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2602 (.A(\line_cache[228][2] ),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2603 (.A(\line_cache[51][1] ),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2604 (.A(\line_cache[44][3] ),
    .X(net3010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2605 (.A(\line_cache[112][1] ),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2606 (.A(\line_cache[305][2] ),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2607 (.A(\line_cache[161][0] ),
    .X(net3013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2608 (.A(\line_cache[140][3] ),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2609 (.A(\line_cache[98][5] ),
    .X(net3015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\line_cache[231][2] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2610 (.A(\line_cache[29][1] ),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2611 (.A(\line_cache[10][5] ),
    .X(net3017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2612 (.A(\res_v_counter[5] ),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2613 (.A(_02712_),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2614 (.A(\line_cache[273][5] ),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2615 (.A(\line_cache[248][7] ),
    .X(net3021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2616 (.A(\line_cache[284][3] ),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2617 (.A(\line_cache[257][6] ),
    .X(net3023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2618 (.A(\line_cache[114][7] ),
    .X(net3024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2619 (.A(\line_cache[61][2] ),
    .X(net3025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_01170_),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2620 (.A(\line_cache[263][0] ),
    .X(net3026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2621 (.A(\line_cache[262][2] ),
    .X(net3027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2622 (.A(\line_cache[47][5] ),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2623 (.A(\line_cache[23][4] ),
    .X(net3029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2624 (.A(\line_cache[262][4] ),
    .X(net3030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2625 (.A(\line_cache[66][6] ),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2626 (.A(\line_cache[66][2] ),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2627 (.A(\line_cache[219][3] ),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2628 (.A(\line_cache[319][7] ),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2629 (.A(\line_cache[5][1] ),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\line_cache[231][0] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2630 (.A(\line_cache[200][4] ),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2631 (.A(\line_cache[182][1] ),
    .X(net3037));
 sky130_fd_sc_hd__clkbuf_2 hold2632 (.A(\res_h_counter[1] ),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2633 (.A(_02698_),
    .X(net3039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2634 (.A(\line_cache[93][4] ),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2635 (.A(\line_cache[179][6] ),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2636 (.A(\line_cache[115][5] ),
    .X(net3042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2637 (.A(\line_cache[276][2] ),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2638 (.A(\line_cache[143][7] ),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2639 (.A(\line_cache[187][7] ),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_01168_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2640 (.A(\line_cache[34][2] ),
    .X(net3046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2641 (.A(\line_cache[277][4] ),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2642 (.A(\line_cache[121][7] ),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2643 (.A(\line_cache[290][4] ),
    .X(net3049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2644 (.A(\line_cache[35][6] ),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2645 (.A(\line_cache[42][4] ),
    .X(net3051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2646 (.A(\line_cache[131][4] ),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2647 (.A(\line_cache[261][2] ),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2648 (.A(\line_cache[50][6] ),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2649 (.A(\line_cache[118][1] ),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\line_cache[317][0] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2650 (.A(\line_cache[76][3] ),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2651 (.A(\line_cache[19][2] ),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2652 (.A(\line_cache[283][7] ),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2653 (.A(\line_cache[317][3] ),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2654 (.A(\line_cache[121][5] ),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2655 (.A(\line_cache[298][3] ),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2656 (.A(\line_cache[260][5] ),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2657 (.A(\line_cache[176][3] ),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2658 (.A(\line_cache[16][2] ),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2659 (.A(\line_cache[47][0] ),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_01928_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2660 (.A(\line_cache[64][3] ),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2661 (.A(\line_cache[57][5] ),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2662 (.A(\line_cache[220][6] ),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2663 (.A(\line_cache[29][3] ),
    .X(net3069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2664 (.A(\line_cache[77][5] ),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2665 (.A(\line_cache[46][5] ),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2666 (.A(\line_cache[141][2] ),
    .X(net3072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2667 (.A(\line_cache[213][4] ),
    .X(net3073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2668 (.A(\line_cache[308][3] ),
    .X(net3074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2669 (.A(\line_cache[4][1] ),
    .X(net3075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\line_cache[227][5] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2670 (.A(\line_cache[274][4] ),
    .X(net3076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2671 (.A(\line_cache[236][7] ),
    .X(net3077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2672 (.A(_10516_),
    .X(net3078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2673 (.A(\line_cache[301][7] ),
    .X(net3079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2674 (.A(\line_cache[178][2] ),
    .X(net3080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2675 (.A(\line_cache[210][2] ),
    .X(net3081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2676 (.A(\line_cache[29][7] ),
    .X(net3082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2677 (.A(\line_cache[115][6] ),
    .X(net3083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2678 (.A(\line_cache[79][7] ),
    .X(net3084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2679 (.A(\line_cache[117][5] ),
    .X(net3085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_01133_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2680 (.A(\line_cache[123][6] ),
    .X(net3086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2681 (.A(\line_cache[52][3] ),
    .X(net3087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2682 (.A(\line_cache[190][3] ),
    .X(net3088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2683 (.A(\line_cache[316][4] ),
    .X(net3089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2684 (.A(\line_cache[45][1] ),
    .X(net3090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2685 (.A(\line_cache[126][1] ),
    .X(net3091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2686 (.A(\line_cache[278][1] ),
    .X(net3092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2687 (.A(\line_cache[59][7] ),
    .X(net3093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2688 (.A(\line_cache[114][0] ),
    .X(net3094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2689 (.A(\line_cache[262][7] ),
    .X(net3095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\line_cache[68][0] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2690 (.A(\line_cache[273][0] ),
    .X(net3096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2691 (.A(\line_cache[262][0] ),
    .X(net3097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2692 (.A(\line_cache[48][3] ),
    .X(net3098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2693 (.A(\line_cache[116][3] ),
    .X(net3099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2694 (.A(\line_cache[279][4] ),
    .X(net3100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2695 (.A(\line_cache[47][1] ),
    .X(net3101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2696 (.A(\line_cache[269][7] ),
    .X(net3102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2697 (.A(\line_cache[282][2] ),
    .X(net3103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2698 (.A(\line_cache[49][5] ),
    .X(net3104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2699 (.A(\line_cache[33][7] ),
    .X(net3105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\line_cache[21][2] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_02272_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2700 (.A(\line_cache[143][5] ),
    .X(net3106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2701 (.A(\line_cache[76][6] ),
    .X(net3107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2702 (.A(_02350_),
    .X(net3108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2703 (.A(\line_cache[216][0] ),
    .X(net3109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2704 (.A(\line_cache[66][1] ),
    .X(net3110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2705 (.A(\line_cache[305][7] ),
    .X(net3111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2706 (.A(\line_cache[58][6] ),
    .X(net3112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2707 (.A(\line_cache[147][5] ),
    .X(net3113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2708 (.A(\line_cache[53][7] ),
    .X(net3114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2709 (.A(\line_cache[130][2] ),
    .X(net3115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\line_cache[20][4] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2710 (.A(\line_cache[161][3] ),
    .X(net3116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2711 (.A(\line_cache[214][2] ),
    .X(net3117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2712 (.A(\line_cache[218][1] ),
    .X(net3118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2713 (.A(\line_cache[6][5] ),
    .X(net3119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2714 (.A(\line_cache[213][5] ),
    .X(net3120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2715 (.A(\line_cache[248][6] ),
    .X(net3121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2716 (.A(\line_cache[282][1] ),
    .X(net3122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2717 (.A(\line_cache[275][6] ),
    .X(net3123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2718 (.A(\line_cache[261][7] ),
    .X(net3124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2719 (.A(\line_cache[285][7] ),
    .X(net3125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_00980_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2720 (.A(\line_cache[294][4] ),
    .X(net3126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2721 (.A(\line_cache[124][6] ),
    .X(net3127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2722 (.A(\line_cache[311][3] ),
    .X(net3128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2723 (.A(net96),
    .X(net3129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2724 (.A(_02585_),
    .X(net3130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2725 (.A(\line_cache[178][0] ),
    .X(net3131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2726 (.A(\line_cache[314][5] ),
    .X(net3132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2727 (.A(\line_cache[186][1] ),
    .X(net3133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2728 (.A(\line_cache[304][3] ),
    .X(net3134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2729 (.A(\line_cache[193][5] ),
    .X(net3135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\line_cache[137][0] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2730 (.A(\base_v_fporch[1] ),
    .X(net3136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2731 (.A(\line_cache[260][2] ),
    .X(net3137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2732 (.A(\line_cache[307][2] ),
    .X(net3138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2733 (.A(\line_cache[176][0] ),
    .X(net3139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2734 (.A(\line_cache[1][5] ),
    .X(net3140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2735 (.A(\line_cache[42][0] ),
    .X(net3141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2736 (.A(\line_cache[67][1] ),
    .X(net3142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2737 (.A(\line_cache[1][4] ),
    .X(net3143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2738 (.A(\line_cache[45][2] ),
    .X(net3144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2739 (.A(\line_cache[14][6] ),
    .X(net3145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_00328_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2740 (.A(\line_cache[9][5] ),
    .X(net3146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2741 (.A(\line_cache[62][1] ),
    .X(net3147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2742 (.A(\line_cache[244][6] ),
    .X(net3148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2743 (.A(\line_cache[217][2] ),
    .X(net3149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2744 (.A(\line_cache[46][1] ),
    .X(net3150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2745 (.A(\line_cache[78][3] ),
    .X(net3151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2746 (.A(\line_cache[84][6] ),
    .X(net3152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2747 (.A(\line_cache[43][2] ),
    .X(net3153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2748 (.A(\line_cache[33][2] ),
    .X(net3154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2749 (.A(\line_cache[4][2] ),
    .X(net3155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\line_cache[244][5] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2750 (.A(\line_cache[184][5] ),
    .X(net3156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2751 (.A(\line_cache[115][3] ),
    .X(net3157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2752 (.A(\line_cache[277][1] ),
    .X(net3158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2753 (.A(\line_cache[88][6] ),
    .X(net3159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2754 (.A(\line_cache[11][7] ),
    .X(net3160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2755 (.A(\line_cache[112][3] ),
    .X(net3161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2756 (.A(\line_cache[187][6] ),
    .X(net3162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2757 (.A(\line_cache[4][0] ),
    .X(net3163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2758 (.A(\line_cache[269][6] ),
    .X(net3164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2759 (.A(\line_cache[82][1] ),
    .X(net3165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_01285_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2760 (.A(\line_cache[215][0] ),
    .X(net3166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2761 (.A(\line_cache[5][6] ),
    .X(net3167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2762 (.A(\line_cache[266][0] ),
    .X(net3168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2763 (.A(\line_cache[317][7] ),
    .X(net3169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2764 (.A(\line_cache[188][6] ),
    .X(net3170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2765 (.A(\line_cache[181][4] ),
    .X(net3171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2766 (.A(\line_cache[233][7] ),
    .X(net3172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2767 (.A(\line_cache[258][2] ),
    .X(net3173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2768 (.A(\line_cache[209][4] ),
    .X(net3174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2769 (.A(\line_cache[46][7] ),
    .X(net3175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\line_cache[111][2] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2770 (.A(\line_cache[61][1] ),
    .X(net3176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2771 (.A(\line_cache[55][2] ),
    .X(net3177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2772 (.A(\line_cache[277][0] ),
    .X(net3178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2773 (.A(\line_cache[278][6] ),
    .X(net3179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2774 (.A(\line_cache[305][5] ),
    .X(net3180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2775 (.A(\line_cache[179][4] ),
    .X(net3181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2776 (.A(\line_cache[281][4] ),
    .X(net3182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2777 (.A(\line_cache[46][6] ),
    .X(net3183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2778 (.A(\line_cache[281][7] ),
    .X(net3184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2779 (.A(\line_cache[88][7] ),
    .X(net3185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_00106_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2780 (.A(\line_cache[61][5] ),
    .X(net3186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2781 (.A(\line_cache[65][7] ),
    .X(net3187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2782 (.A(net103),
    .X(net3188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2783 (.A(_02592_),
    .X(net3189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2784 (.A(\line_cache[283][2] ),
    .X(net3190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2785 (.A(\line_cache[270][7] ),
    .X(net3191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2786 (.A(\line_cache[307][7] ),
    .X(net3192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2787 (.A(\line_cache[143][4] ),
    .X(net3193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2788 (.A(\line_cache[309][6] ),
    .X(net3194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2789 (.A(\line_cache[59][5] ),
    .X(net3195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\line_cache[227][7] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2790 (.A(\line_cache[28][3] ),
    .X(net3196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2791 (.A(\line_cache[261][3] ),
    .X(net3197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2792 (.A(\line_cache[131][0] ),
    .X(net3198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2793 (.A(\line_cache[142][1] ),
    .X(net3199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2794 (.A(\line_cache[295][0] ),
    .X(net3200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2795 (.A(\line_cache[282][7] ),
    .X(net3201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2796 (.A(\line_cache[44][2] ),
    .X(net3202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2797 (.A(\line_cache[113][4] ),
    .X(net3203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2798 (.A(\line_cache[7][7] ),
    .X(net3204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2799 (.A(\line_cache[45][4] ),
    .X(net3205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_01066_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_01135_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2800 (.A(\base_v_sync[1] ),
    .X(net3206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2801 (.A(\line_cache[113][1] ),
    .X(net3207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2802 (.A(\line_cache[81][3] ),
    .X(net3208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2803 (.A(\line_cache[270][1] ),
    .X(net3209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2804 (.A(\line_cache[275][4] ),
    .X(net3210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2805 (.A(\line_cache[213][2] ),
    .X(net3211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2806 (.A(\line_cache[298][4] ),
    .X(net3212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2807 (.A(\line_cache[57][7] ),
    .X(net3213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2808 (.A(\line_cache[239][5] ),
    .X(net3214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2809 (.A(_01237_),
    .X(net3215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\line_cache[156][7] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2810 (.A(\line_cache[285][5] ),
    .X(net3216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2811 (.A(\line_cache[316][3] ),
    .X(net3217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2812 (.A(\line_cache[67][4] ),
    .X(net3218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2813 (.A(\line_cache[83][6] ),
    .X(net3219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2814 (.A(\line_cache[45][6] ),
    .X(net3220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2815 (.A(\line_cache[22][1] ),
    .X(net3221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2816 (.A(\line_cache[44][1] ),
    .X(net3222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2817 (.A(\line_cache[291][2] ),
    .X(net3223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2818 (.A(\line_cache[210][1] ),
    .X(net3224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2819 (.A(\line_cache[185][5] ),
    .X(net3225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_00503_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2820 (.A(\line_cache[227][2] ),
    .X(net3226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2821 (.A(\base_h_bporch[2] ),
    .X(net3227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2822 (.A(\line_cache[283][1] ),
    .X(net3228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2823 (.A(\line_cache[52][1] ),
    .X(net3229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2824 (.A(\line_cache[115][2] ),
    .X(net3230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2825 (.A(\line_cache[68][7] ),
    .X(net3231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2826 (.A(_04002_),
    .X(net3232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2827 (.A(\line_cache[12][6] ),
    .X(net3233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2828 (.A(\line_cache[152][6] ),
    .X(net3234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2829 (.A(\line_cache[192][6] ),
    .X(net3235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\line_cache[167][7] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2830 (.A(_00822_),
    .X(net3236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2831 (.A(\line_cache[5][2] ),
    .X(net3237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2832 (.A(\line_cache[163][3] ),
    .X(net3238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2833 (.A(\line_cache[20][6] ),
    .X(net3239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2834 (.A(\line_cache[48][0] ),
    .X(net3240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2835 (.A(\line_cache[98][2] ),
    .X(net3241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2836 (.A(\line_cache[176][1] ),
    .X(net3242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2837 (.A(\line_cache[130][3] ),
    .X(net3243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2838 (.A(\line_cache[94][7] ),
    .X(net3244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2839 (.A(\line_cache[261][5] ),
    .X(net3245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_00599_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2840 (.A(\line_cache[224][6] ),
    .X(net3246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2841 (.A(_01110_),
    .X(net3247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2842 (.A(\line_cache[17][1] ),
    .X(net3248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2843 (.A(\line_cache[51][7] ),
    .X(net3249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2844 (.A(\line_cache[82][2] ),
    .X(net3250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2845 (.A(\line_cache[192][7] ),
    .X(net3251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2846 (.A(_00823_),
    .X(net3252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2847 (.A(\line_cache[72][6] ),
    .X(net3253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2848 (.A(_03945_),
    .X(net3254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2849 (.A(\line_cache[5][4] ),
    .X(net3255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\line_cache[259][5] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2850 (.A(\line_cache[47][3] ),
    .X(net3256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2851 (.A(\line_cache[186][4] ),
    .X(net3257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2852 (.A(\line_cache[316][2] ),
    .X(net3258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2853 (.A(\line_cache[278][2] ),
    .X(net3259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2854 (.A(\line_cache[63][1] ),
    .X(net3260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2855 (.A(\line_cache[162][2] ),
    .X(net3261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2856 (.A(\line_cache[314][2] ),
    .X(net3262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2857 (.A(\line_cache[52][4] ),
    .X(net3263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2858 (.A(\line_cache[95][2] ),
    .X(net3264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2859 (.A(\line_cache[9][3] ),
    .X(net3265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_01413_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2860 (.A(\line_cache[283][3] ),
    .X(net3266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2861 (.A(\line_cache[19][6] ),
    .X(net3267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2862 (.A(\line_cache[5][0] ),
    .X(net3268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2863 (.A(\line_cache[56][2] ),
    .X(net3269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2864 (.A(\line_cache[131][2] ),
    .X(net3270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2865 (.A(\line_cache[80][4] ),
    .X(net3271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2866 (.A(\line_cache[262][5] ),
    .X(net3272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2867 (.A(\line_cache[193][3] ),
    .X(net3273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2868 (.A(\line_cache[65][0] ),
    .X(net3274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2869 (.A(\line_cache[313][4] ),
    .X(net3275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\line_cache[120][7] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2870 (.A(\line_cache[176][2] ),
    .X(net3276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2871 (.A(\line_cache[185][2] ),
    .X(net3277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2872 (.A(\line_cache[66][0] ),
    .X(net3278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2873 (.A(\line_cache[187][5] ),
    .X(net3279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2874 (.A(\line_cache[301][5] ),
    .X(net3280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2875 (.A(\base_h_bporch[1] ),
    .X(net3281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2876 (.A(\base_h_fporch[0] ),
    .X(net3282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2877 (.A(\line_cache[294][0] ),
    .X(net3283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2878 (.A(\line_cache[45][0] ),
    .X(net3284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2879 (.A(\line_cache[54][3] ),
    .X(net3285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_00191_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2880 (.A(\line_cache[147][3] ),
    .X(net3286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2881 (.A(\line_cache[62][2] ),
    .X(net3287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2882 (.A(\line_cache[279][5] ),
    .X(net3288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2883 (.A(\line_cache[34][4] ),
    .X(net3289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2884 (.A(\line_cache[181][1] ),
    .X(net3290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2885 (.A(\line_cache[184][0] ),
    .X(net3291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2886 (.A(\line_cache[179][1] ),
    .X(net3292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2887 (.A(\line_cache[291][4] ),
    .X(net3293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2888 (.A(\line_cache[118][0] ),
    .X(net3294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2889 (.A(\line_cache[47][2] ),
    .X(net3295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\line_cache[0][4] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2890 (.A(\line_cache[220][4] ),
    .X(net3296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2891 (.A(\line_cache[291][0] ),
    .X(net3297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2892 (.A(\line_cache[14][2] ),
    .X(net3298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2893 (.A(\line_cache[19][5] ),
    .X(net3299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2894 (.A(\line_cache[212][6] ),
    .X(net3300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2895 (.A(\line_cache[224][7] ),
    .X(net3301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2896 (.A(_01111_),
    .X(net3302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2897 (.A(\line_cache[307][0] ),
    .X(net3303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2898 (.A(\line_cache[116][2] ),
    .X(net3304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2899 (.A(\line_cache[104][6] ),
    .X(net3305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\line_cache[130][0] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_00004_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2900 (.A(_03502_),
    .X(net3306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2901 (.A(\line_cache[80][0] ),
    .X(net3307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2902 (.A(\line_cache[5][3] ),
    .X(net3308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2903 (.A(\line_cache[117][2] ),
    .X(net3309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2904 (.A(\line_cache[99][7] ),
    .X(net3310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2905 (.A(\line_cache[305][0] ),
    .X(net3311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2906 (.A(\line_cache[112][5] ),
    .X(net3312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2907 (.A(\line_cache[283][0] ),
    .X(net3313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2908 (.A(\line_cache[19][7] ),
    .X(net3314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2909 (.A(\line_cache[283][4] ),
    .X(net3315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\line_cache[315][2] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2910 (.A(\line_cache[117][7] ),
    .X(net3316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2911 (.A(\line_cache[4][3] ),
    .X(net3317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2912 (.A(\line_cache[197][5] ),
    .X(net3318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2913 (.A(\line_cache[184][3] ),
    .X(net3319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2914 (.A(\line_cache[113][3] ),
    .X(net3320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2915 (.A(\line_cache[193][2] ),
    .X(net3321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2916 (.A(\line_cache[54][0] ),
    .X(net3322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2917 (.A(\line_cache[178][1] ),
    .X(net3323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2918 (.A(\line_cache[257][7] ),
    .X(net3324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2919 (.A(\line_cache[198][1] ),
    .X(net3325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_01914_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2920 (.A(\base_v_bporch[1] ),
    .X(net3326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2921 (.A(\line_cache[99][6] ),
    .X(net3327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2922 (.A(\line_cache[291][1] ),
    .X(net3328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2923 (.A(\line_cache[112][2] ),
    .X(net3329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2924 (.A(\line_cache[10][3] ),
    .X(net3330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2925 (.A(\line_cache[261][4] ),
    .X(net3331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2926 (.A(\line_cache[157][5] ),
    .X(net3332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2927 (.A(\line_cache[42][2] ),
    .X(net3333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2928 (.A(\line_cache[19][3] ),
    .X(net3334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2929 (.A(\line_cache[209][5] ),
    .X(net3335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\line_cache[226][4] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2930 (.A(\line_cache[126][5] ),
    .X(net3336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2931 (.A(\line_cache[288][0] ),
    .X(net3337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2932 (.A(\line_cache[123][0] ),
    .X(net3338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2933 (.A(\line_cache[279][7] ),
    .X(net3339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2934 (.A(\line_cache[6][4] ),
    .X(net3340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2935 (.A(\line_cache[63][4] ),
    .X(net3341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2936 (.A(\line_cache[312][3] ),
    .X(net3342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2937 (.A(\line_cache[279][3] ),
    .X(net3343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2938 (.A(\line_cache[300][3] ),
    .X(net3344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2939 (.A(\line_cache[80][3] ),
    .X(net3345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_01124_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2940 (.A(\line_cache[162][1] ),
    .X(net3346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2941 (.A(\line_cache[278][5] ),
    .X(net3347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2942 (.A(\line_cache[4][4] ),
    .X(net3348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2943 (.A(\line_cache[258][7] ),
    .X(net3349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2944 (.A(\line_cache[81][5] ),
    .X(net3350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2945 (.A(\line_cache[11][5] ),
    .X(net3351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2946 (.A(\line_cache[125][7] ),
    .X(net3352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2947 (.A(\line_cache[143][3] ),
    .X(net3353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2948 (.A(\line_cache[14][1] ),
    .X(net3354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2949 (.A(\line_cache[296][3] ),
    .X(net3355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\line_cache[103][3] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2950 (.A(\line_cache[61][7] ),
    .X(net3356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2951 (.A(\line_cache[35][5] ),
    .X(net3357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2952 (.A(\line_cache[260][7] ),
    .X(net3358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2953 (.A(\line_cache[176][5] ),
    .X(net3359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2954 (.A(\line_cache[277][3] ),
    .X(net3360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2955 (.A(\line_cache[218][6] ),
    .X(net3361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2956 (.A(\line_cache[278][0] ),
    .X(net3362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2957 (.A(\line_cache[119][2] ),
    .X(net3363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2958 (.A(\line_cache[64][1] ),
    .X(net3364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2959 (.A(\line_cache[147][2] ),
    .X(net3365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_00035_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2960 (.A(\line_cache[94][2] ),
    .X(net3366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2961 (.A(\line_cache[277][2] ),
    .X(net3367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2962 (.A(\line_cache[64][0] ),
    .X(net3368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2963 (.A(\line_cache[306][2] ),
    .X(net3369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2964 (.A(\line_cache[44][4] ),
    .X(net3370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2965 (.A(\line_cache[41][0] ),
    .X(net3371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2966 (.A(\base_v_active[1] ),
    .X(net3372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2967 (.A(\line_cache[41][5] ),
    .X(net3373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2968 (.A(\line_cache[234][6] ),
    .X(net3374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2969 (.A(\line_cache[114][5] ),
    .X(net3375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\line_cache[203][1] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2970 (.A(\line_cache[129][4] ),
    .X(net3376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2971 (.A(\line_cache[54][2] ),
    .X(net3377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2972 (.A(\line_cache[300][0] ),
    .X(net3378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2973 (.A(\line_cache[30][7] ),
    .X(net3379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2974 (.A(\line_cache[47][7] ),
    .X(net3380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2975 (.A(\line_cache[178][6] ),
    .X(net3381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2976 (.A(\line_cache[157][3] ),
    .X(net3382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2977 (.A(\line_cache[195][1] ),
    .X(net3383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2978 (.A(\line_cache[30][1] ),
    .X(net3384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2979 (.A(\line_cache[142][0] ),
    .X(net3385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_00921_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2980 (.A(\line_cache[55][6] ),
    .X(net3386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2981 (.A(\line_cache[217][0] ),
    .X(net3387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2982 (.A(\line_cache[130][6] ),
    .X(net3388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2983 (.A(\line_cache[114][3] ),
    .X(net3389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2984 (.A(\line_cache[156][2] ),
    .X(net3390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2985 (.A(\line_cache[20][7] ),
    .X(net3391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2986 (.A(\line_cache[228][7] ),
    .X(net3392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2987 (.A(_01143_),
    .X(net3393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2988 (.A(\line_cache[181][5] ),
    .X(net3394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2989 (.A(\line_cache[160][0] ),
    .X(net3395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\line_cache[244][0] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2990 (.A(\line_cache[189][7] ),
    .X(net3396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2991 (.A(\line_cache[38][4] ),
    .X(net3397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2992 (.A(\line_cache[100][7] ),
    .X(net3398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2993 (.A(_03557_),
    .X(net3399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2994 (.A(\line_cache[260][6] ),
    .X(net3400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2995 (.A(\line_cache[289][1] ),
    .X(net3401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2996 (.A(\line_cache[50][2] ),
    .X(net3402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2997 (.A(\line_cache[315][1] ),
    .X(net3403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2998 (.A(\line_cache[297][5] ),
    .X(net3404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2999 (.A(\line_cache[209][2] ),
    .X(net3405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\line_cache[126][3] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00272_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_01280_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3000 (.A(\line_cache[276][4] ),
    .X(net3406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3001 (.A(\line_cache[80][2] ),
    .X(net3407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3002 (.A(\line_cache[239][3] ),
    .X(net3408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3003 (.A(\line_cache[97][5] ),
    .X(net3409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3004 (.A(\line_cache[50][0] ),
    .X(net3410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3005 (.A(\line_cache[118][7] ),
    .X(net3411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3006 (.A(\line_cache[261][0] ),
    .X(net3412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3007 (.A(\line_cache[84][7] ),
    .X(net3413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3008 (.A(\line_cache[309][7] ),
    .X(net3414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3009 (.A(\line_cache[68][6] ),
    .X(net3415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\line_cache[229][1] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3010 (.A(_04000_),
    .X(net3416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3011 (.A(\line_cache[197][6] ),
    .X(net3417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3012 (.A(\line_cache[315][5] ),
    .X(net3418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3013 (.A(\line_cache[64][2] ),
    .X(net3419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3014 (.A(\line_cache[52][0] ),
    .X(net3420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3015 (.A(\line_cache[180][3] ),
    .X(net3421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3016 (.A(\line_cache[187][2] ),
    .X(net3422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3017 (.A(\line_cache[216][3] ),
    .X(net3423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3018 (.A(\line_cache[58][3] ),
    .X(net3424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3019 (.A(\line_cache[301][4] ),
    .X(net3425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_01145_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3020 (.A(\line_cache[42][1] ),
    .X(net3426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3021 (.A(\line_cache[280][5] ),
    .X(net3427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3022 (.A(_01605_),
    .X(net3428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3023 (.A(\line_cache[123][7] ),
    .X(net3429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3024 (.A(\line_cache[33][5] ),
    .X(net3430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3025 (.A(\line_cache[272][1] ),
    .X(net3431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3026 (.A(\line_cache[264][6] ),
    .X(net3432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3027 (.A(\line_cache[94][1] ),
    .X(net3433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3028 (.A(\line_cache[235][4] ),
    .X(net3434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3029 (.A(\line_cache[304][5] ),
    .X(net3435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\line_cache[281][0] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3030 (.A(\prescaler_counter[0] ),
    .X(net3436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3031 (.A(\line_cache[96][3] ),
    .X(net3437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3032 (.A(\line_cache[45][3] ),
    .X(net3438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3033 (.A(\line_cache[77][4] ),
    .X(net3439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3034 (.A(\line_cache[147][0] ),
    .X(net3440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3035 (.A(\line_cache[143][6] ),
    .X(net3441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3036 (.A(\line_cache[131][6] ),
    .X(net3442));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3037 (.A(\base_h_counter[7] ),
    .X(net3443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3038 (.A(_02684_),
    .X(net3444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3039 (.A(\line_cache[161][5] ),
    .X(net3445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_01608_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3040 (.A(\line_cache[17][5] ),
    .X(net3446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3041 (.A(\line_cache[163][0] ),
    .X(net3447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3042 (.A(\line_cache[203][2] ),
    .X(net3448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3043 (.A(\line_cache[44][7] ),
    .X(net3449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3044 (.A(\line_cache[58][7] ),
    .X(net3450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3045 (.A(\line_cache[52][7] ),
    .X(net3451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3046 (.A(\line_cache[216][1] ),
    .X(net3452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3047 (.A(\line_cache[277][7] ),
    .X(net3453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3048 (.A(\line_cache[35][7] ),
    .X(net3454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3049 (.A(\line_cache[273][7] ),
    .X(net3455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\line_cache[164][5] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3050 (.A(\line_cache[56][3] ),
    .X(net3456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3051 (.A(\line_cache[51][3] ),
    .X(net3457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3052 (.A(\line_cache[157][1] ),
    .X(net3458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3053 (.A(\line_cache[19][4] ),
    .X(net3459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3054 (.A(\line_cache[9][0] ),
    .X(net3460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3055 (.A(\line_cache[117][4] ),
    .X(net3461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3056 (.A(\line_cache[129][2] ),
    .X(net3462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3057 (.A(\line_cache[163][4] ),
    .X(net3463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3058 (.A(\line_cache[201][6] ),
    .X(net3464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3059 (.A(\line_cache[196][1] ),
    .X(net3465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_00573_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3060 (.A(\line_cache[57][4] ),
    .X(net3466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3061 (.A(\line_cache[156][3] ),
    .X(net3467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3062 (.A(\line_cache[232][3] ),
    .X(net3468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3063 (.A(\line_cache[199][4] ),
    .X(net3469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3064 (.A(\line_cache[58][2] ),
    .X(net3470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3065 (.A(\line_cache[217][3] ),
    .X(net3471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3066 (.A(\line_cache[129][5] ),
    .X(net3472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3067 (.A(\line_cache[45][5] ),
    .X(net3473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3068 (.A(\line_cache[265][7] ),
    .X(net3474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3069 (.A(\line_cache[163][5] ),
    .X(net3475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\line_cache[218][0] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3070 (.A(\line_cache[232][4] ),
    .X(net3476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3071 (.A(\line_cache[276][1] ),
    .X(net3477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3072 (.A(\line_cache[298][2] ),
    .X(net3478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3073 (.A(\line_cache[177][7] ),
    .X(net3479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3074 (.A(\line_cache[113][2] ),
    .X(net3480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3075 (.A(\line_cache[131][5] ),
    .X(net3481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3076 (.A(\line_cache[33][6] ),
    .X(net3482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3077 (.A(\line_cache[262][3] ),
    .X(net3483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3078 (.A(\line_cache[290][2] ),
    .X(net3484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3079 (.A(\line_cache[260][0] ),
    .X(net3485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_01048_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3080 (.A(\line_cache[61][4] ),
    .X(net3486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3081 (.A(\line_cache[313][2] ),
    .X(net3487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3082 (.A(\line_cache[120][1] ),
    .X(net3488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3083 (.A(\line_cache[4][5] ),
    .X(net3489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3084 (.A(\line_cache[13][3] ),
    .X(net3490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3085 (.A(\line_cache[9][7] ),
    .X(net3491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3086 (.A(\line_cache[158][1] ),
    .X(net3492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3087 (.A(\line_cache[18][1] ),
    .X(net3493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3088 (.A(\line_cache[78][1] ),
    .X(net3494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3089 (.A(\line_cache[280][2] ),
    .X(net3495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\line_cache[167][5] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3090 (.A(_09848_),
    .X(net3496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3091 (.A(\line_cache[211][0] ),
    .X(net3497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3092 (.A(\line_cache[159][5] ),
    .X(net3498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3093 (.A(\line_cache[230][6] ),
    .X(net3499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3094 (.A(\line_cache[60][2] ),
    .X(net3500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3095 (.A(\line_cache[122][6] ),
    .X(net3501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3096 (.A(\res_v_active[0] ),
    .X(net3502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3097 (.A(\line_cache[33][4] ),
    .X(net3503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3098 (.A(\line_cache[49][0] ),
    .X(net3504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3099 (.A(\line_cache[270][5] ),
    .X(net3505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\line_cache[203][6] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_00597_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3100 (.A(\line_cache[195][0] ),
    .X(net3506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3101 (.A(\line_cache[279][0] ),
    .X(net3507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3102 (.A(\base_h_fporch[2] ),
    .X(net3508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3103 (.A(\line_cache[17][4] ),
    .X(net3509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3104 (.A(\line_cache[34][5] ),
    .X(net3510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3105 (.A(\line_cache[18][2] ),
    .X(net3511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3106 (.A(\line_cache[44][5] ),
    .X(net3512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3107 (.A(\line_cache[96][0] ),
    .X(net3513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3108 (.A(\line_cache[16][6] ),
    .X(net3514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3109 (.A(_00622_),
    .X(net3515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\line_cache[137][6] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3110 (.A(\line_cache[123][1] ),
    .X(net3516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3111 (.A(\res_v_counter[4] ),
    .X(net3517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3112 (.A(_02711_),
    .X(net3518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3113 (.A(\line_cache[58][1] ),
    .X(net3519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3114 (.A(\line_cache[269][0] ),
    .X(net3520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3115 (.A(\line_cache[47][6] ),
    .X(net3521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3116 (.A(\line_cache[32][3] ),
    .X(net3522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3117 (.A(\line_cache[195][5] ),
    .X(net3523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3118 (.A(\line_cache[266][1] ),
    .X(net3524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3119 (.A(\line_cache[131][7] ),
    .X(net3525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_00334_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3120 (.A(\line_cache[147][7] ),
    .X(net3526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3121 (.A(\res_v_active[1] ),
    .X(net3527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3122 (.A(\line_cache[306][1] ),
    .X(net3528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3123 (.A(\line_cache[292][6] ),
    .X(net3529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3124 (.A(\line_cache[17][2] ),
    .X(net3530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3125 (.A(\line_cache[157][4] ),
    .X(net3531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3126 (.A(\line_cache[257][4] ),
    .X(net3532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3127 (.A(\line_cache[235][5] ),
    .X(net3533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3128 (.A(\line_cache[23][6] ),
    .X(net3534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3129 (.A(\line_cache[33][1] ),
    .X(net3535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\line_cache[211][4] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3130 (.A(\line_cache[130][1] ),
    .X(net3536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3131 (.A(\line_cache[283][5] ),
    .X(net3537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3132 (.A(\line_cache[282][4] ),
    .X(net3538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3133 (.A(\line_cache[272][3] ),
    .X(net3539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3134 (.A(\line_cache[313][5] ),
    .X(net3540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3135 (.A(\line_cache[148][6] ),
    .X(net3541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3136 (.A(_02875_),
    .X(net3542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3137 (.A(\line_cache[300][4] ),
    .X(net3543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3138 (.A(\line_cache[5][5] ),
    .X(net3544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3139 (.A(\line_cache[136][6] ),
    .X(net3545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_00996_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3140 (.A(_03050_),
    .X(net3546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3141 (.A(\line_cache[212][7] ),
    .X(net3547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3142 (.A(\line_cache[96][5] ),
    .X(net3548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3143 (.A(\line_cache[288][6] ),
    .X(net3549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3144 (.A(_01670_),
    .X(net3550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3145 (.A(\line_cache[196][6] ),
    .X(net3551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3146 (.A(_00854_),
    .X(net3552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3147 (.A(\line_cache[77][0] ),
    .X(net3553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3148 (.A(\line_cache[60][6] ),
    .X(net3554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3149 (.A(\line_cache[50][1] ),
    .X(net3555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\line_cache[166][7] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3150 (.A(\line_cache[161][2] ),
    .X(net3556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3151 (.A(\line_cache[78][2] ),
    .X(net3557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3152 (.A(\line_cache[32][0] ),
    .X(net3558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3153 (.A(\line_cache[37][0] ),
    .X(net3559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3154 (.A(\line_cache[112][4] ),
    .X(net3560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3155 (.A(\line_cache[55][4] ),
    .X(net3561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3156 (.A(\line_cache[297][0] ),
    .X(net3562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3157 (.A(\line_cache[13][7] ),
    .X(net3563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3158 (.A(\line_cache[292][2] ),
    .X(net3564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3159 (.A(\line_cache[188][7] ),
    .X(net3565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_00591_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3160 (.A(\line_cache[52][5] ),
    .X(net3566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3161 (.A(\line_cache[300][5] ),
    .X(net3567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3162 (.A(\line_cache[164][6] ),
    .X(net3568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3163 (.A(_11558_),
    .X(net3569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3164 (.A(\line_cache[115][1] ),
    .X(net3570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3165 (.A(\line_cache[219][5] ),
    .X(net3571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3166 (.A(\line_cache[194][2] ),
    .X(net3572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3167 (.A(\line_cache[298][1] ),
    .X(net3573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3168 (.A(\line_cache[120][3] ),
    .X(net3574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3169 (.A(\line_cache[216][4] ),
    .X(net3575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\line_cache[100][0] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3170 (.A(\line_cache[35][4] ),
    .X(net3576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3171 (.A(\line_cache[116][7] ),
    .X(net3577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3172 (.A(\line_cache[208][3] ),
    .X(net3578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3173 (.A(\line_cache[63][5] ),
    .X(net3579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3174 (.A(\line_cache[288][7] ),
    .X(net3580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3175 (.A(_01671_),
    .X(net3581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3176 (.A(\line_cache[20][3] ),
    .X(net3582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3177 (.A(\line_cache[189][5] ),
    .X(net3583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3178 (.A(\line_cache[286][2] ),
    .X(net3584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3179 (.A(\line_cache[181][7] ),
    .X(net3585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_00008_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3180 (.A(\line_cache[158][2] ),
    .X(net3586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3181 (.A(\line_cache[24][6] ),
    .X(net3587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3182 (.A(_01334_),
    .X(net3588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3183 (.A(\line_cache[262][1] ),
    .X(net3589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3184 (.A(\line_cache[156][5] ),
    .X(net3590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3185 (.A(\line_cache[16][3] ),
    .X(net3591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3186 (.A(_04738_),
    .X(net3592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3187 (.A(\line_cache[195][3] ),
    .X(net3593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3188 (.A(\line_cache[272][2] ),
    .X(net3594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3189 (.A(\line_cache[208][1] ),
    .X(net3595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\line_cache[180][1] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3190 (.A(\line_cache[60][3] ),
    .X(net3596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3191 (.A(\line_cache[131][3] ),
    .X(net3597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3192 (.A(\line_cache[36][7] ),
    .X(net3598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3193 (.A(\line_cache[136][7] ),
    .X(net3599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3194 (.A(_03052_),
    .X(net3600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3195 (.A(\line_cache[276][7] ),
    .X(net3601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3196 (.A(\line_cache[194][1] ),
    .X(net3602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3197 (.A(\line_cache[22][2] ),
    .X(net3603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3198 (.A(\line_cache[195][4] ),
    .X(net3604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3199 (.A(\line_cache[81][7] ),
    .X(net3605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_00926_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_00713_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3200 (.A(\line_cache[198][2] ),
    .X(net3606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3201 (.A(\line_cache[6][3] ),
    .X(net3607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3202 (.A(\line_cache[187][1] ),
    .X(net3608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3203 (.A(\line_cache[300][6] ),
    .X(net3609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3204 (.A(\line_cache[284][6] ),
    .X(net3610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3205 (.A(\line_cache[128][6] ),
    .X(net3611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3206 (.A(\line_cache[310][6] ),
    .X(net3612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3207 (.A(\line_cache[279][2] ),
    .X(net3613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3208 (.A(\line_cache[294][6] ),
    .X(net3614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3209 (.A(\line_cache[253][5] ),
    .X(net3615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\line_cache[303][1] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3210 (.A(\line_cache[234][0] ),
    .X(net3616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3211 (.A(\line_cache[122][2] ),
    .X(net3617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3212 (.A(\line_cache[239][1] ),
    .X(net3618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3213 (.A(_01233_),
    .X(net3619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3214 (.A(\line_cache[28][6] ),
    .X(net3620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3215 (.A(\line_cache[100][6] ),
    .X(net3621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3216 (.A(_03555_),
    .X(net3622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3217 (.A(\line_cache[265][5] ),
    .X(net3623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3218 (.A(\line_cache[260][3] ),
    .X(net3624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3219 (.A(\line_cache[190][2] ),
    .X(net3625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_01809_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3220 (.A(\line_cache[316][5] ),
    .X(net3626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3221 (.A(_01925_),
    .X(net3627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3222 (.A(\line_cache[92][6] ),
    .X(net3628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3223 (.A(\line_cache[4][7] ),
    .X(net3629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3224 (.A(\line_cache[52][2] ),
    .X(net3630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3225 (.A(\line_cache[82][0] ),
    .X(net3631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3226 (.A(\line_cache[79][6] ),
    .X(net3632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3227 (.A(\resolution[1] ),
    .X(net3633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3228 (.A(\line_cache[160][3] ),
    .X(net3634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3229 (.A(\line_cache[98][1] ),
    .X(net3635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\line_cache[307][4] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3230 (.A(\line_cache[17][7] ),
    .X(net3636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3231 (.A(\line_cache[279][1] ),
    .X(net3637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3232 (.A(\line_cache[6][1] ),
    .X(net3638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3233 (.A(\line_cache[36][6] ),
    .X(net3639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3234 (.A(\line_cache[128][7] ),
    .X(net3640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3235 (.A(\line_cache[76][7] ),
    .X(net3641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3236 (.A(_02351_),
    .X(net3642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3237 (.A(\line_cache[21][5] ),
    .X(net3643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3238 (.A(\line_cache[310][1] ),
    .X(net3644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3239 (.A(\line_cache[233][5] ),
    .X(net3645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_01844_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3240 (.A(\line_cache[231][3] ),
    .X(net3646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3241 (.A(\line_cache[252][3] ),
    .X(net3647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3242 (.A(\line_cache[276][0] ),
    .X(net3648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3243 (.A(\line_cache[254][1] ),
    .X(net3649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3244 (.A(\line_cache[288][3] ),
    .X(net3650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3245 (.A(\line_cache[230][2] ),
    .X(net3651));
 sky130_fd_sc_hd__clkbuf_2 hold3246 (.A(\res_h_counter[7] ),
    .X(net3652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3247 (.A(_02704_),
    .X(net3653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3248 (.A(\line_cache[37][7] ),
    .X(net3654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3249 (.A(\line_cache[278][7] ),
    .X(net3655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\line_cache[161][4] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3250 (.A(\line_cache[239][0] ),
    .X(net3656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3251 (.A(_01232_),
    .X(net3657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3252 (.A(\line_cache[216][6] ),
    .X(net3658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3253 (.A(_01038_),
    .X(net3659));
 sky130_fd_sc_hd__buf_1 hold3254 (.A(\base_h_counter[4] ),
    .X(net3660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3255 (.A(_02681_),
    .X(net3661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3256 (.A(\line_cache[44][6] ),
    .X(net3662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3257 (.A(\line_cache[228][6] ),
    .X(net3663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3258 (.A(_01142_),
    .X(net3664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3259 (.A(\line_cache[292][4] ),
    .X(net3665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_00548_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3260 (.A(\line_cache[273][1] ),
    .X(net3666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3261 (.A(\line_cache[122][1] ),
    .X(net3667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3262 (.A(\line_cache[312][5] ),
    .X(net3668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3263 (.A(_01893_),
    .X(net3669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3264 (.A(\line_cache[304][6] ),
    .X(net3670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3265 (.A(_01822_),
    .X(net3671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3266 (.A(\line_cache[298][6] ),
    .X(net3672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3267 (.A(\line_cache[80][7] ),
    .X(net3673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3268 (.A(\line_cache[308][6] ),
    .X(net3674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3269 (.A(\line_cache[292][5] ),
    .X(net3675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\line_cache[244][4] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3270 (.A(\line_cache[265][4] ),
    .X(net3676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3271 (.A(\line_cache[285][1] ),
    .X(net3677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3272 (.A(\line_cache[272][7] ),
    .X(net3678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3273 (.A(_01535_),
    .X(net3679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3274 (.A(\line_cache[54][1] ),
    .X(net3680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3275 (.A(\line_cache[253][7] ),
    .X(net3681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3276 (.A(\line_cache[308][7] ),
    .X(net3682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3277 (.A(\line_cache[199][5] ),
    .X(net3683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3278 (.A(\line_cache[4][6] ),
    .X(net3684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3279 (.A(\line_cache[159][7] ),
    .X(net3685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_01284_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3280 (.A(\line_cache[34][7] ),
    .X(net3686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3281 (.A(\line_cache[200][3] ),
    .X(net3687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3282 (.A(\line_cache[37][5] ),
    .X(net3688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3283 (.A(\line_cache[24][2] ),
    .X(net3689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3284 (.A(\line_cache[183][3] ),
    .X(net3690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3285 (.A(\line_cache[21][0] ),
    .X(net3691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3286 (.A(\line_cache[276][5] ),
    .X(net3692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3287 (.A(\line_cache[146][2] ),
    .X(net3693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3288 (.A(\line_cache[196][7] ),
    .X(net3694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3289 (.A(_00855_),
    .X(net3695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\line_cache[122][3] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3290 (.A(\line_cache[312][1] ),
    .X(net3696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3291 (.A(\line_cache[201][5] ),
    .X(net3697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3292 (.A(\line_cache[43][3] ),
    .X(net3698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3293 (.A(\line_cache[236][6] ),
    .X(net3699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3294 (.A(_10514_),
    .X(net3700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3295 (.A(\line_cache[22][7] ),
    .X(net3701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3296 (.A(\line_cache[219][2] ),
    .X(net3702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3297 (.A(\line_cache[40][3] ),
    .X(net3703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3298 (.A(\line_cache[211][5] ),
    .X(net3704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3299 (.A(\line_cache[56][6] ),
    .X(net3705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\line_cache[228][1] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_00203_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3300 (.A(_02174_),
    .X(net3706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3301 (.A(\line_cache[254][2] ),
    .X(net3707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3302 (.A(\line_cache[257][5] ),
    .X(net3708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3303 (.A(\line_cache[296][5] ),
    .X(net3709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3304 (.A(_01741_),
    .X(net3710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3305 (.A(\line_cache[38][2] ),
    .X(net3711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3306 (.A(\line_cache[97][3] ),
    .X(net3712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3307 (.A(\line_cache[228][3] ),
    .X(net3713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3308 (.A(\line_cache[294][3] ),
    .X(net3714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3309 (.A(\line_cache[120][6] ),
    .X(net3715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\line_cache[227][4] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3310 (.A(\line_cache[280][6] ),
    .X(net3716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3311 (.A(_01606_),
    .X(net3717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3312 (.A(\line_cache[203][7] ),
    .X(net3718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3313 (.A(\line_cache[36][3] ),
    .X(net3719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3314 (.A(\line_cache[197][7] ),
    .X(net3720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3315 (.A(\line_cache[238][2] ),
    .X(net3721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3316 (.A(_01226_),
    .X(net3722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3317 (.A(\line_cache[316][6] ),
    .X(net3723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3318 (.A(_01926_),
    .X(net3724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3319 (.A(\line_cache[276][6] ),
    .X(net3725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_01132_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3320 (.A(\line_cache[176][6] ),
    .X(net3726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3321 (.A(\line_cache[275][3] ),
    .X(net3727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3322 (.A(\line_cache[188][1] ),
    .X(net3728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3323 (.A(\line_cache[30][6] ),
    .X(net3729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3324 (.A(\line_cache[163][2] ),
    .X(net3730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3325 (.A(\line_cache[266][2] ),
    .X(net3731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3326 (.A(\line_cache[56][7] ),
    .X(net3732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3327 (.A(_02175_),
    .X(net3733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3328 (.A(\line_cache[290][1] ),
    .X(net3734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3329 (.A(\base_h_sync[5] ),
    .X(net3735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\line_cache[306][4] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3330 (.A(\line_cache[203][5] ),
    .X(net3736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3331 (.A(\line_cache[124][3] ),
    .X(net3737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3332 (.A(\line_cache[52][6] ),
    .X(net3738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3333 (.A(\line_cache[209][7] ),
    .X(net3739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3334 (.A(\line_cache[292][3] ),
    .X(net3740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3335 (.A(\line_cache[201][3] ),
    .X(net3741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3336 (.A(\line_cache[128][3] ),
    .X(net3742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3337 (.A(\base_v_bporch[3] ),
    .X(net3743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3338 (.A(\line_cache[26][7] ),
    .X(net3744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3339 (.A(\line_cache[176][7] ),
    .X(net3745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_01836_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3340 (.A(\line_cache[309][5] ),
    .X(net3746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3341 (.A(\line_cache[311][6] ),
    .X(net3747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3342 (.A(\line_cache[48][7] ),
    .X(net3748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3343 (.A(_02103_),
    .X(net3749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3344 (.A(\line_cache[237][5] ),
    .X(net3750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3345 (.A(_01221_),
    .X(net3751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3346 (.A(\line_cache[210][6] ),
    .X(net3752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3347 (.A(\line_cache[196][3] ),
    .X(net3753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3348 (.A(\base_h_sync[0] ),
    .X(net3754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3349 (.A(\line_cache[201][7] ),
    .X(net3755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\line_cache[135][3] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3350 (.A(\line_cache[312][6] ),
    .X(net3756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3351 (.A(_01894_),
    .X(net3757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3352 (.A(\line_cache[313][7] ),
    .X(net3758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3353 (.A(\line_cache[53][5] ),
    .X(net3759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3354 (.A(\line_cache[200][6] ),
    .X(net3760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3355 (.A(_00902_),
    .X(net3761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3356 (.A(\line_cache[232][5] ),
    .X(net3762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3357 (.A(\line_cache[112][7] ),
    .X(net3763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3358 (.A(\line_cache[221][1] ),
    .X(net3764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3359 (.A(\line_cache[48][6] ),
    .X(net3765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_00315_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3360 (.A(_02102_),
    .X(net3766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3361 (.A(\line_cache[116][6] ),
    .X(net3767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3362 (.A(\line_cache[14][4] ),
    .X(net3768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3363 (.A(\line_cache[96][4] ),
    .X(net3769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3364 (.A(\line_cache[200][7] ),
    .X(net3770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3365 (.A(_00903_),
    .X(net3771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3366 (.A(\line_cache[195][2] ),
    .X(net3772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3367 (.A(\line_cache[67][2] ),
    .X(net3773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3368 (.A(\line_cache[26][0] ),
    .X(net3774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3369 (.A(\line_cache[286][1] ),
    .X(net3775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\line_cache[106][4] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3370 (.A(\line_cache[293][7] ),
    .X(net3776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3371 (.A(\line_cache[308][5] ),
    .X(net3777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3372 (.A(\line_cache[300][7] ),
    .X(net3778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3373 (.A(\line_cache[219][4] ),
    .X(net3779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3374 (.A(\line_cache[157][7] ),
    .X(net3780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3375 (.A(\line_cache[93][5] ),
    .X(net3781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3376 (.A(\line_cache[264][5] ),
    .X(net3782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3377 (.A(\base_h_bporch[3] ),
    .X(net3783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3378 (.A(\line_cache[64][6] ),
    .X(net3784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3379 (.A(_02246_),
    .X(net3785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_00060_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3380 (.A(\line_cache[78][7] ),
    .X(net3786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3381 (.A(\line_cache[182][5] ),
    .X(net3787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3382 (.A(\prescaler[0] ),
    .X(net3788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3383 (.A(\line_cache[24][5] ),
    .X(net3789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3384 (.A(_01333_),
    .X(net3790));
 sky130_fd_sc_hd__buf_4 hold3385 (.A(\line_cache_idx[4] ),
    .X(net3791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3386 (.A(_02576_),
    .X(net3792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3387 (.A(\line_cache[127][3] ),
    .X(net3793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3388 (.A(\line_cache[292][7] ),
    .X(net3794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3389 (.A(net97),
    .X(net3795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\line_cache[313][0] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3390 (.A(_07683_),
    .X(net3796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3391 (.A(_02586_),
    .X(net3797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3392 (.A(\line_cache[31][3] ),
    .X(net3798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3393 (.A(\line_cache[40][5] ),
    .X(net3799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3394 (.A(_02037_),
    .X(net3800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3395 (.A(\line_cache[13][5] ),
    .X(net3801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3396 (.A(\line_cache[145][5] ),
    .X(net3802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3397 (.A(\line_cache[289][7] ),
    .X(net3803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3398 (.A(\line_cache[24][7] ),
    .X(net3804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3399 (.A(_01335_),
    .X(net3805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_01137_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_01896_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3400 (.A(\line_cache[140][6] ),
    .X(net3806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3401 (.A(_00366_),
    .X(net3807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3402 (.A(\line_cache[296][6] ),
    .X(net3808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3403 (.A(_01742_),
    .X(net3809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3404 (.A(\line_cache[112][6] ),
    .X(net3810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3405 (.A(\line_cache[31][1] ),
    .X(net3811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3406 (.A(\line_cache[148][7] ),
    .X(net3812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3407 (.A(_02877_),
    .X(net3813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3408 (.A(\line_cache[64][7] ),
    .X(net3814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3409 (.A(\line_cache[304][7] ),
    .X(net3815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\line_cache[173][3] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3410 (.A(_01823_),
    .X(net3816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3411 (.A(\line_cache[63][6] ),
    .X(net3817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3412 (.A(\line_cache[80][6] ),
    .X(net3818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3413 (.A(\prescaler[2] ),
    .X(net3819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3414 (.A(\line_cache[272][6] ),
    .X(net3820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3415 (.A(_01534_),
    .X(net3821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3416 (.A(\base_v_active[6] ),
    .X(net3822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3417 (.A(\line_cache[32][6] ),
    .X(net3823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3418 (.A(_01966_),
    .X(net3824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3419 (.A(\line_cache[232][2] ),
    .X(net3825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_00651_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3420 (.A(\line_cache[7][6] ),
    .X(net3826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3421 (.A(\line_cache[222][1] ),
    .X(net3827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3422 (.A(\line_cache[195][7] ),
    .X(net3828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3423 (.A(\line_cache[32][7] ),
    .X(net3829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3424 (.A(_01967_),
    .X(net3830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3425 (.A(\line_cache[96][6] ),
    .X(net3831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3426 (.A(\line_cache[208][7] ),
    .X(net3832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3427 (.A(\line_cache[93][0] ),
    .X(net3833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3428 (.A(\line_cache[199][0] ),
    .X(net3834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3429 (.A(\line_cache[286][6] ),
    .X(net3835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\line_cache[139][1] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3430 (.A(\line_cache[25][7] ),
    .X(net3836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3431 (.A(\line_cache[145][6] ),
    .X(net3837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3432 (.A(\base_h_sync[6] ),
    .X(net3838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3433 (.A(\line_cache[156][6] ),
    .X(net3839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3434 (.A(_00502_),
    .X(net3840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3435 (.A(\line_cache[27][7] ),
    .X(net3841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3436 (.A(\line_cache[13][2] ),
    .X(net3842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3437 (.A(\line_cache[199][7] ),
    .X(net3843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3438 (.A(\line_cache[10][7] ),
    .X(net3844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3439 (.A(\line_cache[161][7] ),
    .X(net3845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_00345_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3440 (.A(\line_cache[6][2] ),
    .X(net3846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3441 (.A(\line_cache[56][5] ),
    .X(net3847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3442 (.A(_02173_),
    .X(net3848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3443 (.A(\line_cache[92][3] ),
    .X(net3849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3444 (.A(\line_cache[235][6] ),
    .X(net3850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3445 (.A(\line_cache[203][0] ),
    .X(net3851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3446 (.A(\line_cache[277][5] ),
    .X(net3852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3447 (.A(\line_cache[238][5] ),
    .X(net3853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3448 (.A(\line_cache[256][5] ),
    .X(net3854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3449 (.A(_01389_),
    .X(net3855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\line_cache[69][0] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3450 (.A(\line_cache[160][4] ),
    .X(net3856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3451 (.A(\line_cache[289][5] ),
    .X(net3857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3452 (.A(\line_cache[232][1] ),
    .X(net3858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3453 (.A(\line_cache[183][5] ),
    .X(net3859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3454 (.A(\line_cache[281][5] ),
    .X(net3860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3455 (.A(\line_cache[206][6] ),
    .X(net3861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3456 (.A(\line_cache[238][1] ),
    .X(net3862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3457 (.A(\line_cache[7][3] ),
    .X(net3863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3458 (.A(\line_cache[297][7] ),
    .X(net3864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3459 (.A(\line_cache[7][4] ),
    .X(net3865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_02280_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3460 (.A(\line_cache[215][6] ),
    .X(net3866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3461 (.A(\line_cache[293][5] ),
    .X(net3867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3462 (.A(\line_cache[102][1] ),
    .X(net3868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3463 (.A(\line_cache[268][5] ),
    .X(net3869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3464 (.A(\line_cache[219][0] ),
    .X(net3870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3465 (.A(\base_h_active[0] ),
    .X(net3871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3466 (.A(\line_cache[221][7] ),
    .X(net3872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3467 (.A(\line_cache[237][7] ),
    .X(net3873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3468 (.A(\line_cache[200][1] ),
    .X(net3874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3469 (.A(\line_cache[162][6] ),
    .X(net3875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\line_cache[111][1] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3470 (.A(\line_cache[220][1] ),
    .X(net3876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3471 (.A(\line_cache[169][4] ),
    .X(net3877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3472 (.A(\line_cache[237][1] ),
    .X(net3878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3473 (.A(\line_cache[229][5] ),
    .X(net3879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3474 (.A(\line_cache[302][0] ),
    .X(net3880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3475 (.A(\res_v_active[7] ),
    .X(net3881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3476 (.A(\line_cache[230][1] ),
    .X(net3882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3477 (.A(\line_cache[230][3] ),
    .X(net3883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3478 (.A(\line_cache[180][6] ),
    .X(net3884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3479 (.A(_00718_),
    .X(net3885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_00105_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3480 (.A(\line_cache[36][5] ),
    .X(net3886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3481 (.A(\line_cache[202][1] ),
    .X(net3887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3482 (.A(\line_cache[146][1] ),
    .X(net3888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3483 (.A(\line_cache[222][4] ),
    .X(net3889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3484 (.A(\line_cache[204][2] ),
    .X(net3890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3485 (.A(\line_cache[31][4] ),
    .X(net3891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3486 (.A(\line_cache[204][1] ),
    .X(net3892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3487 (.A(\line_cache[263][7] ),
    .X(net3893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3488 (.A(\line_cache[263][3] ),
    .X(net3894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3489 (.A(\line_cache[8][3] ),
    .X(net3895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\line_cache[149][3] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3490 (.A(\line_cache[309][0] ),
    .X(net3896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3491 (.A(\line_cache[144][1] ),
    .X(net3897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3492 (.A(\res_h_active[3] ),
    .X(net3898));
 sky130_fd_sc_hd__buf_2 hold3493 (.A(\line_cache_idx[6] ),
    .X(net3899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3494 (.A(_02578_),
    .X(net3900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3495 (.A(\line_cache[282][0] ),
    .X(net3901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3496 (.A(\line_cache[96][7] ),
    .X(net3902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3497 (.A(\line_cache[235][1] ),
    .X(net3903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3498 (.A(\line_cache[268][3] ),
    .X(net3904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3499 (.A(\line_cache[125][4] ),
    .X(net3905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\line_cache[258][3] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_00435_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3500 (.A(\line_cache[264][4] ),
    .X(net3906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3501 (.A(\line_cache[263][4] ),
    .X(net3907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3502 (.A(\line_cache[180][7] ),
    .X(net3908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3503 (.A(\line_cache[7][2] ),
    .X(net3909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3504 (.A(\prescaler[1] ),
    .X(net3910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3505 (.A(\base_v_active[2] ),
    .X(net3911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3506 (.A(\line_cache[155][7] ),
    .X(net3912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3507 (.A(\line_cache[244][1] ),
    .X(net3913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3508 (.A(\line_cache[87][5] ),
    .X(net3914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3509 (.A(\line_cache[25][5] ),
    .X(net3915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\line_cache[19][0] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3510 (.A(\line_cache[133][5] ),
    .X(net3916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3511 (.A(\base_h_active[7] ),
    .X(net3917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3512 (.A(\line_cache[263][1] ),
    .X(net3918));
 sky130_fd_sc_hd__buf_1 hold3513 (.A(\res_h_counter[2] ),
    .X(net3919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3514 (.A(_02699_),
    .X(net3920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3515 (.A(\line_cache[264][3] ),
    .X(net3921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3516 (.A(\base_h_bporch[6] ),
    .X(net3922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3517 (.A(\res_h_active[1] ),
    .X(net3923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3518 (.A(\line_cache[88][3] ),
    .X(net3924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3519 (.A(\line_cache[86][1] ),
    .X(net3925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_00880_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3520 (.A(\line_cache[87][1] ),
    .X(net3926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3521 (.A(\line_cache[102][5] ),
    .X(net3927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3522 (.A(\line_cache[255][6] ),
    .X(net3928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3523 (.A(\line_cache[8][4] ),
    .X(net3929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3524 (.A(\line_cache[241][7] ),
    .X(net3930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3525 (.A(\line_cache[124][1] ),
    .X(net3931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3526 (.A(\line_cache[170][2] ),
    .X(net3932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3527 (.A(\line_cache[277][6] ),
    .X(net3933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3528 (.A(\line_cache[74][4] ),
    .X(net3934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3529 (.A(\line_cache[184][6] ),
    .X(net3935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\line_cache[214][0] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3530 (.A(\line_cache[71][3] ),
    .X(net3936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3531 (.A(\base_v_active[4] ),
    .X(net3937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3532 (.A(\line_cache[70][4] ),
    .X(net3938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3533 (.A(\line_cache[264][1] ),
    .X(net3939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3534 (.A(\base_v_active[0] ),
    .X(net3940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3535 (.A(\line_cache[204][4] ),
    .X(net3941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3536 (.A(\base_v_active[8] ),
    .X(net3942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3537 (.A(\line_cache[75][5] ),
    .X(net3943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3538 (.A(\line_cache[237][4] ),
    .X(net3944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3539 (.A(\line_cache[168][1] ),
    .X(net3945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_01016_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3540 (.A(\line_cache[170][4] ),
    .X(net3946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3541 (.A(\line_cache[103][5] ),
    .X(net3947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3542 (.A(\line_cache[148][4] ),
    .X(net3948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3543 (.A(\line_cache[106][1] ),
    .X(net3949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3544 (.A(\line_cache[247][7] ),
    .X(net3950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3545 (.A(\line_cache[110][2] ),
    .X(net3951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3546 (.A(\line_cache[199][6] ),
    .X(net3952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3547 (.A(\line_cache[242][1] ),
    .X(net3953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3548 (.A(\line_cache[160][1] ),
    .X(net3954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3549 (.A(\line_cache[204][0] ),
    .X(net3955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\line_cache[219][1] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3550 (.A(\line_cache[168][0] ),
    .X(net3956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3551 (.A(\line_cache[252][6] ),
    .X(net3957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3552 (.A(_01358_),
    .X(net3958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3553 (.A(\line_cache[133][7] ),
    .X(net3959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3554 (.A(\line_cache[16][7] ),
    .X(net3960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3555 (.A(_00623_),
    .X(net3961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3556 (.A(\line_cache[104][2] ),
    .X(net3962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3557 (.A(\line_cache[243][3] ),
    .X(net3963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3558 (.A(\line_cache[74][1] ),
    .X(net3964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3559 (.A(\line_cache[248][5] ),
    .X(net3965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_01057_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3560 (.A(\base_h_bporch[5] ),
    .X(net3966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3561 (.A(\line_cache[171][3] ),
    .X(net3967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3562 (.A(\line_cache[168][3] ),
    .X(net3968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3563 (.A(\line_cache[101][5] ),
    .X(net3969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3564 (.A(\line_cache[230][7] ),
    .X(net3970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3565 (.A(\line_cache[139][0] ),
    .X(net3971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3566 (.A(\line_cache[105][7] ),
    .X(net3972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3567 (.A(\line_cache[75][1] ),
    .X(net3973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3568 (.A(\line_cache[104][3] ),
    .X(net3974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3569 (.A(\line_cache[169][5] ),
    .X(net3975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\line_cache[103][4] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3570 (.A(\line_cache[169][7] ),
    .X(net3976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3571 (.A(\line_cache[170][6] ),
    .X(net3977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3572 (.A(\line_cache[75][2] ),
    .X(net3978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3573 (.A(\line_cache[243][0] ),
    .X(net3979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3574 (.A(\line_cache[204][5] ),
    .X(net3980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3575 (.A(\line_cache[169][3] ),
    .X(net3981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3576 (.A(\line_cache[173][7] ),
    .X(net3982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3577 (.A(\line_cache[172][3] ),
    .X(net3983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3578 (.A(\line_cache[138][2] ),
    .X(net3984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3579 (.A(\line_cache[71][0] ),
    .X(net3985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_00036_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3580 (.A(\line_cache[6][0] ),
    .X(net3986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3581 (.A(\line_cache[86][4] ),
    .X(net3987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3582 (.A(\line_cache[220][3] ),
    .X(net3988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3583 (.A(\line_cache[204][3] ),
    .X(net3989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3584 (.A(\line_cache[148][3] ),
    .X(net3990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3585 (.A(\line_cache[242][6] ),
    .X(net3991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3586 (.A(\line_cache[245][0] ),
    .X(net3992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3587 (.A(\line_cache[169][2] ),
    .X(net3993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3588 (.A(\line_cache[205][6] ),
    .X(net3994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3589 (.A(\line_cache[40][6] ),
    .X(net3995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\line_cache[3][1] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3590 (.A(_02038_),
    .X(net3996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3591 (.A(\line_cache[109][4] ),
    .X(net3997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3592 (.A(\line_cache[87][2] ),
    .X(net3998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3593 (.A(\line_cache[136][0] ),
    .X(net3999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3594 (.A(\line_cache[154][3] ),
    .X(net4000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3595 (.A(\line_cache[109][0] ),
    .X(net4001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3596 (.A(\line_cache[171][6] ),
    .X(net4002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3597 (.A(\line_cache[107][7] ),
    .X(net4003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3598 (.A(\line_cache[223][3] ),
    .X(net4004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3599 (.A(\line_cache[111][4] ),
    .X(net4005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_01403_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_02025_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3600 (.A(\line_cache[106][2] ),
    .X(net4006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3601 (.A(\base_h_fporch[1] ),
    .X(net4007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3602 (.A(\line_cache[268][6] ),
    .X(net4008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3603 (.A(_01494_),
    .X(net4009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3604 (.A(\line_cache[132][3] ),
    .X(net4010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3605 (.A(\line_cache[166][0] ),
    .X(net4011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3606 (.A(\line_cache[167][3] ),
    .X(net4012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3607 (.A(\line_cache[170][3] ),
    .X(net4013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3608 (.A(\line_cache[105][3] ),
    .X(net4014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3609 (.A(\line_cache[190][1] ),
    .X(net4015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\line_cache[78][0] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3610 (.A(\line_cache[208][6] ),
    .X(net4016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3611 (.A(\line_cache[8][6] ),
    .X(net4017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3612 (.A(_02470_),
    .X(net4018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3613 (.A(\line_cache[91][2] ),
    .X(net4019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3614 (.A(\line_cache[169][1] ),
    .X(net4020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3615 (.A(\line_cache[170][1] ),
    .X(net4021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3616 (.A(\line_cache[189][4] ),
    .X(net4022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3617 (.A(\line_cache[232][6] ),
    .X(net4023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3618 (.A(\line_cache[85][7] ),
    .X(net4024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3619 (.A(\line_cache[240][3] ),
    .X(net4025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_02360_),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3620 (.A(\res_h_active[0] ),
    .X(net4026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3621 (.A(\line_cache[150][0] ),
    .X(net4027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3622 (.A(\line_cache[242][3] ),
    .X(net4028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3623 (.A(\line_cache[73][4] ),
    .X(net4029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3624 (.A(\line_cache[86][2] ),
    .X(net4030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3625 (.A(\line_cache[89][5] ),
    .X(net4031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3626 (.A(\line_cache[242][2] ),
    .X(net4032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3627 (.A(\line_cache[152][5] ),
    .X(net4033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3628 (.A(\line_cache[166][4] ),
    .X(net4034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3629 (.A(\line_cache[165][1] ),
    .X(net4035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\line_cache[101][3] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3630 (.A(\line_cache[88][0] ),
    .X(net4036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3631 (.A(\base_h_active[4] ),
    .X(net4037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3632 (.A(\line_cache[160][6] ),
    .X(net4038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3633 (.A(_00542_),
    .X(net4039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3634 (.A(\line_cache[86][6] ),
    .X(net4040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3635 (.A(\line_cache[171][0] ),
    .X(net4041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3636 (.A(\line_cache[109][2] ),
    .X(net4042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3637 (.A(\line_cache[164][1] ),
    .X(net4043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3638 (.A(\line_cache[109][1] ),
    .X(net4044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3639 (.A(\line_cache[170][7] ),
    .X(net4045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_00019_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3640 (.A(\line_cache[68][2] ),
    .X(net4046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3641 (.A(\line_cache[231][7] ),
    .X(net4047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3642 (.A(\base_h_sync[4] ),
    .X(net4048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3643 (.A(\line_cache[166][1] ),
    .X(net4049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3644 (.A(\line_cache[134][1] ),
    .X(net4050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3645 (.A(\line_cache[232][0] ),
    .X(net4051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3646 (.A(\line_cache[70][1] ),
    .X(net4052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3647 (.A(\line_cache[106][7] ),
    .X(net4053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3648 (.A(\line_cache[138][1] ),
    .X(net4054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3649 (.A(\line_cache[144][7] ),
    .X(net4055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\line_cache[259][3] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3650 (.A(\line_cache[145][7] ),
    .X(net4056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3651 (.A(\line_cache[87][4] ),
    .X(net4057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3652 (.A(\line_double_counter[0] ),
    .X(net4058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3653 (.A(\line_cache[109][7] ),
    .X(net4059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3654 (.A(\line_cache[154][2] ),
    .X(net4060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3655 (.A(\line_cache[144][4] ),
    .X(net4061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3656 (.A(\base_h_sync[1] ),
    .X(net4062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3657 (.A(\res_h_active[7] ),
    .X(net4063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3658 (.A(\line_cache[74][6] ),
    .X(net4064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3659 (.A(\line_cache[171][2] ),
    .X(net4065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_01411_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3660 (.A(\line_cache[110][1] ),
    .X(net4066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3661 (.A(\base_v_sync[2] ),
    .X(net4067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3662 (.A(\line_cache[69][1] ),
    .X(net4068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3663 (.A(\line_cache[107][3] ),
    .X(net4069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3664 (.A(\line_cache[160][7] ),
    .X(net4070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3665 (.A(\line_cache[154][1] ),
    .X(net4071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3666 (.A(\line_cache[151][6] ),
    .X(net4072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3667 (.A(\line_cache[100][5] ),
    .X(net4073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3668 (.A(\line_cache[108][2] ),
    .X(net4074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3669 (.A(\line_cache[84][2] ),
    .X(net4075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\line_cache[67][0] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3670 (.A(\line_cache[153][3] ),
    .X(net4076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3671 (.A(\line_cache[166][6] ),
    .X(net4077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3672 (.A(\line_cache[173][5] ),
    .X(net4078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3673 (.A(\line_cache[171][4] ),
    .X(net4079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3674 (.A(\line_cache[188][3] ),
    .X(net4080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3675 (.A(\line_cache[84][3] ),
    .X(net4081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3676 (.A(\line_cache[275][7] ),
    .X(net4082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3677 (.A(\line_cache[69][5] ),
    .X(net4083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3678 (.A(\line_cache[68][4] ),
    .X(net4084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3679 (.A(\line_cache[85][5] ),
    .X(net4085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_02264_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3680 (.A(\res_h_active[2] ),
    .X(net4086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3681 (.A(\line_cache[134][2] ),
    .X(net4087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3682 (.A(\line_cache[101][7] ),
    .X(net4088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3683 (.A(\line_cache[152][3] ),
    .X(net4089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3684 (.A(\line_cache[70][2] ),
    .X(net4090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3685 (.A(\line_cache[171][1] ),
    .X(net4091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3686 (.A(\line_cache[168][5] ),
    .X(net4092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3687 (.A(\line_cache[72][0] ),
    .X(net4093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3688 (.A(\line_cache[153][7] ),
    .X(net4094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3689 (.A(\line_cache[165][0] ),
    .X(net4095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\line_cache[230][5] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3690 (.A(\line_cache[191][1] ),
    .X(net4096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3691 (.A(\line_cache[191][5] ),
    .X(net4097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3692 (.A(\line_cache[286][7] ),
    .X(net4098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3693 (.A(\line_cache[174][2] ),
    .X(net4099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3694 (.A(\line_cache[87][3] ),
    .X(net4100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3695 (.A(\line_cache[155][0] ),
    .X(net4101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3696 (.A(\line_cache[68][5] ),
    .X(net4102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3697 (.A(\line_cache[166][2] ),
    .X(net4103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3698 (.A(\line_cache[89][7] ),
    .X(net4104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3699 (.A(\line_cache[8][5] ),
    .X(net4105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\line_cache[2][0] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_01165_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3700 (.A(_02469_),
    .X(net4106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3701 (.A(\line_cache[90][2] ),
    .X(net4107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3702 (.A(\line_cache[149][6] ),
    .X(net4108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3703 (.A(\line_cache[247][5] ),
    .X(net4109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3704 (.A(\line_cache[168][2] ),
    .X(net4110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3705 (.A(\line_cache[148][5] ),
    .X(net4111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3706 (.A(\line_cache[256][7] ),
    .X(net4112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3707 (.A(_01391_),
    .X(net4113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3708 (.A(\line_cache[148][2] ),
    .X(net4114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3709 (.A(\line_cache[205][0] ),
    .X(net4115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\line_cache[37][4] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3710 (.A(\line_cache[236][3] ),
    .X(net4116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3711 (.A(\line_cache[256][3] ),
    .X(net4117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3712 (.A(\line_cache[207][6] ),
    .X(net4118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3713 (.A(\line_cache[256][6] ),
    .X(net4119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3714 (.A(_01390_),
    .X(net4120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3715 (.A(\line_cache[70][0] ),
    .X(net4121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3716 (.A(\line_cache[134][6] ),
    .X(net4122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3717 (.A(\line_cache[137][7] ),
    .X(net4123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3718 (.A(\res_h_active[5] ),
    .X(net4124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3719 (.A(\line_cache[137][5] ),
    .X(net4125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_02004_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3720 (.A(\line_cache[73][2] ),
    .X(net4126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3721 (.A(\line_cache[250][2] ),
    .X(net4127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3722 (.A(\line_cache[154][7] ),
    .X(net4128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3723 (.A(\line_cache[249][5] ),
    .X(net4129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3724 (.A(\line_cache[134][3] ),
    .X(net4130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3725 (.A(\line_cache[244][3] ),
    .X(net4131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3726 (.A(\line_cache[248][0] ),
    .X(net4132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3727 (.A(\line_cache[125][5] ),
    .X(net4133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3728 (.A(\line_cache[136][4] ),
    .X(net4134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3729 (.A(\line_cache[87][7] ),
    .X(net4135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\line_cache[318][4] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3730 (.A(\line_cache[310][2] ),
    .X(net4136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3731 (.A(\base_h_sync[2] ),
    .X(net4137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3732 (.A(\line_cache[164][3] ),
    .X(net4138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3733 (.A(\line_cache[169][6] ),
    .X(net4139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3734 (.A(\line_cache[101][1] ),
    .X(net4140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3735 (.A(\line_cache[164][4] ),
    .X(net4141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3736 (.A(\line_cache[241][5] ),
    .X(net4142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3737 (.A(\line_cache[248][4] ),
    .X(net4143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3738 (.A(\line_cache[206][2] ),
    .X(net4144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3739 (.A(\res_h_active[6] ),
    .X(net4145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_01940_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3740 (.A(\line_cache[135][5] ),
    .X(net4146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3741 (.A(\line_cache[152][0] ),
    .X(net4147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3742 (.A(\line_cache[175][2] ),
    .X(net4148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3743 (.A(\line_cache[73][5] ),
    .X(net4149));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3744 (.A(\base_h_counter[8] ),
    .X(net4150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3745 (.A(_08077_),
    .X(net4151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3746 (.A(_02685_),
    .X(net4152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3747 (.A(\line_cache[241][2] ),
    .X(net4153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3748 (.A(\line_cache[250][0] ),
    .X(net4154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3749 (.A(\line_cache[89][2] ),
    .X(net4155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\line_cache[71][4] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3750 (.A(\line_cache[153][5] ),
    .X(net4156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3751 (.A(\base_v_active[5] ),
    .X(net4157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3752 (.A(\line_cache[138][5] ),
    .X(net4158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3753 (.A(\line_cache[168][6] ),
    .X(net4159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3754 (.A(\line_cache[170][0] ),
    .X(net4160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3755 (.A(\base_v_active[3] ),
    .X(net4161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3756 (.A(\line_cache[74][2] ),
    .X(net4162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3757 (.A(\line_cache[108][4] ),
    .X(net4163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3758 (.A(\line_cache[91][7] ),
    .X(net4164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3759 (.A(\line_cache[149][7] ),
    .X(net4165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_02308_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3760 (.A(\line_cache[110][5] ),
    .X(net4166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3761 (.A(\line_cache[71][5] ),
    .X(net4167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3762 (.A(\line_cache[126][2] ),
    .X(net4168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3763 (.A(\line_cache[207][5] ),
    .X(net4169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3764 (.A(\line_cache[87][0] ),
    .X(net4170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3765 (.A(_03729_),
    .X(net4171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3766 (.A(\line_cache[168][4] ),
    .X(net4172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3767 (.A(\line_cache[149][5] ),
    .X(net4173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3768 (.A(\line_cache[165][5] ),
    .X(net4174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3769 (.A(\line_cache[206][1] ),
    .X(net4175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\line_cache[25][6] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3770 (.A(\line_cache[91][4] ),
    .X(net4176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3771 (.A(\line_cache[90][1] ),
    .X(net4177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3772 (.A(\line_cache[107][6] ),
    .X(net4178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3773 (.A(net115),
    .X(net4179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3774 (.A(_02604_),
    .X(net4180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3775 (.A(\line_cache[174][7] ),
    .X(net4181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3776 (.A(net114),
    .X(net4182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3777 (.A(_02603_),
    .X(net4183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3778 (.A(\line_cache[108][3] ),
    .X(net4184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3779 (.A(\base_h_active[9] ),
    .X(net4185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_01422_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3780 (.A(\res_h_counter[5] ),
    .X(net4186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3781 (.A(_02702_),
    .X(net4187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3782 (.A(\base_v_bporch[2] ),
    .X(net4188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3783 (.A(\line_cache[149][0] ),
    .X(net4189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3784 (.A(\line_cache[154][5] ),
    .X(net4190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3785 (.A(\line_cache[21][7] ),
    .X(net4191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3786 (.A(\line_cache[174][0] ),
    .X(net4192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3787 (.A(net112),
    .X(net4193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3788 (.A(_02601_),
    .X(net4194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3789 (.A(\line_cache[222][2] ),
    .X(net4195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\line_cache[124][7] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3790 (.A(\line_cache[202][2] ),
    .X(net4196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3791 (.A(\line_cache[139][7] ),
    .X(net4197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3792 (.A(\base_h_bporch[4] ),
    .X(net4198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3793 (.A(\line_cache[246][1] ),
    .X(net4199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3794 (.A(\line_cache[171][7] ),
    .X(net4200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3795 (.A(\line_cache[241][4] ),
    .X(net4201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3796 (.A(\line_cache[15][0] ),
    .X(net4202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3797 (.A(\base_h_active[3] ),
    .X(net4203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3798 (.A(\line_cache[105][5] ),
    .X(net4204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3799 (.A(\base_h_active[6] ),
    .X(net4205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_01776_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_00223_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3800 (.A(\line_cache[87][6] ),
    .X(net4206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3801 (.A(\line_cache[109][5] ),
    .X(net4207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3802 (.A(\line_cache[73][7] ),
    .X(net4208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3803 (.A(\base_h_active[2] ),
    .X(net4209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3804 (.A(\base_h_fporch[3] ),
    .X(net4210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3805 (.A(net113),
    .X(net4211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3806 (.A(_02602_),
    .X(net4212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3807 (.A(\line_cache[138][0] ),
    .X(net4213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3808 (.A(\line_cache[150][2] ),
    .X(net4214));
 sky130_fd_sc_hd__clkbuf_4 hold3809 (.A(\fb_read_state[2] ),
    .X(net4215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\line_cache[299][0] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3810 (.A(_07631_),
    .X(net4216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3811 (.A(\line_cache[172][2] ),
    .X(net4217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3812 (.A(\line_cache[250][1] ),
    .X(net4218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3813 (.A(\base_h_sync[3] ),
    .X(net4219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3814 (.A(\line_cache[70][5] ),
    .X(net4220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3815 (.A(net123),
    .X(net4221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3816 (.A(_02573_),
    .X(net4222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3817 (.A(net116),
    .X(net4223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3818 (.A(_02605_),
    .X(net4224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3819 (.A(\line_cache[171][5] ),
    .X(net4225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_01760_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3820 (.A(\line_cache[246][3] ),
    .X(net4226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3821 (.A(\line_cache[68][3] ),
    .X(net4227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3822 (.A(\line_cache[169][0] ),
    .X(net4228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3823 (.A(\base_v_counter[9] ),
    .X(net4229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3824 (.A(_02696_),
    .X(net4230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3825 (.A(\line_cache[245][5] ),
    .X(net4231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3826 (.A(\line_cache[249][7] ),
    .X(net4232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3827 (.A(\line_cache[144][6] ),
    .X(net4233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3828 (.A(\base_h_active[8] ),
    .X(net4234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3829 (.A(\line_cache[102][2] ),
    .X(net4235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\line_cache[297][4] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3830 (.A(\base_h_active[5] ),
    .X(net4236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3831 (.A(\base_v_active[7] ),
    .X(net4237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3832 (.A(\line_cache[250][6] ),
    .X(net4238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3833 (.A(\line_cache[248][3] ),
    .X(net4239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3834 (.A(\line_cache[245][7] ),
    .X(net4240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3835 (.A(\line_cache[165][7] ),
    .X(net4241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3836 (.A(net109),
    .X(net4242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3837 (.A(_02598_),
    .X(net4243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3838 (.A(\line_cache[136][3] ),
    .X(net4244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3839 (.A(\line_cache[221][5] ),
    .X(net4245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_01748_),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3840 (.A(\line_cache[150][1] ),
    .X(net4246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3841 (.A(\base_h_active[1] ),
    .X(net4247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3842 (.A(\line_cache[100][3] ),
    .X(net4248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3843 (.A(\line_cache[15][6] ),
    .X(net4249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3844 (.A(\line_cache[100][2] ),
    .X(net4250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3845 (.A(\line_cache[271][6] ),
    .X(net4251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3846 (.A(\line_cache[168][7] ),
    .X(net4252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3847 (.A(_11503_),
    .X(net4253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3848 (.A(\line_cache[107][4] ),
    .X(net4254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3849 (.A(\line_cache[145][3] ),
    .X(net4255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\line_cache[134][5] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3850 (.A(\line_cache[86][0] ),
    .X(net4256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3851 (.A(net118),
    .X(net4257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3852 (.A(_02607_),
    .X(net4258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3853 (.A(\line_cache[170][5] ),
    .X(net4259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3854 (.A(\line_cache[150][7] ),
    .X(net4260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3855 (.A(\line_cache[26][2] ),
    .X(net4261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3856 (.A(\line_cache[174][1] ),
    .X(net4262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3857 (.A(\line_cache[205][7] ),
    .X(net4263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3858 (.A(\line_cache[175][1] ),
    .X(net4264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3859 (.A(\line_cache[144][3] ),
    .X(net4265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_00309_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3860 (.A(\base_h_counter[6] ),
    .X(net4266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3861 (.A(_02683_),
    .X(net4267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3862 (.A(\line_cache[175][4] ),
    .X(net4268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3863 (.A(\line_cache[89][0] ),
    .X(net4269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3864 (.A(net94),
    .X(net4270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3865 (.A(_02583_),
    .X(net4271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3866 (.A(\line_cache[26][1] ),
    .X(net4272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3867 (.A(net117),
    .X(net4273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3868 (.A(_02606_),
    .X(net4274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3869 (.A(\line_cache[27][3] ),
    .X(net4275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\line_cache[173][2] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3870 (.A(\prescaler_counter[4] ),
    .X(net4276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3871 (.A(_04983_),
    .X(net4277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3872 (.A(_04985_),
    .X(net4278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3873 (.A(\line_cache[246][2] ),
    .X(net4279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3874 (.A(\line_cache[205][5] ),
    .X(net4280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3875 (.A(\line_cache_idx[9] ),
    .X(net4281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3876 (.A(\line_cache[101][4] ),
    .X(net4282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3877 (.A(\line_cache[26][3] ),
    .X(net4283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3878 (.A(\line_cache[69][7] ),
    .X(net4284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3879 (.A(net119),
    .X(net4285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_00650_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3880 (.A(_02608_),
    .X(net4286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3881 (.A(\res_h_active[4] ),
    .X(net4287));
 sky130_fd_sc_hd__buf_1 hold3882 (.A(\res_h_counter[4] ),
    .X(net4288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3883 (.A(\base_v_counter[2] ),
    .X(net4289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3884 (.A(_02689_),
    .X(net4290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3885 (.A(\line_cache[72][3] ),
    .X(net4291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3886 (.A(\resolution[0] ),
    .X(net4292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3887 (.A(\line_cache[255][0] ),
    .X(net4293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3888 (.A(\prescaler_counter[1] ),
    .X(net4294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3889 (.A(\line_cache[0][7] ),
    .X(net4295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\line_cache[39][2] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3890 (.A(_00007_),
    .X(net4296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3891 (.A(\line_cache_idx[2] ),
    .X(net4297));
 sky130_fd_sc_hd__buf_1 hold3892 (.A(\base_v_counter[6] ),
    .X(net4298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3893 (.A(_02693_),
    .X(net4299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3894 (.A(\base_v_counter[3] ),
    .X(net4300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3895 (.A(_02690_),
    .X(net4301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3896 (.A(\line_cache[0][6] ),
    .X(net4302));
 sky130_fd_sc_hd__clkbuf_2 hold3897 (.A(\base_v_counter[0] ),
    .X(net4303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3898 (.A(_02687_),
    .X(net4304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3899 (.A(\line_cache[251][0] ),
    .X(net4305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\line_cache[211][1] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_02018_),
    .X(net796));
 sky130_fd_sc_hd__buf_1 hold3900 (.A(\base_v_counter[4] ),
    .X(net4306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3901 (.A(_02691_),
    .X(net4307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3902 (.A(\line_cache[271][7] ),
    .X(net4308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3903 (.A(\line_cache[255][5] ),
    .X(net4309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3904 (.A(\base_h_counter[1] ),
    .X(net4310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3905 (.A(_02678_),
    .X(net4311));
 sky130_fd_sc_hd__buf_1 hold3906 (.A(\base_v_counter[1] ),
    .X(net4312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3907 (.A(_02688_),
    .X(net4313));
 sky130_fd_sc_hd__buf_1 hold3908 (.A(\prescaler_counter[3] ),
    .X(net4314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3909 (.A(_08625_),
    .X(net4315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\line_cache[247][6] ),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_2 hold3910 (.A(_08632_),
    .X(net4316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3911 (.A(_02570_),
    .X(net4317));
 sky130_fd_sc_hd__clkbuf_2 hold3912 (.A(\base_v_counter[8] ),
    .X(net4318));
 sky130_fd_sc_hd__buf_1 hold3913 (.A(\base_h_counter[0] ),
    .X(net4319));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3914 (.A(\base_h_counter[2] ),
    .X(net4320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3915 (.A(\base_v_counter[7] ),
    .X(net4321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3916 (.A(\prescaler_counter[2] ),
    .X(net4322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3917 (.A(\base_h_counter[3] ),
    .X(net4323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3918 (.A(\prescaler_counter[6] ),
    .X(net4324));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3919 (.A(\base_v_counter[5] ),
    .X(net4325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_01310_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3920 (.A(\line_cache[287][6] ),
    .X(net4326));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3921 (.A(\base_h_counter[5] ),
    .X(net4327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3922 (.A(\line_cache[287][1] ),
    .X(net4328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3923 (.A(\line_cache[287][7] ),
    .X(net4329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3924 (.A(\line_cache[271][0] ),
    .X(net4330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3925 (.A(net98),
    .X(net4331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3926 (.A(_07687_),
    .X(net4332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3927 (.A(net121),
    .X(net4333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3928 (.A(_07777_),
    .X(net4334));
 sky130_fd_sc_hd__buf_1 hold3929 (.A(_08632_),
    .X(net4335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\line_cache[29][4] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3930 (.A(\line_cache_idx[2] ),
    .X(net4336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3931 (.A(\line_cache_idx[6] ),
    .X(net4337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_01772_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\line_cache[153][0] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_00472_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\line_cache[77][6] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_02358_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\line_cache[184][7] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00235_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_00993_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_00751_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\line_cache[25][0] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_01416_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\line_cache[2][7] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_01783_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\line_cache[259][1] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_01409_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\line_cache[177][2] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_00682_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\line_cache[259][4] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\line_cache[242][7] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_01412_),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\line_cache[312][7] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_01895_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\line_cache[42][5] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_02053_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\line_cache[84][1] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_02417_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\line_cache[206][3] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_00947_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\line_cache[245][3] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_01271_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_01291_),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\line_cache[135][1] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_00313_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\line_cache[315][6] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_01918_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\line_cache[71][2] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_02306_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\line_cache[98][4] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_02540_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\line_cache[12][5] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\line_cache[214][5] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_00269_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\line_cache[240][5] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_01253_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\line_cache[81][2] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_02394_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\line_cache[85][3] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_02427_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\line_cache[150][4] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_00452_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\line_cache[189][6] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_01021_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_00790_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\line_cache[295][1] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_01729_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\line_cache[3][5] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_02029_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\line_cache[218][3] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_01051_),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\line_cache[86][3] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_02435_),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\line_cache[38][7] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\line_cache[74][3] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_02015_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\line_cache[136][2] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_00322_),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\line_cache[275][0] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_01552_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\line_cache[288][1] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_01665_),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\line_cache[11][0] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_00176_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\line_cache[303][0] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_02331_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_01808_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\line_cache[102][7] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_00031_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\line_cache[69][4] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_02284_),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\line_cache[198][4] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_00868_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\line_cache[280][7] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_01607_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\line_cache[33][0] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\line_cache[242][4] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_01968_),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\line_cache[282][5] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_01621_),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\line_cache[81][4] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_02396_),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\line_cache[38][5] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_02013_),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\line_cache[84][5] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_02421_),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\line_cache[246][7] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_01268_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_01303_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\line_cache[21][4] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_01068_),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\line_cache[159][2] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_00522_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\line_cache[162][7] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_00559_),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\line_cache[167][4] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_00596_),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\line_cache[66][5] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\line_cache[214][3] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_02261_),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\line_cache[108][7] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_00079_),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\line_cache[86][5] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_02437_),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\line_cache[259][0] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_01408_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\line_cache[166][3] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_00587_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\line_cache[70][3] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\line_cache[162][0] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_01019_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_02299_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\line_cache[109][3] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_00083_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\line_cache[235][0] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_01200_),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\line_cache[265][0] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_01464_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\line_cache[70][6] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_02302_),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\line_cache[258][5] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\line_cache[243][6] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_01405_),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\line_cache[125][1] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_00225_),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\line_cache[125][0] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_00224_),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\line_cache[165][3] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_00579_),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\line_cache[102][4] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_00028_),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\line_cache[220][2] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_01278_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_01074_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\line_cache[177][0] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_00680_),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\line_cache[3][3] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_02027_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\line_cache[267][1] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_01481_),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\line_cache[158][5] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_00517_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\line_cache[246][0] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\line_cache[25][4] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_01296_),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\line_cache[102][6] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_00030_),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\line_cache[155][5] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_00493_),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\line_cache[104][1] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_00041_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\line_cache[191][3] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_00811_),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\line_cache[132][0] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_01420_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_00288_),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\line_cache[81][0] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_02392_),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\line_cache[188][2] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_00778_),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\line_cache[173][6] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_00654_),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\line_cache[62][3] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_02227_),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\line_cache[234][5] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\line_cache[133][4] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_01197_),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\line_cache[9][2] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_02554_),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\line_cache[66][4] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_02260_),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\line_cache[224][2] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_01106_),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\line_cache[218][7] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_01055_),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\line_cache[158][7] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_00300_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_00519_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\line_cache[150][6] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_00454_),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\line_cache[99][1] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_02545_),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\line_cache[306][0] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_01832_),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\line_cache[72][5] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_02317_),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\line_cache[125][2] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\line_cache[132][2] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_00226_),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\line_cache[293][2] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_01714_),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\line_cache[91][1] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_02481_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\line_cache[206][5] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_00949_),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\line_cache[85][4] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_02428_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\line_cache[303][6] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_00290_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_01814_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\line_cache[239][7] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_01239_),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\line_cache[69][2] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_02282_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\line_cache[151][4] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_00460_),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\line_cache[125][6] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_00230_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\line_cache[108][1] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\line_cache[211][6] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_00073_),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\line_cache[206][7] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_00951_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\line_cache[294][5] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_01725_),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\line_cache[62][7] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_02231_),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\line_cache[290][5] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_01693_),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\line_cache[307][1] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_00552_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_00998_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_01841_),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\line_cache[167][1] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_00593_),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\line_cache[62][5] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_02229_),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\line_cache[246][5] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_01301_),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\line_cache[238][7] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_01231_),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\line_cache[49][4] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\line_cache[186][0] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_02108_),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\line_cache[138][7] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_00343_),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\line_cache[309][2] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_01858_),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\line_cache[302][6] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_01806_),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\line_cache[254][5] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_01373_),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\line_cache[220][0] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_00760_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_01072_),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\line_cache[141][4] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_00372_),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\line_cache[234][4] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_01196_),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\line_cache[134][4] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_00308_),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\line_cache[178][5] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_00693_),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\line_cache[201][4] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\line_cache[243][1] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_00908_),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\line_cache[307][3] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_01843_),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\line_cache[318][2] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_01938_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\line_cache[56][1] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_02169_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\line_cache[91][3] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_02483_),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\line_cache[51][2] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_01273_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_02130_),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\line_cache[310][7] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_01879_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\line_cache[18][4] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_00796_),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\line_cache[244][2] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_01282_),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\line_cache[211][3] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_00995_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\line_cache[249][4] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\line_cache[1][2] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_01324_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\line_cache[205][3] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_00939_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\line_cache[294][7] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_01727_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\line_cache[138][4] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_00340_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\line_cache[84][0] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_02416_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\line_cache[174][3] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_00890_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_00659_),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\line_cache[9][6] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_02558_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\line_cache[172][0] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_00640_),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\line_cache[42][6] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_02054_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\line_cache[177][4] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_00684_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\line_cache[210][4] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\line_cache[137][2] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_00988_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\line_cache[90][4] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_02476_),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\line_cache[97][2] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_02530_),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\line_cache[99][4] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_02548_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\line_cache[230][4] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_01164_),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\line_cache[43][5] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_00330_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_02061_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\line_cache[134][0] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_00304_),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\line_cache[311][1] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_01881_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\line_cache[175][7] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_00671_),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\line_cache[59][0] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_02192_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\line_cache[66][3] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\line_cache[318][0] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_02259_),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\line_cache[34][0] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_01976_),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\line_cache[77][2] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_02354_),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\line_cache[59][1] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_02193_),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\line_cache[128][1] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_00249_),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\line_cache[163][6] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\line_cache[137][1] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_01936_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_00566_),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\line_cache[10][0] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_00088_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\line_cache[30][3] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_01867_),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\line_cache[202][0] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_00912_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\line_cache[245][2] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_01290_),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\line_cache[79][0] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\line_cache[126][6] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_02368_),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\line_cache[42][7] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_02055_),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\line_cache[88][5] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(_02453_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\line_cache[25][1] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_01417_),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\line_cache[140][7] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_00367_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\line_cache[148][1] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_00238_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_00425_),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\line_cache[166][5] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_00589_),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\line_cache[266][5] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_01477_),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\line_cache[317][4] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_01932_),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\line_cache[153][6] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_00478_),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\line_cache[106][6] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\line_cache[241][6] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_00062_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\line_cache[79][1] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_02369_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\line_cache[133][6] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_00302_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\line_cache[314][6] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_01910_),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\line_cache[303][2] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_01810_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\line_cache[245][4] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_01262_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_01292_),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\line_cache[141][0] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_00368_),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\line_cache[189][1] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_00785_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\line_cache[109][6] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_00086_),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\line_cache[270][4] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_01516_),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\line_cache[212][1] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\line_cache[229][0] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_01001_),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\line_cache[164][2] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_00570_),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\line_cache[103][1] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_00033_),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\line_cache[146][0] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_00408_),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\line_cache[153][4] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_00476_),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\line_cache[111][5] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_01144_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_00109_),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\line_cache[104][5] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_00045_),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\line_cache[82][6] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_02406_),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\line_cache[75][7] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_02343_),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\line_cache[312][4] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_01892_),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\line_cache[297][2] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\line_cache[319][0] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_01746_),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\line_cache[50][4] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_02124_),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\line_cache[267][4] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_01484_),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\line_cache[149][2] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_00434_),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\line_cache[182][0] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_00728_),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\line_cache[135][0] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_01944_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_00312_),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\line_cache[11][6] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_00182_),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\line_cache[165][2] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_00578_),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\line_cache[94][0] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_02504_),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\line_cache[90][6] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_02478_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\line_cache[246][6] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\line_cache[132][4] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_01302_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\line_cache[39][6] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_02022_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\line_cache[142][5] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_00381_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\line_cache[54][5] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_02157_),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\line_cache[119][1] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_00169_),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\line_cache[22][4] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00329_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_00292_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_01156_),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\line_cache[299][2] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_01762_),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\line_cache[311][2] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_01882_),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\line_cache[290][3] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_01691_),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\line_cache[162][4] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_00556_),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\line_cache[39][1] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\line_cache[226][5] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_02017_),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\line_cache[231][6] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_01174_),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\line_cache[12][2] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_00266_),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\line_cache[83][2] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_02410_),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\line_cache[148][0] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_00424_),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\line_cache[253][0] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_01125_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_01360_),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\line_cache[131][1] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_00281_),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\line_cache[106][5] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_00061_),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\line_cache[165][4] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_00580_),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\line_cache[211][2] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_00994_),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\line_cache[152][2] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\line_cache[121][4] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_00466_),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\line_cache[139][2] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_00346_),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\line_cache[246][4] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_01300_),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\line_cache[110][3] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_00099_),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\line_cache[198][3] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_00867_),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\line_cache[228][0] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_00196_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(_01136_),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\line_cache[108][0] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_00072_),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\line_cache[51][0] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_02128_),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\line_cache[91][6] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_02486_),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\line_cache[76][2] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_02346_),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\line_cache[189][0] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\line_cache[3][2] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_00784_),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\line_cache[18][3] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_00795_),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\line_cache[301][2] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_01794_),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\line_cache[282][3] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_01619_),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\line_cache[50][7] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_02127_),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\line_cache[18][7] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_02026_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_00799_),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\line_cache[257][1] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_01393_),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\line_cache[41][6] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_02046_),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\line_cache[35][1] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_01985_),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\line_cache[299][6] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_01766_),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\line_cache[124][0] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\line_cache[230][0] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_00216_),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\line_cache[105][4] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(_00052_),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\line_cache[172][1] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_00641_),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\line_cache[76][0] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_02344_),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\line_cache[58][5] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_02189_),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\line_cache[200][0] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_01160_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_00896_),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\line_cache[264][2] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_01458_),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\line_cache[175][3] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_00667_),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\line_cache[97][4] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_02532_),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\line_cache[203][4] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_00924_),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\line_cache[127][5] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\line_cache[206][0] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_00245_),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\line_cache[83][7] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_02415_),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\line_cache[159][6] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_00526_),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\line_cache[167][0] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_00592_),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\line_cache[101][6] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_00022_),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\line_cache[308][1] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\line_cache[121][2] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_00944_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_01849_),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\line_cache[127][2] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_00242_),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\line_cache[33][3] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_01971_),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\line_cache[238][0] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_01224_),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\line_cache[309][4] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_01860_),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\line_cache[110][7] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\line_cache[30][0] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_00103_),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\line_cache[179][2] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_00698_),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\line_cache[107][2] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_00066_),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\line_cache[50][3] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_02123_),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\line_cache[73][3] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_02323_),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\line_cache[23][2] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_01864_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_01242_),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\line_cache[91][5] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_02485_),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\line_cache[40][2] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_02034_),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\line_cache[266][7] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_01479_),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\line_cache[80][1] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_02385_),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\line_cache[202][3] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\line_cache[40][0] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_00915_),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\line_cache[304][1] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_01817_),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\line_cache[81][1] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_02393_),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\line_cache[107][5] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_00069_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\line_cache[70][7] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_02303_),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\line_cache[79][5] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_02032_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_02373_),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\line_cache[75][6] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_02342_),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\line_cache[269][4] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_01500_),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\line_cache[30][5] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_01869_),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\line_cache[245][6] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_01294_),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\line_cache[130][7] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\line_cache[243][4] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_00279_),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\line_cache[310][3] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_01875_),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\line_cache[1][3] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_00891_),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\line_cache[88][4] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(_02452_),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\line_cache[111][6] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_00110_),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\line_cache[223][6] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_01276_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_01102_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\line_cache[43][0] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_02056_),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\line_cache[181][2] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_00722_),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\line_cache[185][0] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_00752_),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\line_cache[29][6] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_01774_),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\line_cache[251][1] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\line_cache[65][4] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_01345_),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\line_cache[313][6] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_01902_),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\line_cache[191][2] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_00810_),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\line_cache[221][4] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_01084_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\line_cache[50][5] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_02125_),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\line_cache[24][0] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_02252_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_01328_),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\line_cache[303][7] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_01815_),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\line_cache[43][7] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_02063_),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\line_cache[178][4] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_00692_),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\line_cache[136][5] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_00325_),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\line_cache[134][7] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\line_cache[2][3] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_00311_),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\line_cache[62][4] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_02228_),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\line_cache[38][6] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_02014_),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\line_cache[247][0] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_01304_),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\line_cache[306][7] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_01839_),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\line_cache[149][1] ),
    .X(net1405));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(base_h_active_i[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(base_h_active_i[9]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(base_h_bporch_i[0]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(base_h_bporch_i[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(base_h_bporch_i[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(base_h_bporch_i[3]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(base_h_bporch_i[4]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(base_h_bporch_i[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(base_h_bporch_i[6]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(base_h_fporch_i[0]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(base_h_fporch_i[1]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(base_h_active_i[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(base_h_fporch_i[2]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(base_h_fporch_i[3]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(base_h_fporch_i[4]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(base_h_sync_i[0]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(base_h_sync_i[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(base_h_sync_i[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(base_h_sync_i[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(base_h_sync_i[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(base_h_sync_i[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(base_h_sync_i[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(base_h_active_i[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(base_v_active_i[0]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(base_v_active_i[1]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(base_v_active_i[2]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(base_v_active_i[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(base_v_active_i[4]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(base_v_active_i[5]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(base_v_active_i[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(base_v_active_i[7]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(base_v_active_i[8]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(base_v_bporch_i[0]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(base_h_active_i[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(base_v_bporch_i[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(base_v_bporch_i[2]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(base_v_bporch_i[3]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(base_v_fporch_i[0]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(base_v_fporch_i[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(base_v_fporch_i[2]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(base_v_sync_i[0]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(base_v_sync_i[1]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(base_v_sync_i[2]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(enable_i),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(base_h_active_i[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_8 input50 (.A(mport_i[0]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 input51 (.A(mport_i[10]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_16 input52 (.A(mport_i[11]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(mport_i[12]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(mport_i[13]),
    .X(net54));
 sky130_fd_sc_hd__buf_8 input55 (.A(mport_i[14]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(mport_i[15]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(mport_i[16]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(mport_i[17]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(mport_i[18]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(base_h_active_i[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input60 (.A(mport_i[19]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(mport_i[1]),
    .X(net61));
 sky130_fd_sc_hd__buf_6 input62 (.A(mport_i[20]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(mport_i[21]),
    .X(net63));
 sky130_fd_sc_hd__buf_12 input64 (.A(mport_i[22]),
    .X(net64));
 sky130_fd_sc_hd__buf_6 input65 (.A(mport_i[23]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(mport_i[24]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(mport_i[25]),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input68 (.A(mport_i[26]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_16 input69 (.A(mport_i[27]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(base_h_active_i[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input70 (.A(mport_i[28]),
    .X(net70));
 sky130_fd_sc_hd__buf_8 input71 (.A(mport_i[29]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 input72 (.A(mport_i[2]),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(mport_i[30]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_16 input74 (.A(mport_i[31]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(mport_i[33]),
    .X(net75));
 sky130_fd_sc_hd__buf_4 input76 (.A(mport_i[3]),
    .X(net76));
 sky130_fd_sc_hd__buf_6 input77 (.A(mport_i[4]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_16 input78 (.A(mport_i[5]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(mport_i[6]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(base_h_active_i[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input80 (.A(mport_i[7]),
    .X(net80));
 sky130_fd_sc_hd__buf_6 input81 (.A(mport_i[8]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_16 input82 (.A(mport_i[9]),
    .X(net82));
 sky130_fd_sc_hd__buf_2 input83 (.A(nrst_i),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(prescaler_i[0]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(prescaler_i[1]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(prescaler_i[2]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(prescaler_i[3]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(resolution_i[0]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(resolution_i[1]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(base_h_active_i[8]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(resolution_i[2]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(resolution_i[3]),
    .X(net91));
 sky130_fd_sc_hd__buf_12 load_slew137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 load_slew138 (.A(_09414_),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_16 load_slew139 (.A(_09287_),
    .X(net139));
 sky130_fd_sc_hd__buf_12 load_slew141 (.A(_09494_),
    .X(net141));
 sky130_fd_sc_hd__buf_6 load_slew142 (.A(_09440_),
    .X(net142));
 sky130_fd_sc_hd__buf_8 load_slew146 (.A(_09218_),
    .X(net146));
 sky130_fd_sc_hd__buf_12 max_cap135 (.A(_09530_),
    .X(net135));
 sky130_fd_sc_hd__buf_12 max_cap136 (.A(_09504_),
    .X(net136));
 sky130_fd_sc_hd__buf_12 max_cap140 (.A(_09283_),
    .X(net140));
 sky130_fd_sc_hd__buf_8 max_cap143 (.A(_09331_),
    .X(net143));
 sky130_fd_sc_hd__buf_12 max_cap144 (.A(_09268_),
    .X(net144));
 sky130_fd_sc_hd__buf_12 max_cap145 (.A(_09262_),
    .X(net145));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(mport_o[41]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(mport_o[42]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(mport_o[43]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(mport_o[44]));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(mport_o[45]));
 sky130_fd_sc_hd__buf_12 output105 (.A(net105),
    .X(mport_o[46]));
 sky130_fd_sc_hd__buf_12 output106 (.A(net106),
    .X(mport_o[47]));
 sky130_fd_sc_hd__buf_12 output107 (.A(net107),
    .X(mport_o[48]));
 sky130_fd_sc_hd__buf_12 output108 (.A(net108),
    .X(mport_o[49]));
 sky130_fd_sc_hd__buf_12 output109 (.A(net109),
    .X(mport_o[50]));
 sky130_fd_sc_hd__buf_12 output110 (.A(net110),
    .X(mport_o[51]));
 sky130_fd_sc_hd__buf_12 output111 (.A(net111),
    .X(mport_o[52]));
 sky130_fd_sc_hd__buf_12 output112 (.A(net112),
    .X(mport_o[53]));
 sky130_fd_sc_hd__buf_12 output113 (.A(net113),
    .X(mport_o[54]));
 sky130_fd_sc_hd__buf_12 output114 (.A(net114),
    .X(mport_o[55]));
 sky130_fd_sc_hd__buf_12 output115 (.A(net115),
    .X(mport_o[56]));
 sky130_fd_sc_hd__buf_12 output116 (.A(net116),
    .X(mport_o[57]));
 sky130_fd_sc_hd__buf_12 output117 (.A(net117),
    .X(mport_o[58]));
 sky130_fd_sc_hd__buf_12 output118 (.A(net118),
    .X(mport_o[59]));
 sky130_fd_sc_hd__buf_12 output119 (.A(net119),
    .X(mport_o[60]));
 sky130_fd_sc_hd__buf_12 output120 (.A(net120),
    .X(mport_o[61]));
 sky130_fd_sc_hd__buf_12 output121 (.A(net121),
    .X(mport_o[62]));
 sky130_fd_sc_hd__buf_12 output122 (.A(net122),
    .X(mport_o[63]));
 sky130_fd_sc_hd__buf_12 output123 (.A(net123),
    .X(mport_o[64]));
 sky130_fd_sc_hd__buf_12 output124 (.A(net124),
    .X(mport_o[66]));
 sky130_fd_sc_hd__buf_12 output125 (.A(net125),
    .X(mport_o[67]));
 sky130_fd_sc_hd__buf_12 output126 (.A(net126),
    .X(pixel_o[0]));
 sky130_fd_sc_hd__buf_12 output127 (.A(net127),
    .X(pixel_o[1]));
 sky130_fd_sc_hd__buf_12 output128 (.A(net128),
    .X(pixel_o[2]));
 sky130_fd_sc_hd__buf_12 output129 (.A(net129),
    .X(pixel_o[3]));
 sky130_fd_sc_hd__buf_12 output130 (.A(net130),
    .X(pixel_o[4]));
 sky130_fd_sc_hd__buf_12 output131 (.A(net131),
    .X(pixel_o[5]));
 sky130_fd_sc_hd__buf_12 output132 (.A(net132),
    .X(pixel_o[6]));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(pixel_o[7]));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(vsync_o));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(hsync_o));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(mport_o[34]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(mport_o[35]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(mport_o[36]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(mport_o[37]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(mport_o[38]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(mport_o[39]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(mport_o[40]));
 sky130_fd_sc_hd__conb_1 vga_m_371 (.LO(net371));
 sky130_fd_sc_hd__conb_1 vga_m_372 (.LO(net372));
 sky130_fd_sc_hd__conb_1 vga_m_373 (.LO(net373));
 sky130_fd_sc_hd__conb_1 vga_m_374 (.LO(net374));
 sky130_fd_sc_hd__conb_1 vga_m_375 (.LO(net375));
 sky130_fd_sc_hd__conb_1 vga_m_376 (.LO(net376));
 sky130_fd_sc_hd__conb_1 vga_m_377 (.LO(net377));
 sky130_fd_sc_hd__conb_1 vga_m_378 (.LO(net378));
 sky130_fd_sc_hd__conb_1 vga_m_379 (.LO(net379));
 sky130_fd_sc_hd__conb_1 vga_m_380 (.LO(net380));
 sky130_fd_sc_hd__conb_1 vga_m_381 (.LO(net381));
 sky130_fd_sc_hd__conb_1 vga_m_382 (.LO(net382));
 sky130_fd_sc_hd__conb_1 vga_m_383 (.LO(net383));
 sky130_fd_sc_hd__conb_1 vga_m_384 (.LO(net384));
 sky130_fd_sc_hd__conb_1 vga_m_385 (.LO(net385));
 sky130_fd_sc_hd__conb_1 vga_m_386 (.LO(net386));
 sky130_fd_sc_hd__conb_1 vga_m_387 (.LO(net387));
 sky130_fd_sc_hd__conb_1 vga_m_388 (.LO(net388));
 sky130_fd_sc_hd__conb_1 vga_m_389 (.LO(net389));
 sky130_fd_sc_hd__conb_1 vga_m_390 (.LO(net390));
 sky130_fd_sc_hd__conb_1 vga_m_391 (.LO(net391));
 sky130_fd_sc_hd__conb_1 vga_m_392 (.LO(net392));
 sky130_fd_sc_hd__conb_1 vga_m_393 (.LO(net393));
 sky130_fd_sc_hd__conb_1 vga_m_394 (.LO(net394));
 sky130_fd_sc_hd__conb_1 vga_m_395 (.LO(net395));
 sky130_fd_sc_hd__conb_1 vga_m_396 (.LO(net396));
 sky130_fd_sc_hd__conb_1 vga_m_397 (.LO(net397));
 sky130_fd_sc_hd__conb_1 vga_m_398 (.LO(net398));
 sky130_fd_sc_hd__conb_1 vga_m_399 (.LO(net399));
 sky130_fd_sc_hd__conb_1 vga_m_400 (.LO(net400));
 sky130_fd_sc_hd__conb_1 vga_m_401 (.LO(net401));
 sky130_fd_sc_hd__conb_1 vga_m_402 (.LO(net402));
 sky130_fd_sc_hd__conb_1 vga_m_403 (.LO(net403));
 sky130_fd_sc_hd__conb_1 vga_m_404 (.LO(net404));
 sky130_fd_sc_hd__conb_1 vga_m_405 (.LO(net405));
 sky130_fd_sc_hd__conb_1 vga_m_406 (.LO(net406));
 assign mport_o[0] = net371;
 assign mport_o[10] = net381;
 assign mport_o[11] = net382;
 assign mport_o[12] = net383;
 assign mport_o[13] = net384;
 assign mport_o[14] = net385;
 assign mport_o[15] = net386;
 assign mport_o[16] = net387;
 assign mport_o[17] = net388;
 assign mport_o[18] = net389;
 assign mport_o[19] = net390;
 assign mport_o[1] = net372;
 assign mport_o[20] = net391;
 assign mport_o[21] = net392;
 assign mport_o[22] = net393;
 assign mport_o[23] = net394;
 assign mport_o[24] = net395;
 assign mport_o[25] = net396;
 assign mport_o[26] = net397;
 assign mport_o[27] = net398;
 assign mport_o[28] = net399;
 assign mport_o[29] = net400;
 assign mport_o[2] = net373;
 assign mport_o[30] = net401;
 assign mport_o[31] = net402;
 assign mport_o[32] = net403;
 assign mport_o[33] = net404;
 assign mport_o[3] = net374;
 assign mport_o[4] = net375;
 assign mport_o[5] = net376;
 assign mport_o[65] = net405;
 assign mport_o[68] = net406;
 assign mport_o[6] = net377;
 assign mport_o[7] = net378;
 assign mport_o[8] = net379;
 assign mport_o[9] = net380;
endmodule

