// This is the unpowered netlist.
module mac (clk,
    nrst,
    a_i,
    b_i,
    y_o);
 input clk;
 input nrst;
 input [31:0] a_i;
 input [31:0] b_i;
 output [31:0] y_o;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire \absum[0] ;
 wire \absum[10] ;
 wire \absum[11] ;
 wire \absum[12] ;
 wire \absum[13] ;
 wire \absum[14] ;
 wire \absum[15] ;
 wire \absum[16] ;
 wire \absum[17] ;
 wire \absum[18] ;
 wire \absum[19] ;
 wire \absum[1] ;
 wire \absum[20] ;
 wire \absum[21] ;
 wire \absum[22] ;
 wire \absum[23] ;
 wire \absum[24] ;
 wire \absum[25] ;
 wire \absum[26] ;
 wire \absum[27] ;
 wire \absum[28] ;
 wire \absum[29] ;
 wire \absum[2] ;
 wire \absum[30] ;
 wire \absum[31] ;
 wire \absum[3] ;
 wire \absum[4] ;
 wire \absum[5] ;
 wire \absum[6] ;
 wire \absum[7] ;
 wire \absum[8] ;
 wire \absum[9] ;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__05341__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05341__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05343__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__05345__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05345__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05351__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05351__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05358__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05358__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05360__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05360__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05362__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05362__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05371__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05375__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05375__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05381__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05398__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05398__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05400__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05400__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05402__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05407__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05407__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05409__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05409__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05414__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05414__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05424__A (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05424__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05427__A (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05427__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05433__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05434__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05434__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05445__A (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05445__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05447__A (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05447__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05451__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05452__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05452__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05465__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05465__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05482__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05482__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05485__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05485__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05490__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05490__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05505__A (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05505__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05507__A (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05507__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05513__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05514__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05514__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05539__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05539__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05545__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05545__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05549__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05549__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05551__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05551__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__05556__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05557__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05557__B (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05567__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05567__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05568__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05568__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05574__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05574__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__05586__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05586__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05588__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__05589__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05589__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05594__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05595__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05595__B (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05606__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05606__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05607__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05608__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05608__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05613__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05613__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__05641__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05641__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05643__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05643__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05644__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05644__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05658__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05658__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05659__A (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05659__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05661__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05661__B (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05686__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05686__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05687__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05688__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05688__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05690__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05704__A (.DIODE(_03611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05704__B (.DIODE(_04304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05719__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05719__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05728__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05728__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05734__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__05735__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05735__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05747__A (.DIODE(_04304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05747__B (.DIODE(_03611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05751__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05751__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__05753__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05753__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__05760__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05760__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05767__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05767__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05780__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05780__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05781__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05781__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__05783__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05783__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__05805__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05805__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05808__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05808__B (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05813__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__05813__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__05819__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05819__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05820__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05820__B (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05822__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05822__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05829__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05830__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__05830__B (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05845__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05845__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05845__C (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05845__D (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05863__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05863__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05864__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05864__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05866__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05866__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05871__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05871__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05872__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05872__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05874__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05874__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__05901__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__05901__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05903__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05903__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05908__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05908__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05919__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05919__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05921__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05921__B (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05926__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05926__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05938__A (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05938__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05939__A (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05940__A (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05940__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05944__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05944__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05967__A (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05968__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05968__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05970__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05970__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05975__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05975__B (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05984__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05985__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05986__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05986__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05987__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05987__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06023__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06023__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06025__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06025__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06030__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06031__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06031__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06047__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06047__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06048__B (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06048__C (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06049__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06050__A (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06053__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06053__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06063__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06063__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__B (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06127__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06127__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__06128__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06128__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06130__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06130__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__B (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__B (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06148__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06148__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06149__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06150__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06150__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__06152__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06152__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06181__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__A1 (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__A2 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__B1 (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__B2 (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06191__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06191__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06192__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06192__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06194__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06194__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__06204__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06204__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06205__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06205__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06207__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06207__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06224__A (.DIODE(_03611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06225__A (.DIODE(_04304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06228__B (.DIODE(_04304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06229__B (.DIODE(_03611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06270__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06270__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06271__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06271__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06326__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06326__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06327__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06327__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06329__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06329__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__B (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06336__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06336__B (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06339__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06339__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06347__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06347__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06348__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__06351__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06351__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06389__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06389__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06390__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06390__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06397__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06398__A (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06399__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06399__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06400__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06400__B (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06405__A (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06405__B (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__A (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06444__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06512__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06515__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06516__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06516__B (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__A (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__B (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__B (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06536__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06537__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06537__B (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06539__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06539__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A1 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A2 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__B (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06630__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__A (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__B (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__A (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__A (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__A (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06748__A1 (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__B (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__B (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__C (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__B (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__B (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__B (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__B (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__B (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__B (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__B (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__B (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__B (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__B (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__B (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__B (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__B (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__B (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__B (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__B (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__B (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A1 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A2 (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__B (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__B (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__B (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__B (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__B (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__B (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__B (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__C (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__D (.DIODE(_02522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__B (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__B (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__B (.DIODE(_01257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A (.DIODE(_01727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__B (.DIODE(_01727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A1 (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A2 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B1 (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B2 (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07881__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B (.DIODE(_01224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__B (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__B (.DIODE(_01893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A (.DIODE(_01893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__B (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__B (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__B (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__B (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__B (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__A (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__B (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A (.DIODE(_01893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B (.DIODE(_01893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__B (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__B (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__B (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A1 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A2 (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__B (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__A (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__B (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__B (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__B (.DIODE(_00641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__B (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__B (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__B (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__B (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A_N (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A_N (.DIODE(_02177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__B (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__B (.DIODE(_02177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A1 (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A2 (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__B1 (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__B2 (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__B (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__C (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__D (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__C (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__D (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A2 (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__B1 (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__B2 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__C (.DIODE(_02177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__B (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__B (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__C (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__A (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__B (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__C (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__A1 (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__C (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__B (.DIODE(_02177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__B1 (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__B (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__A (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A_N (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__A (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A1 (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__A (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__B (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A2 (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__B (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__B (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A1 (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__B (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__A (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__A (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__A (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A1 (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__B (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A2 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08724__A (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__B (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__A (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__B (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__B (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08900__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08900__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__C (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A2 (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__B2 (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__B (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__A (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__A1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__A2 (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__C (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__A (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__A (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09165__A (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A1 (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__A (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A1 (.DIODE(_01267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__B (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__B (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__B (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__B (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__B (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__B (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A1 (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__B1 (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__B (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__C (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__D (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A1 (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A2 (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B2 (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__B (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__C (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__D (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__A1 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__A2 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B1 (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B2 (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__C (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__D (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A2 (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__B1 (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__B2 (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__B (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__C (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__D (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A1 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A2 (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__B2 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__A (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__B (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__C (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__D (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A1 (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A2 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__B1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__B2 (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__B (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__C (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__D (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__A2 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__B1 (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__B2 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__C (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__D (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A2 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__B2 (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__C (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__D (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A2 (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__B2 (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__B (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__C (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__D (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A1 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A2 (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__B1 (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__B2 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__B (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__C (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__D (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A2 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__B1 (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__B2 (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__B (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A1 (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__B1 (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A2 (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A1 (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__B1 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09644__A2 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__A (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__B (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__C (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__A1 (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__B2 (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A2 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A3 (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A2 (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A3 (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__A (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__B (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__C (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__D (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__A1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__A2 (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__B1 (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__B2 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__A2 (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__A3 (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A1 (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A2 (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__B1 (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__B2 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__B (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__B (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__C (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__D (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A2 (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__B1 (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__B2 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__C (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__D (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__A2 (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__B2 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A2 (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A3 (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__C (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__D (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__A2 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__B2 (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__B (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A2 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09820__A (.DIODE(_03939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09820__B (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__B (.DIODE(_03939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__C (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__B (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A2 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__B2 (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__D (.DIODE(_02309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A2 (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__B2 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__C (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A2 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__B (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__B (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__D (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A2 (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__B1 (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__B2 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A2 (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09956__A1 (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09956__B1 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__B (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__A (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A1 (.DIODE(_00560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__A (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__A (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__C (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A1 (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A2 (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B1 (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B2 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__A1 (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__A2 (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__B1 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__B2 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__B (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__C (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__A (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__B (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__B (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__C (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__D (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A2 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B1 (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B2 (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A (.DIODE(_04236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__B (.DIODE(_04239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B (.DIODE(_04236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__C (.DIODE(_04239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A1 (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__B1 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__B (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A1 (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__A (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__A (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__A (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__B (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__B (.DIODE(_01895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__B (.DIODE(_05049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__A (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__B (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__B (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A1 (.DIODE(_00960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A2 (.DIODE(_04899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__B2 (.DIODE(_00520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__A1 (.DIODE(_01334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__A2 (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__B2 (.DIODE(_04936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__B (.DIODE(_05278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__A (.DIODE(_05191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__B (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__B (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A2 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B2 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A2 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__B2 (.DIODE(_00384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__A3 (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__B (.DIODE(_04236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A_N (.DIODE(_04236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__B (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__B (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__B (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10715__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10733__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net65));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__buf_6 _05339_ (.A(net58),
    .X(_00300_));
 sky130_fd_sc_hd__clkbuf_8 _05340_ (.A(net9),
    .X(_00311_));
 sky130_fd_sc_hd__nand2_1 _05341_ (.A(_00300_),
    .B(_00311_),
    .Y(_00322_));
 sky130_fd_sc_hd__inv_2 _05342_ (.A(_00322_),
    .Y(_00333_));
 sky130_fd_sc_hd__buf_6 _05343_ (.A(net55),
    .X(_00344_));
 sky130_fd_sc_hd__buf_6 _05344_ (.A(net10),
    .X(_00355_));
 sky130_fd_sc_hd__nand2_1 _05345_ (.A(_00344_),
    .B(_00355_),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _05346_ (.A(_00333_),
    .B(_00366_),
    .Y(_00377_));
 sky130_fd_sc_hd__inv_2 _05347_ (.A(_00366_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _05348_ (.A(_00388_),
    .B(_00322_),
    .Y(_00399_));
 sky130_fd_sc_hd__buf_6 _05349_ (.A(net44),
    .X(_00410_));
 sky130_fd_sc_hd__buf_4 _05350_ (.A(net11),
    .X(_00421_));
 sky130_fd_sc_hd__nand2_1 _05351_ (.A(_00410_),
    .B(_00421_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand3_1 _05352_ (.A(_00377_),
    .B(_00399_),
    .C(_00432_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _05353_ (.A(_00388_),
    .B(_00333_),
    .Y(_00454_));
 sky130_fd_sc_hd__inv_2 _05354_ (.A(_00432_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _05355_ (.A(_00366_),
    .B(_00322_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand3_1 _05356_ (.A(_00454_),
    .B(_00465_),
    .C(_00476_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _05357_ (.A(_00443_),
    .B(_00487_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _05358_ (.A(_00344_),
    .B(_00311_),
    .Y(_00509_));
 sky130_fd_sc_hd__clkbuf_8 _05359_ (.A(net8),
    .X(_00520_));
 sky130_fd_sc_hd__nand2_1 _05360_ (.A(_00300_),
    .B(_00520_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _05361_ (.A(_00509_),
    .B(_00531_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _05362_ (.A(_00410_),
    .B(_00355_),
    .Y(_00553_));
 sky130_fd_sc_hd__inv_2 _05363_ (.A(_00553_),
    .Y(_00564_));
 sky130_fd_sc_hd__nor2_1 _05364_ (.A(_00509_),
    .B(_00531_),
    .Y(_00575_));
 sky130_fd_sc_hd__a21oi_2 _05365_ (.A1(_00542_),
    .A2(_00564_),
    .B1(_00575_),
    .Y(_00586_));
 sky130_fd_sc_hd__inv_2 _05366_ (.A(_00586_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _05367_ (.A(_00498_),
    .B(_00597_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand3_1 _05368_ (.A(_00586_),
    .B(_00443_),
    .C(_00487_),
    .Y(_00619_));
 sky130_fd_sc_hd__nand2_1 _05369_ (.A(_00608_),
    .B(_00619_),
    .Y(_00630_));
 sky130_fd_sc_hd__clkbuf_8 _05370_ (.A(net59),
    .X(_00641_));
 sky130_fd_sc_hd__nand2_1 _05371_ (.A(_00641_),
    .B(net8),
    .Y(_00652_));
 sky130_fd_sc_hd__inv_2 _05372_ (.A(_00652_),
    .Y(_00663_));
 sky130_fd_sc_hd__buf_8 _05373_ (.A(net33),
    .X(_00674_));
 sky130_fd_sc_hd__buf_6 _05374_ (.A(net13),
    .X(_00685_));
 sky130_fd_sc_hd__nand2_1 _05375_ (.A(_00674_),
    .B(_00685_),
    .Y(_00696_));
 sky130_fd_sc_hd__inv_2 _05376_ (.A(_00696_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand2_1 _05377_ (.A(_00663_),
    .B(_00707_),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_2 _05378_ (.A(_00652_),
    .B(_00696_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _05379_ (.A(_00718_),
    .B(_00729_),
    .Y(_00740_));
 sky130_fd_sc_hd__clkbuf_8 _05380_ (.A(net60),
    .X(_00751_));
 sky130_fd_sc_hd__nand2_1 _05381_ (.A(_00751_),
    .B(net7),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _05382_ (.A(_00740_),
    .B(_00762_),
    .Y(_00773_));
 sky130_fd_sc_hd__inv_2 _05383_ (.A(_00762_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand3_1 _05384_ (.A(_00718_),
    .B(_00784_),
    .C(_00729_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand2_1 _05385_ (.A(_00773_),
    .B(_00795_),
    .Y(_00806_));
 sky130_fd_sc_hd__inv_2 _05386_ (.A(_00806_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_1 _05387_ (.A(_00630_),
    .B(_00817_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand3_1 _05388_ (.A(_00608_),
    .B(_00619_),
    .C(_00806_),
    .Y(_00839_));
 sky130_fd_sc_hd__nand2_1 _05389_ (.A(_00828_),
    .B(_00839_),
    .Y(_00850_));
 sky130_fd_sc_hd__inv_2 _05390_ (.A(_00531_),
    .Y(_00861_));
 sky130_fd_sc_hd__nand2_1 _05391_ (.A(_00861_),
    .B(_00509_),
    .Y(_00872_));
 sky130_fd_sc_hd__inv_2 _05392_ (.A(_00509_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand2_1 _05393_ (.A(_00883_),
    .B(_00531_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand3_1 _05394_ (.A(_00872_),
    .B(_00894_),
    .C(_00553_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_1 _05395_ (.A(_00883_),
    .B(_00861_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand3_1 _05396_ (.A(_00916_),
    .B(_00564_),
    .C(_00542_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand2_1 _05397_ (.A(_00905_),
    .B(_00927_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _05398_ (.A(_00344_),
    .B(_00520_),
    .Y(_00949_));
 sky130_fd_sc_hd__clkbuf_8 _05399_ (.A(net7),
    .X(_00960_));
 sky130_fd_sc_hd__nand2_1 _05400_ (.A(_00300_),
    .B(_00960_),
    .Y(_00971_));
 sky130_fd_sc_hd__nand2_1 _05401_ (.A(_00949_),
    .B(_00971_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _05402_ (.A(_00410_),
    .B(net9),
    .Y(_00993_));
 sky130_fd_sc_hd__inv_2 _05403_ (.A(_00993_),
    .Y(_01004_));
 sky130_fd_sc_hd__nor2_1 _05404_ (.A(_00949_),
    .B(_00971_),
    .Y(_01015_));
 sky130_fd_sc_hd__a21oi_2 _05405_ (.A1(_00982_),
    .A2(_01004_),
    .B1(_01015_),
    .Y(_01026_));
 sky130_fd_sc_hd__nand2_1 _05406_ (.A(_00938_),
    .B(_01026_),
    .Y(_01037_));
 sky130_fd_sc_hd__nand2_1 _05407_ (.A(_00641_),
    .B(_00960_),
    .Y(_01048_));
 sky130_fd_sc_hd__inv_2 _05408_ (.A(_01048_),
    .Y(_01059_));
 sky130_fd_sc_hd__nand2_1 _05409_ (.A(_00674_),
    .B(_00421_),
    .Y(_01070_));
 sky130_fd_sc_hd__inv_2 _05410_ (.A(_01070_),
    .Y(_01081_));
 sky130_fd_sc_hd__nand2_1 _05411_ (.A(_01059_),
    .B(_01081_),
    .Y(_01092_));
 sky130_fd_sc_hd__nand2_1 _05412_ (.A(_01048_),
    .B(_01070_),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _05413_ (.A(_01092_),
    .B(_01103_),
    .Y(_01114_));
 sky130_fd_sc_hd__nand2_1 _05414_ (.A(_00751_),
    .B(net6),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _05415_ (.A(_01114_),
    .B(_01125_),
    .Y(_01136_));
 sky130_fd_sc_hd__inv_2 _05416_ (.A(_01125_),
    .Y(_01147_));
 sky130_fd_sc_hd__nand3_1 _05417_ (.A(_01092_),
    .B(_01147_),
    .C(_01103_),
    .Y(_01158_));
 sky130_fd_sc_hd__nand2_1 _05418_ (.A(_01136_),
    .B(_01158_),
    .Y(_01169_));
 sky130_fd_sc_hd__inv_2 _05419_ (.A(_01169_),
    .Y(_01180_));
 sky130_fd_sc_hd__nor2_1 _05420_ (.A(_01026_),
    .B(_00938_),
    .Y(_01191_));
 sky130_fd_sc_hd__a21oi_1 _05421_ (.A1(_01037_),
    .A2(_01180_),
    .B1(_01191_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _05422_ (.A(_00850_),
    .B(_01202_),
    .Y(_01213_));
 sky130_fd_sc_hd__clkbuf_8 _05423_ (.A(net62),
    .X(_01224_));
 sky130_fd_sc_hd__nand2_1 _05424_ (.A(_01224_),
    .B(net5),
    .Y(_01235_));
 sky130_fd_sc_hd__inv_2 _05425_ (.A(_01235_),
    .Y(_01246_));
 sky130_fd_sc_hd__buf_6 _05426_ (.A(net61),
    .X(_01257_));
 sky130_fd_sc_hd__nand2_1 _05427_ (.A(_01257_),
    .B(net6),
    .Y(_01268_));
 sky130_fd_sc_hd__inv_2 _05428_ (.A(_01268_),
    .Y(_01279_));
 sky130_fd_sc_hd__nand2_1 _05429_ (.A(_01246_),
    .B(_01279_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _05430_ (.A(_01235_),
    .B(_01268_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_1 _05431_ (.A(_01290_),
    .B(_01301_),
    .Y(_01312_));
 sky130_fd_sc_hd__buf_4 _05432_ (.A(net63),
    .X(_01323_));
 sky130_fd_sc_hd__buf_6 _05433_ (.A(net4),
    .X(_01334_));
 sky130_fd_sc_hd__nand2_1 _05434_ (.A(_01323_),
    .B(_01334_),
    .Y(_01345_));
 sky130_fd_sc_hd__nand2_1 _05435_ (.A(_01312_),
    .B(_01345_),
    .Y(_01356_));
 sky130_fd_sc_hd__inv_2 _05436_ (.A(_01345_),
    .Y(_01367_));
 sky130_fd_sc_hd__nand3_1 _05437_ (.A(_01290_),
    .B(_01367_),
    .C(_01301_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _05438_ (.A(_01356_),
    .B(_01378_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _05439_ (.A(_01048_),
    .B(_01070_),
    .Y(_01400_));
 sky130_fd_sc_hd__a21oi_2 _05440_ (.A1(_01103_),
    .A2(_01147_),
    .B1(_01400_),
    .Y(_01411_));
 sky130_fd_sc_hd__inv_2 _05441_ (.A(_01411_),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _05442_ (.A(_01389_),
    .B(_01422_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand3_1 _05443_ (.A(_01356_),
    .B(_01411_),
    .C(_01378_),
    .Y(_01444_));
 sky130_fd_sc_hd__nand2_1 _05444_ (.A(_01433_),
    .B(_01444_),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _05445_ (.A(_01257_),
    .B(net5),
    .Y(_01466_));
 sky130_fd_sc_hd__inv_2 _05446_ (.A(_01466_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_1 _05447_ (.A(_01224_),
    .B(net4),
    .Y(_01488_));
 sky130_fd_sc_hd__inv_2 _05448_ (.A(_01488_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_1 _05449_ (.A(_01477_),
    .B(_01499_),
    .Y(_01510_));
 sky130_fd_sc_hd__buf_6 _05450_ (.A(net3),
    .X(_01521_));
 sky130_fd_sc_hd__clkbuf_8 _05451_ (.A(_01521_),
    .X(_01532_));
 sky130_fd_sc_hd__nand2_1 _05452_ (.A(_01532_),
    .B(_01323_),
    .Y(_01543_));
 sky130_fd_sc_hd__inv_2 _05453_ (.A(_01543_),
    .Y(_01554_));
 sky130_fd_sc_hd__nand2_1 _05454_ (.A(_01466_),
    .B(_01488_),
    .Y(_01565_));
 sky130_fd_sc_hd__nand3_1 _05455_ (.A(_01510_),
    .B(_01554_),
    .C(_01565_),
    .Y(_01576_));
 sky130_fd_sc_hd__nand2_2 _05456_ (.A(_01576_),
    .B(_01510_),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _05457_ (.A(_01455_),
    .B(_01587_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand3b_1 _05458_ (.A_N(_01587_),
    .B(_01433_),
    .C(_01444_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_1 _05459_ (.A(_01598_),
    .B(_01609_),
    .Y(_01620_));
 sky130_fd_sc_hd__inv_2 _05460_ (.A(_01620_),
    .Y(_01631_));
 sky130_fd_sc_hd__nor2_1 _05461_ (.A(_01202_),
    .B(_00850_),
    .Y(_01642_));
 sky130_fd_sc_hd__a21o_1 _05462_ (.A1(_01213_),
    .A2(_01631_),
    .B1(_01642_),
    .X(_01653_));
 sky130_fd_sc_hd__nand2_1 _05463_ (.A(_00344_),
    .B(_00421_),
    .Y(_01664_));
 sky130_fd_sc_hd__inv_2 _05464_ (.A(_01664_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_1 _05465_ (.A(_00300_),
    .B(_00355_),
    .Y(_01686_));
 sky130_fd_sc_hd__nand2_1 _05466_ (.A(_01675_),
    .B(_01686_),
    .Y(_01697_));
 sky130_fd_sc_hd__inv_2 _05467_ (.A(_01686_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand2_1 _05468_ (.A(_01708_),
    .B(_01664_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _05469_ (.A(_00410_),
    .B(_00685_),
    .Y(_01730_));
 sky130_fd_sc_hd__nand3_1 _05470_ (.A(_01697_),
    .B(_01719_),
    .C(_01730_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _05471_ (.A(_01708_),
    .B(_01675_),
    .Y(_01752_));
 sky130_fd_sc_hd__inv_2 _05472_ (.A(_01730_),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _05473_ (.A(_01686_),
    .B(_01664_),
    .Y(_01774_));
 sky130_fd_sc_hd__nand3_1 _05474_ (.A(_01752_),
    .B(_01763_),
    .C(_01774_),
    .Y(_01785_));
 sky130_fd_sc_hd__nand2_1 _05475_ (.A(_01741_),
    .B(_01785_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _05476_ (.A(_00366_),
    .B(_00322_),
    .Y(_01807_));
 sky130_fd_sc_hd__a21oi_2 _05477_ (.A1(_00476_),
    .A2(_00465_),
    .B1(_01807_),
    .Y(_01818_));
 sky130_fd_sc_hd__inv_2 _05478_ (.A(_01818_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_1 _05479_ (.A(_01796_),
    .B(_01829_),
    .Y(_01840_));
 sky130_fd_sc_hd__nand3_1 _05480_ (.A(_01818_),
    .B(_01741_),
    .C(_01785_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _05481_ (.A(_01840_),
    .B(_01851_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_1 _05482_ (.A(_00641_),
    .B(_00311_),
    .Y(_01873_));
 sky130_fd_sc_hd__inv_2 _05483_ (.A(_01873_),
    .Y(_01884_));
 sky130_fd_sc_hd__clkbuf_4 _05484_ (.A(net14),
    .X(_01895_));
 sky130_fd_sc_hd__nand2_1 _05485_ (.A(_00674_),
    .B(_01895_),
    .Y(_01906_));
 sky130_fd_sc_hd__inv_2 _05486_ (.A(_01906_),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _05487_ (.A(_01884_),
    .B(_01917_),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _05488_ (.A(_01873_),
    .B(_01906_),
    .Y(_01939_));
 sky130_fd_sc_hd__nand2_1 _05489_ (.A(_01928_),
    .B(_01939_),
    .Y(_01950_));
 sky130_fd_sc_hd__nand2_1 _05490_ (.A(_00751_),
    .B(_00520_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_1 _05491_ (.A(_01950_),
    .B(_01961_),
    .Y(_01972_));
 sky130_fd_sc_hd__inv_2 _05492_ (.A(_01961_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand3_1 _05493_ (.A(_01928_),
    .B(_01983_),
    .C(_01939_),
    .Y(_01994_));
 sky130_fd_sc_hd__nand2_1 _05494_ (.A(_01972_),
    .B(_01994_),
    .Y(_02005_));
 sky130_fd_sc_hd__inv_2 _05495_ (.A(_02005_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_1 _05496_ (.A(_01862_),
    .B(_02016_),
    .Y(_02027_));
 sky130_fd_sc_hd__nand3_1 _05497_ (.A(_01840_),
    .B(_01851_),
    .C(_02005_),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _05498_ (.A(_02027_),
    .B(_02038_),
    .Y(_02049_));
 sky130_fd_sc_hd__inv_2 _05499_ (.A(_02049_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand2_1 _05500_ (.A(_00498_),
    .B(_00586_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_1 _05501_ (.A(_00586_),
    .B(_00498_),
    .Y(_02082_));
 sky130_fd_sc_hd__a21oi_4 _05502_ (.A1(_02071_),
    .A2(_00817_),
    .B1(_02082_),
    .Y(_02093_));
 sky130_fd_sc_hd__inv_2 _05503_ (.A(_02093_),
    .Y(_02104_));
 sky130_fd_sc_hd__nand2_1 _05504_ (.A(_02060_),
    .B(_02104_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _05505_ (.A(_01224_),
    .B(net6),
    .Y(_02126_));
 sky130_fd_sc_hd__inv_2 _05506_ (.A(_02126_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_1 _05507_ (.A(_01257_),
    .B(_00960_),
    .Y(_02148_));
 sky130_fd_sc_hd__inv_2 _05508_ (.A(_02148_),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_1 _05509_ (.A(_02137_),
    .B(_02159_),
    .Y(_02170_));
 sky130_fd_sc_hd__nand2_1 _05510_ (.A(_02126_),
    .B(_02148_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _05511_ (.A(_02170_),
    .B(_02181_),
    .Y(_02192_));
 sky130_fd_sc_hd__clkbuf_8 _05512_ (.A(_01323_),
    .X(_02203_));
 sky130_fd_sc_hd__clkbuf_8 _05513_ (.A(net5),
    .X(_02214_));
 sky130_fd_sc_hd__nand2_1 _05514_ (.A(_02203_),
    .B(_02214_),
    .Y(_02225_));
 sky130_fd_sc_hd__nand2_1 _05515_ (.A(_02192_),
    .B(_02225_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand3b_1 _05516_ (.A_N(_02225_),
    .B(_02170_),
    .C(_02181_),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _05517_ (.A(_02236_),
    .B(_02247_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _05518_ (.A(_00652_),
    .B(_00696_),
    .Y(_02269_));
 sky130_fd_sc_hd__a21oi_4 _05519_ (.A1(_00729_),
    .A2(_00784_),
    .B1(_02269_),
    .Y(_02280_));
 sky130_fd_sc_hd__inv_2 _05520_ (.A(_02280_),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_1 _05521_ (.A(_02258_),
    .B(_02291_),
    .Y(_02302_));
 sky130_fd_sc_hd__nand3_1 _05522_ (.A(_02236_),
    .B(_02247_),
    .C(_02280_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_1 _05523_ (.A(_02302_),
    .B(_02313_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_1 _05524_ (.A(_01378_),
    .B(_01290_),
    .Y(_02335_));
 sky130_fd_sc_hd__nand2_1 _05525_ (.A(_02324_),
    .B(_02335_),
    .Y(_02346_));
 sky130_fd_sc_hd__nand3b_1 _05526_ (.A_N(_02335_),
    .B(_02302_),
    .C(_02313_),
    .Y(_02357_));
 sky130_fd_sc_hd__nand2_1 _05527_ (.A(_02346_),
    .B(_02357_),
    .Y(_02368_));
 sky130_fd_sc_hd__inv_2 _05528_ (.A(_02368_),
    .Y(_02379_));
 sky130_fd_sc_hd__nand2_1 _05529_ (.A(_02049_),
    .B(_02093_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand3_1 _05530_ (.A(_02115_),
    .B(_02379_),
    .C(_02390_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand2_1 _05531_ (.A(_02060_),
    .B(_02093_),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _05532_ (.A(_02104_),
    .B(_02049_),
    .Y(_02423_));
 sky130_fd_sc_hd__nand3_1 _05533_ (.A(_02412_),
    .B(_02368_),
    .C(_02423_),
    .Y(_02434_));
 sky130_fd_sc_hd__nand3_1 _05534_ (.A(_01653_),
    .B(_02401_),
    .C(_02434_),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _05535_ (.A(_02401_),
    .B(_02434_),
    .Y(_02456_));
 sky130_fd_sc_hd__a21oi_2 _05536_ (.A1(_01213_),
    .A2(_01631_),
    .B1(_01642_),
    .Y(_02467_));
 sky130_fd_sc_hd__nand2_1 _05537_ (.A(_02456_),
    .B(_02467_),
    .Y(_02478_));
 sky130_fd_sc_hd__buf_6 _05538_ (.A(net2),
    .X(_02489_));
 sky130_fd_sc_hd__nand2_1 _05539_ (.A(_02489_),
    .B(net64),
    .Y(_02500_));
 sky130_fd_sc_hd__buf_6 _05540_ (.A(net32),
    .X(_02511_));
 sky130_fd_sc_hd__buf_6 _05541_ (.A(net34),
    .X(_02522_));
 sky130_fd_sc_hd__nand2_1 _05542_ (.A(_02511_),
    .B(_02522_),
    .Y(_02533_));
 sky130_fd_sc_hd__nand2_1 _05543_ (.A(_02500_),
    .B(_02533_),
    .Y(_02544_));
 sky130_fd_sc_hd__buf_6 _05544_ (.A(net31),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _05545_ (.A(_02555_),
    .B(net35),
    .Y(_02566_));
 sky130_fd_sc_hd__inv_2 _05546_ (.A(_02566_),
    .Y(_02577_));
 sky130_fd_sc_hd__nor2_1 _05547_ (.A(_02500_),
    .B(_02533_),
    .Y(_02588_));
 sky130_fd_sc_hd__a21oi_2 _05548_ (.A1(_02544_),
    .A2(_02577_),
    .B1(_02588_),
    .Y(_02599_));
 sky130_fd_sc_hd__nand2_1 _05549_ (.A(_02489_),
    .B(_02522_),
    .Y(_02610_));
 sky130_fd_sc_hd__inv_2 _05550_ (.A(_02610_),
    .Y(_02621_));
 sky130_fd_sc_hd__nand2_1 _05551_ (.A(_01521_),
    .B(net64),
    .Y(_02632_));
 sky130_fd_sc_hd__inv_2 _05552_ (.A(_02632_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _05553_ (.A(_02621_),
    .B(_02643_),
    .Y(_02654_));
 sky130_fd_sc_hd__nand2_1 _05554_ (.A(_02610_),
    .B(_02632_),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _05555_ (.A(_02654_),
    .B(_02665_),
    .Y(_02676_));
 sky130_fd_sc_hd__clkbuf_8 _05556_ (.A(net35),
    .X(_02687_));
 sky130_fd_sc_hd__nand2_1 _05557_ (.A(_02511_),
    .B(_02687_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_1 _05558_ (.A(_02676_),
    .B(_02698_),
    .Y(_02709_));
 sky130_fd_sc_hd__inv_2 _05559_ (.A(_02698_),
    .Y(_02720_));
 sky130_fd_sc_hd__nand3_1 _05560_ (.A(_02654_),
    .B(_02720_),
    .C(_02665_),
    .Y(_02731_));
 sky130_fd_sc_hd__nand2_1 _05561_ (.A(_02709_),
    .B(_02731_),
    .Y(_02742_));
 sky130_fd_sc_hd__inv_2 _05562_ (.A(_02599_),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _05563_ (.A(_02742_),
    .B(_02753_),
    .Y(_02764_));
 sky130_fd_sc_hd__nand3_1 _05564_ (.A(_02709_),
    .B(_02599_),
    .C(_02731_),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2_1 _05565_ (.A(_02764_),
    .B(_02775_),
    .Y(_02786_));
 sky130_fd_sc_hd__clkbuf_8 _05566_ (.A(net30),
    .X(_02797_));
 sky130_fd_sc_hd__nand2_1 _05567_ (.A(_02797_),
    .B(net37),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _05568_ (.A(_02555_),
    .B(net36),
    .Y(_02819_));
 sky130_fd_sc_hd__nor2_1 _05569_ (.A(_02808_),
    .B(_02819_),
    .Y(_02830_));
 sky130_fd_sc_hd__inv_2 _05570_ (.A(_02830_),
    .Y(_02841_));
 sky130_fd_sc_hd__nand2_1 _05571_ (.A(_02808_),
    .B(_02819_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand2_1 _05572_ (.A(_02841_),
    .B(_02852_),
    .Y(_02863_));
 sky130_fd_sc_hd__buf_6 _05573_ (.A(net29),
    .X(_02874_));
 sky130_fd_sc_hd__nand2_1 _05574_ (.A(_02874_),
    .B(net38),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_1 _05575_ (.A(_02863_),
    .B(_02885_),
    .Y(_02896_));
 sky130_fd_sc_hd__inv_2 _05576_ (.A(_02885_),
    .Y(_02907_));
 sky130_fd_sc_hd__nand3_1 _05577_ (.A(_02841_),
    .B(_02907_),
    .C(_02852_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand2_1 _05578_ (.A(_02896_),
    .B(_02918_),
    .Y(_02929_));
 sky130_fd_sc_hd__inv_2 _05579_ (.A(_02929_),
    .Y(_02940_));
 sky130_fd_sc_hd__nand2_1 _05580_ (.A(_02786_),
    .B(_02940_),
    .Y(_02951_));
 sky130_fd_sc_hd__o21ai_2 _05581_ (.A1(_02599_),
    .A2(_02742_),
    .B1(_02951_),
    .Y(_02962_));
 sky130_fd_sc_hd__nand2_1 _05582_ (.A(_01389_),
    .B(_01411_),
    .Y(_02973_));
 sky130_fd_sc_hd__nor2_1 _05583_ (.A(_01411_),
    .B(_01389_),
    .Y(_02984_));
 sky130_fd_sc_hd__a21oi_4 _05584_ (.A1(_02973_),
    .A2(_01587_),
    .B1(_02984_),
    .Y(_02995_));
 sky130_fd_sc_hd__inv_2 _05585_ (.A(_02995_),
    .Y(_03006_));
 sky130_fd_sc_hd__nand2_1 _05586_ (.A(_01532_),
    .B(_02522_),
    .Y(_03017_));
 sky130_fd_sc_hd__inv_2 _05587_ (.A(_03017_),
    .Y(_03028_));
 sky130_fd_sc_hd__clkbuf_8 _05588_ (.A(net64),
    .X(_03039_));
 sky130_fd_sc_hd__nand2_1 _05589_ (.A(_03039_),
    .B(net4),
    .Y(_03050_));
 sky130_fd_sc_hd__inv_2 _05590_ (.A(_03050_),
    .Y(_03061_));
 sky130_fd_sc_hd__nand2_1 _05591_ (.A(_03028_),
    .B(_03061_),
    .Y(_03072_));
 sky130_fd_sc_hd__nand2_1 _05592_ (.A(_03017_),
    .B(_03050_),
    .Y(_03083_));
 sky130_fd_sc_hd__nand2_1 _05593_ (.A(_03072_),
    .B(_03083_),
    .Y(_03094_));
 sky130_fd_sc_hd__clkbuf_8 _05594_ (.A(_02489_),
    .X(_03105_));
 sky130_fd_sc_hd__nand2_1 _05595_ (.A(_03105_),
    .B(_02687_),
    .Y(_03116_));
 sky130_fd_sc_hd__nand2_1 _05596_ (.A(_03094_),
    .B(_03116_),
    .Y(_03127_));
 sky130_fd_sc_hd__inv_2 _05597_ (.A(_03116_),
    .Y(_03138_));
 sky130_fd_sc_hd__nand3_1 _05598_ (.A(_03072_),
    .B(_03138_),
    .C(_03083_),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _05599_ (.A(_03127_),
    .B(_03149_),
    .Y(_03160_));
 sky130_fd_sc_hd__nor2_1 _05600_ (.A(_02610_),
    .B(_02632_),
    .Y(_03171_));
 sky130_fd_sc_hd__a21oi_2 _05601_ (.A1(_02665_),
    .A2(_02720_),
    .B1(_03171_),
    .Y(_03182_));
 sky130_fd_sc_hd__inv_2 _05602_ (.A(_03182_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2_1 _05603_ (.A(_03160_),
    .B(_03193_),
    .Y(_03204_));
 sky130_fd_sc_hd__nand3_1 _05604_ (.A(_03127_),
    .B(_03182_),
    .C(_03149_),
    .Y(_03215_));
 sky130_fd_sc_hd__nand2_1 _05605_ (.A(_03204_),
    .B(_03215_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand2_1 _05606_ (.A(_02555_),
    .B(net37),
    .Y(_03237_));
 sky130_fd_sc_hd__clkbuf_8 _05607_ (.A(net36),
    .X(_03248_));
 sky130_fd_sc_hd__nand2_1 _05608_ (.A(_02511_),
    .B(_03248_),
    .Y(_03259_));
 sky130_fd_sc_hd__nor2_1 _05609_ (.A(_03237_),
    .B(_03259_),
    .Y(_03270_));
 sky130_fd_sc_hd__inv_2 _05610_ (.A(_03270_),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_1 _05611_ (.A(_03237_),
    .B(_03259_),
    .Y(_03292_));
 sky130_fd_sc_hd__nand2_1 _05612_ (.A(_03281_),
    .B(_03292_),
    .Y(_03303_));
 sky130_fd_sc_hd__nand2_1 _05613_ (.A(_02797_),
    .B(net38),
    .Y(_03314_));
 sky130_fd_sc_hd__nand2_1 _05614_ (.A(_03303_),
    .B(_03314_),
    .Y(_03325_));
 sky130_fd_sc_hd__inv_2 _05615_ (.A(_03314_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand3_1 _05616_ (.A(_03281_),
    .B(_03336_),
    .C(_03292_),
    .Y(_03347_));
 sky130_fd_sc_hd__nand2_1 _05617_ (.A(_03325_),
    .B(_03347_),
    .Y(_03358_));
 sky130_fd_sc_hd__inv_2 _05618_ (.A(_03358_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand2_1 _05619_ (.A(_03226_),
    .B(_03369_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand3_1 _05620_ (.A(_03204_),
    .B(_03215_),
    .C(_03358_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand2_1 _05621_ (.A(_03380_),
    .B(_03391_),
    .Y(_03402_));
 sky130_fd_sc_hd__nand2_1 _05622_ (.A(_03006_),
    .B(_03402_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand3_1 _05623_ (.A(_02995_),
    .B(_03380_),
    .C(_03391_),
    .Y(_03424_));
 sky130_fd_sc_hd__nand3b_1 _05624_ (.A_N(_02962_),
    .B(_03413_),
    .C(_03424_),
    .Y(_03435_));
 sky130_fd_sc_hd__nand2_1 _05625_ (.A(_03413_),
    .B(_03424_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _05626_ (.A(_03446_),
    .B(_02962_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_1 _05627_ (.A(_03435_),
    .B(_03457_),
    .Y(_03468_));
 sky130_fd_sc_hd__inv_2 _05628_ (.A(_03468_),
    .Y(_03479_));
 sky130_fd_sc_hd__nand3_2 _05629_ (.A(_02445_),
    .B(_02478_),
    .C(_03479_),
    .Y(_03490_));
 sky130_fd_sc_hd__nand2_1 _05630_ (.A(_02456_),
    .B(_01653_),
    .Y(_03501_));
 sky130_fd_sc_hd__nand3_1 _05631_ (.A(_02467_),
    .B(_02401_),
    .C(_02434_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand3_1 _05632_ (.A(_03501_),
    .B(_03512_),
    .C(_03468_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _05633_ (.A(_03490_),
    .B(_03523_),
    .Y(_03534_));
 sky130_fd_sc_hd__nand3_1 _05634_ (.A(_01202_),
    .B(_00828_),
    .C(_00839_),
    .Y(_03545_));
 sky130_fd_sc_hd__a21o_1 _05635_ (.A1(_01037_),
    .A2(_01180_),
    .B1(_01191_),
    .X(_03556_));
 sky130_fd_sc_hd__nand2_1 _05636_ (.A(_03556_),
    .B(_00850_),
    .Y(_03567_));
 sky130_fd_sc_hd__nand2_1 _05637_ (.A(_03545_),
    .B(_03567_),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_1 _05638_ (.A(_03578_),
    .B(_01631_),
    .Y(_03589_));
 sky130_fd_sc_hd__nand3_1 _05639_ (.A(_03545_),
    .B(_03567_),
    .C(_01620_),
    .Y(_03600_));
 sky130_fd_sc_hd__nand2_2 _05640_ (.A(_03589_),
    .B(_03600_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand2_1 _05641_ (.A(_00751_),
    .B(net5),
    .Y(_03622_));
 sky130_fd_sc_hd__clkinvlp_2 _05642_ (.A(_03622_),
    .Y(_03633_));
 sky130_fd_sc_hd__nand2_1 _05643_ (.A(_00641_),
    .B(net6),
    .Y(_03644_));
 sky130_fd_sc_hd__nand2_1 _05644_ (.A(_00674_),
    .B(_00355_),
    .Y(_03655_));
 sky130_fd_sc_hd__nand2_1 _05645_ (.A(_03644_),
    .B(_03655_),
    .Y(_03666_));
 sky130_fd_sc_hd__inv_2 _05646_ (.A(_03644_),
    .Y(_03677_));
 sky130_fd_sc_hd__inv_2 _05647_ (.A(_03655_),
    .Y(_03688_));
 sky130_fd_sc_hd__nand2_1 _05648_ (.A(_03677_),
    .B(_03688_),
    .Y(_03699_));
 sky130_fd_sc_hd__a21boi_1 _05649_ (.A1(_03633_),
    .A2(_03666_),
    .B1_N(_03699_),
    .Y(_03710_));
 sky130_fd_sc_hd__nand2_1 _05650_ (.A(_01510_),
    .B(_01565_),
    .Y(_03721_));
 sky130_fd_sc_hd__nand2_1 _05651_ (.A(_03721_),
    .B(_01543_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand3_1 _05652_ (.A(_03710_),
    .B(_01576_),
    .C(_03732_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand2_1 _05653_ (.A(_03732_),
    .B(_01576_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand3_1 _05654_ (.A(_03699_),
    .B(_03633_),
    .C(_03666_),
    .Y(_03765_));
 sky130_fd_sc_hd__nand2_1 _05655_ (.A(_03765_),
    .B(_03699_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand2_1 _05656_ (.A(_03754_),
    .B(_03776_),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _05657_ (.A(_03743_),
    .B(_03787_),
    .Y(_03798_));
 sky130_fd_sc_hd__nand2_1 _05658_ (.A(_02489_),
    .B(_01323_),
    .Y(_03809_));
 sky130_fd_sc_hd__nand2_1 _05659_ (.A(_01257_),
    .B(net4),
    .Y(_03820_));
 sky130_fd_sc_hd__inv_2 _05660_ (.A(_03820_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_1 _05661_ (.A(_01521_),
    .B(_01224_),
    .Y(_03842_));
 sky130_fd_sc_hd__inv_2 _05662_ (.A(_03842_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_1 _05663_ (.A(_03831_),
    .B(_03853_),
    .Y(_03864_));
 sky130_fd_sc_hd__nand2_1 _05664_ (.A(_03820_),
    .B(_03842_),
    .Y(_03875_));
 sky130_fd_sc_hd__nand3b_2 _05665_ (.A_N(_03809_),
    .B(_03864_),
    .C(_03875_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand2_2 _05666_ (.A(_03886_),
    .B(_03864_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_1 _05667_ (.A(_03798_),
    .B(_03897_),
    .Y(_03908_));
 sky130_fd_sc_hd__nand3b_1 _05668_ (.A_N(_03897_),
    .B(_03743_),
    .C(_03787_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _05669_ (.A(_03908_),
    .B(_03919_),
    .Y(_03930_));
 sky130_fd_sc_hd__inv_2 _05670_ (.A(_03930_),
    .Y(_03941_));
 sky130_fd_sc_hd__inv_2 _05671_ (.A(_01026_),
    .Y(_03952_));
 sky130_fd_sc_hd__nand2_1 _05672_ (.A(_00938_),
    .B(_03952_),
    .Y(_03963_));
 sky130_fd_sc_hd__nand3_1 _05673_ (.A(_01026_),
    .B(_00905_),
    .C(_00927_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _05674_ (.A(_03963_),
    .B(_03974_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _05675_ (.A(_03985_),
    .B(_01180_),
    .Y(_03996_));
 sky130_fd_sc_hd__nand3_1 _05676_ (.A(_03963_),
    .B(_03974_),
    .C(_01169_),
    .Y(_04007_));
 sky130_fd_sc_hd__nand2_1 _05677_ (.A(_03996_),
    .B(_04007_),
    .Y(_04018_));
 sky130_fd_sc_hd__inv_2 _05678_ (.A(_00971_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _05679_ (.A(_04029_),
    .B(_00949_),
    .Y(_04040_));
 sky130_fd_sc_hd__inv_2 _05680_ (.A(_00949_),
    .Y(_04051_));
 sky130_fd_sc_hd__nand2_1 _05681_ (.A(_04051_),
    .B(_00971_),
    .Y(_04062_));
 sky130_fd_sc_hd__nand3_1 _05682_ (.A(_04040_),
    .B(_04062_),
    .C(_00993_),
    .Y(_04073_));
 sky130_fd_sc_hd__nand2_1 _05683_ (.A(_04051_),
    .B(_04029_),
    .Y(_04084_));
 sky130_fd_sc_hd__nand3_1 _05684_ (.A(_04084_),
    .B(_01004_),
    .C(_00982_),
    .Y(_04095_));
 sky130_fd_sc_hd__nand2_1 _05685_ (.A(_04073_),
    .B(_04095_),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_1 _05686_ (.A(_00344_),
    .B(_00960_),
    .Y(_04117_));
 sky130_fd_sc_hd__clkbuf_8 _05687_ (.A(net6),
    .X(_04128_));
 sky130_fd_sc_hd__nand2_1 _05688_ (.A(_00300_),
    .B(_04128_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _05689_ (.A(_04117_),
    .B(_04139_),
    .Y(_04150_));
 sky130_fd_sc_hd__nand2_1 _05690_ (.A(_00410_),
    .B(net8),
    .Y(_04161_));
 sky130_fd_sc_hd__inv_2 _05691_ (.A(_04161_),
    .Y(_04172_));
 sky130_fd_sc_hd__nor2_1 _05692_ (.A(_04117_),
    .B(_04139_),
    .Y(_04183_));
 sky130_fd_sc_hd__a21oi_2 _05693_ (.A1(_04150_),
    .A2(_04172_),
    .B1(_04183_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _05694_ (.A(_04106_),
    .B(_04194_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand2_1 _05695_ (.A(_03699_),
    .B(_03666_),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_1 _05696_ (.A(_04216_),
    .B(_03622_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand2_1 _05697_ (.A(_04227_),
    .B(_03765_),
    .Y(_04238_));
 sky130_fd_sc_hd__clkinvlp_2 _05698_ (.A(_04238_),
    .Y(_04249_));
 sky130_fd_sc_hd__nor2_1 _05699_ (.A(_04194_),
    .B(_04106_),
    .Y(_04260_));
 sky130_fd_sc_hd__a21oi_1 _05700_ (.A1(_04205_),
    .A2(_04249_),
    .B1(_04260_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand2_1 _05701_ (.A(_04018_),
    .B(_04271_),
    .Y(_04282_));
 sky130_fd_sc_hd__nor2_1 _05702_ (.A(_04271_),
    .B(_04018_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21oi_4 _05703_ (.A1(_03941_),
    .A2(_04282_),
    .B1(_04293_),
    .Y(_04304_));
 sky130_fd_sc_hd__nand2_1 _05704_ (.A(_03611_),
    .B(_04304_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _05705_ (.A(_03754_),
    .B(_03710_),
    .Y(_04326_));
 sky130_fd_sc_hd__nor2_1 _05706_ (.A(_03710_),
    .B(_03754_),
    .Y(_04337_));
 sky130_fd_sc_hd__a21oi_4 _05707_ (.A1(_04326_),
    .A2(_03897_),
    .B1(_04337_),
    .Y(_04348_));
 sky130_fd_sc_hd__inv_2 _05708_ (.A(_04348_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand3_1 _05709_ (.A(_02764_),
    .B(_02775_),
    .C(_02929_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_1 _05710_ (.A(_02951_),
    .B(_04370_),
    .Y(_04381_));
 sky130_fd_sc_hd__nand2_1 _05711_ (.A(_04359_),
    .B(_04381_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand3_1 _05712_ (.A(_04348_),
    .B(_02951_),
    .C(_04370_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_1 _05713_ (.A(_04392_),
    .B(_04403_),
    .Y(_04414_));
 sky130_fd_sc_hd__inv_2 _05714_ (.A(_02544_),
    .Y(_04425_));
 sky130_fd_sc_hd__o21ai_1 _05715_ (.A1(_02588_),
    .A2(_04425_),
    .B1(_02566_),
    .Y(_04436_));
 sky130_fd_sc_hd__nand3b_1 _05716_ (.A_N(_02588_),
    .B(_02577_),
    .C(_02544_),
    .Y(_04447_));
 sky130_fd_sc_hd__nand2_1 _05717_ (.A(_04436_),
    .B(_04447_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand2_1 _05718_ (.A(_02555_),
    .B(_02522_),
    .Y(_04469_));
 sky130_fd_sc_hd__nand2_1 _05719_ (.A(_02511_),
    .B(net64),
    .Y(_04480_));
 sky130_fd_sc_hd__nand2_1 _05720_ (.A(_04469_),
    .B(_04480_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand2_1 _05721_ (.A(_02797_),
    .B(net35),
    .Y(_04502_));
 sky130_fd_sc_hd__inv_2 _05722_ (.A(_04502_),
    .Y(_04513_));
 sky130_fd_sc_hd__nor2_1 _05723_ (.A(_04469_),
    .B(_04480_),
    .Y(_04524_));
 sky130_fd_sc_hd__a21oi_2 _05724_ (.A1(_04491_),
    .A2(_04513_),
    .B1(_04524_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2_1 _05725_ (.A(_04458_),
    .B(_04535_),
    .Y(_04546_));
 sky130_fd_sc_hd__inv_2 _05726_ (.A(_04535_),
    .Y(_04557_));
 sky130_fd_sc_hd__nand3_1 _05727_ (.A(_04447_),
    .B(_04436_),
    .C(_04557_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand2_1 _05728_ (.A(_02874_),
    .B(net37),
    .Y(_04579_));
 sky130_fd_sc_hd__nand2_1 _05729_ (.A(_02797_),
    .B(net36),
    .Y(_04590_));
 sky130_fd_sc_hd__nor2_1 _05730_ (.A(_04579_),
    .B(_04590_),
    .Y(_04601_));
 sky130_fd_sc_hd__nand2_1 _05731_ (.A(_04579_),
    .B(_04590_),
    .Y(_04612_));
 sky130_fd_sc_hd__inv_2 _05732_ (.A(_04612_),
    .Y(_04623_));
 sky130_fd_sc_hd__buf_6 _05733_ (.A(net28),
    .X(_04634_));
 sky130_fd_sc_hd__clkbuf_8 _05734_ (.A(net38),
    .X(_04645_));
 sky130_fd_sc_hd__nand2_1 _05735_ (.A(_04634_),
    .B(_04645_),
    .Y(_04656_));
 sky130_fd_sc_hd__o21ai_1 _05736_ (.A1(_04601_),
    .A2(_04623_),
    .B1(_04656_),
    .Y(_04667_));
 sky130_fd_sc_hd__inv_2 _05737_ (.A(_04656_),
    .Y(_04678_));
 sky130_fd_sc_hd__nand3b_1 _05738_ (.A_N(_04601_),
    .B(_04678_),
    .C(_04612_),
    .Y(_04689_));
 sky130_fd_sc_hd__nand2_1 _05739_ (.A(_04667_),
    .B(_04689_),
    .Y(_04700_));
 sky130_fd_sc_hd__inv_2 _05740_ (.A(_04700_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand3_1 _05741_ (.A(_04546_),
    .B(_04568_),
    .C(_04711_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _05742_ (.A(_04722_),
    .B(_04568_),
    .Y(_04733_));
 sky130_fd_sc_hd__nand2_1 _05743_ (.A(_04414_),
    .B(_04733_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand3b_1 _05744_ (.A_N(_04733_),
    .B(_04392_),
    .C(_04403_),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _05745_ (.A(_04744_),
    .B(_04755_),
    .Y(_04766_));
 sky130_fd_sc_hd__inv_2 _05746_ (.A(_04766_),
    .Y(_04776_));
 sky130_fd_sc_hd__nor2_1 _05747_ (.A(_04304_),
    .B(_03611_),
    .Y(_04785_));
 sky130_fd_sc_hd__a21oi_1 _05748_ (.A1(_04315_),
    .A2(_04776_),
    .B1(_04785_),
    .Y(_04796_));
 sky130_fd_sc_hd__nand2_1 _05749_ (.A(_03534_),
    .B(_04796_),
    .Y(_04805_));
 sky130_fd_sc_hd__buf_12 _05750_ (.A(net27),
    .X(_04814_));
 sky130_fd_sc_hd__nand2_1 _05751_ (.A(_04814_),
    .B(net40),
    .Y(_04823_));
 sky130_fd_sc_hd__inv_2 _05752_ (.A(_04823_),
    .Y(_04832_));
 sky130_fd_sc_hd__nand2_1 _05753_ (.A(_04634_),
    .B(net39),
    .Y(_04839_));
 sky130_fd_sc_hd__inv_2 _05754_ (.A(_04839_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _05755_ (.A(_04832_),
    .B(_04847_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_1 _05756_ (.A(_04823_),
    .B(_04839_),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_1 _05757_ (.A(_04855_),
    .B(_04864_),
    .Y(_04872_));
 sky130_fd_sc_hd__buf_12 _05758_ (.A(net26),
    .X(_04880_));
 sky130_fd_sc_hd__clkbuf_8 _05759_ (.A(net41),
    .X(_04888_));
 sky130_fd_sc_hd__nand2_1 _05760_ (.A(_04880_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__nand2_1 _05761_ (.A(_04872_),
    .B(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand3b_1 _05762_ (.A_N(_04889_),
    .B(_04855_),
    .C(_04864_),
    .Y(_04891_));
 sky130_fd_sc_hd__nand2_1 _05763_ (.A(_04890_),
    .B(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21oi_2 _05764_ (.A1(_04612_),
    .A2(_04678_),
    .B1(_04601_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand2_1 _05765_ (.A(_04892_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__buf_6 _05766_ (.A(net23),
    .X(_04895_));
 sky130_fd_sc_hd__nand2_1 _05767_ (.A(_04895_),
    .B(_04888_),
    .Y(_04896_));
 sky130_fd_sc_hd__clkbuf_8 _05768_ (.A(net39),
    .X(_04897_));
 sky130_fd_sc_hd__nand2_1 _05769_ (.A(_04814_),
    .B(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__clkbuf_8 _05770_ (.A(net40),
    .X(_04899_));
 sky130_fd_sc_hd__nand2_1 _05771_ (.A(_04880_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__or2_1 _05772_ (.A(_04898_),
    .B(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__nand2_1 _05773_ (.A(_04898_),
    .B(_04900_),
    .Y(_04902_));
 sky130_fd_sc_hd__nand3b_1 _05774_ (.A_N(_04896_),
    .B(_04901_),
    .C(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__nand2_1 _05775_ (.A(_04903_),
    .B(_04901_),
    .Y(_04904_));
 sky130_fd_sc_hd__nor2_1 _05776_ (.A(_04893_),
    .B(_04892_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21oi_2 _05777_ (.A1(_04894_),
    .A2(_04904_),
    .B1(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__a21oi_2 _05778_ (.A1(_02852_),
    .A2(_02907_),
    .B1(_02830_),
    .Y(_04907_));
 sky130_fd_sc_hd__inv_2 _05779_ (.A(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand2_1 _05780_ (.A(_04814_),
    .B(_04888_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand2_1 _05781_ (.A(_04634_),
    .B(net40),
    .Y(_04910_));
 sky130_fd_sc_hd__inv_2 _05782_ (.A(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__nand2_1 _05783_ (.A(_02874_),
    .B(net39),
    .Y(_04912_));
 sky130_fd_sc_hd__inv_2 _05784_ (.A(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__nand2_1 _05785_ (.A(_04911_),
    .B(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_1 _05786_ (.A(_04910_),
    .B(_04912_),
    .Y(_04915_));
 sky130_fd_sc_hd__nand3b_2 _05787_ (.A_N(_04909_),
    .B(_04914_),
    .C(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__nand2_1 _05788_ (.A(_04914_),
    .B(_04915_),
    .Y(_04917_));
 sky130_fd_sc_hd__nand2_1 _05789_ (.A(_04917_),
    .B(_04909_),
    .Y(_04918_));
 sky130_fd_sc_hd__nand3_1 _05790_ (.A(_04908_),
    .B(_04916_),
    .C(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__nand2_1 _05791_ (.A(_04918_),
    .B(_04916_),
    .Y(_04920_));
 sky130_fd_sc_hd__nand2_1 _05792_ (.A(_04920_),
    .B(_04907_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_1 _05793_ (.A(_04891_),
    .B(_04855_),
    .Y(_04922_));
 sky130_fd_sc_hd__nand3_1 _05794_ (.A(_04919_),
    .B(_04921_),
    .C(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _05795_ (.A(_04920_),
    .B(_04908_),
    .Y(_04924_));
 sky130_fd_sc_hd__nand3_1 _05796_ (.A(_04918_),
    .B(_04916_),
    .C(_04907_),
    .Y(_04925_));
 sky130_fd_sc_hd__inv_2 _05797_ (.A(_04922_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand3_1 _05798_ (.A(_04924_),
    .B(_04925_),
    .C(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand3_1 _05799_ (.A(_04906_),
    .B(_04923_),
    .C(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__inv_2 _05800_ (.A(_04906_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _05801_ (.A(_04923_),
    .B(_04927_),
    .Y(_04930_));
 sky130_fd_sc_hd__nand2_1 _05802_ (.A(_04929_),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand2_1 _05803_ (.A(_04928_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__buf_4 _05804_ (.A(net43),
    .X(_04933_));
 sky130_fd_sc_hd__nand2_1 _05805_ (.A(_04895_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__inv_2 _05806_ (.A(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__buf_4 _05807_ (.A(net42),
    .X(_04936_));
 sky130_fd_sc_hd__nand2_1 _05808_ (.A(_04880_),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__inv_2 _05809_ (.A(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_1 _05810_ (.A(_04935_),
    .B(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _05811_ (.A(_04934_),
    .B(_04937_),
    .Y(_04940_));
 sky130_fd_sc_hd__buf_4 _05812_ (.A(net45),
    .X(_04941_));
 sky130_fd_sc_hd__nand2_1 _05813_ (.A(net12),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__inv_2 _05814_ (.A(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__a21o_1 _05815_ (.A1(_04939_),
    .A2(_04940_),
    .B1(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__nand3_1 _05816_ (.A(_04939_),
    .B(_04943_),
    .C(_04940_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _05817_ (.A(_04944_),
    .B(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__buf_6 _05818_ (.A(net12),
    .X(_04947_));
 sky130_fd_sc_hd__nand2_1 _05819_ (.A(_04947_),
    .B(_04933_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_1 _05820_ (.A(_04895_),
    .B(_04936_),
    .Y(_04949_));
 sky130_fd_sc_hd__nand2_1 _05821_ (.A(_04948_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nand2_1 _05822_ (.A(net1),
    .B(_04941_),
    .Y(_04951_));
 sky130_fd_sc_hd__inv_2 _05823_ (.A(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__nor2_1 _05824_ (.A(_04948_),
    .B(_04949_),
    .Y(_04953_));
 sky130_fd_sc_hd__a21oi_1 _05825_ (.A1(_04950_),
    .A2(_04952_),
    .B1(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _05826_ (.A(_04946_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand3b_1 _05827_ (.A_N(_04954_),
    .B(_04944_),
    .C(_04945_),
    .Y(_04956_));
 sky130_fd_sc_hd__nand2_1 _05828_ (.A(_04955_),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__buf_6 _05829_ (.A(net1),
    .X(_04958_));
 sky130_fd_sc_hd__nand2_1 _05830_ (.A(net46),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__nand2_1 _05831_ (.A(_04957_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand3b_1 _05832_ (.A_N(_04959_),
    .B(_04955_),
    .C(_04956_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand2_1 _05833_ (.A(_04960_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__inv_2 _05834_ (.A(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__nand2_1 _05835_ (.A(_04932_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand3_1 _05836_ (.A(_04928_),
    .B(_04931_),
    .C(_04962_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_1 _05837_ (.A(_04964_),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__nand2_1 _05838_ (.A(_04381_),
    .B(_04348_),
    .Y(_04967_));
 sky130_fd_sc_hd__nor2_1 _05839_ (.A(_04348_),
    .B(_04381_),
    .Y(_04968_));
 sky130_fd_sc_hd__a21oi_2 _05840_ (.A1(_04967_),
    .A2(_04733_),
    .B1(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__inv_2 _05841_ (.A(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__nand2_1 _05842_ (.A(_04966_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand3_1 _05843_ (.A(_04969_),
    .B(_04964_),
    .C(_04965_),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_1 _05844_ (.A(_04971_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__and4_1 _05845_ (.A(_04947_),
    .B(net1),
    .C(_04936_),
    .D(_04933_),
    .X(_04974_));
 sky130_fd_sc_hd__inv_2 _05846_ (.A(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__nor2b_1 _05847_ (.A(_04953_),
    .B_N(_04950_),
    .Y(_04976_));
 sky130_fd_sc_hd__xor2_1 _05848_ (.A(_04951_),
    .B(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__or2_1 _05849_ (.A(_04975_),
    .B(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__nand2_1 _05850_ (.A(_04977_),
    .B(_04975_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _05851_ (.A(_04978_),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__inv_2 _05852_ (.A(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand3_1 _05853_ (.A(_04890_),
    .B(_04893_),
    .C(_04891_),
    .Y(_04982_));
 sky130_fd_sc_hd__inv_2 _05854_ (.A(_04893_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_1 _05855_ (.A(_04892_),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__nand3b_1 _05856_ (.A_N(_04904_),
    .B(_04982_),
    .C(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_1 _05857_ (.A(_04984_),
    .B(_04982_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_1 _05858_ (.A(_04986_),
    .B(_04904_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand2_1 _05859_ (.A(_04985_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand2_1 _05860_ (.A(_04901_),
    .B(_04902_),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_1 _05861_ (.A(_04989_),
    .B(_04896_),
    .Y(_04990_));
 sky130_fd_sc_hd__nand2_1 _05862_ (.A(_04990_),
    .B(_04903_),
    .Y(_04991_));
 sky130_fd_sc_hd__nand2_1 _05863_ (.A(_04634_),
    .B(net37),
    .Y(_04992_));
 sky130_fd_sc_hd__nand2_1 _05864_ (.A(_02874_),
    .B(_03248_),
    .Y(_04993_));
 sky130_fd_sc_hd__nand2_1 _05865_ (.A(_04992_),
    .B(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nand2_1 _05866_ (.A(_04814_),
    .B(_04645_),
    .Y(_04995_));
 sky130_fd_sc_hd__inv_2 _05867_ (.A(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nor2_1 _05868_ (.A(_04992_),
    .B(_04993_),
    .Y(_04997_));
 sky130_fd_sc_hd__a21oi_2 _05869_ (.A1(_04994_),
    .A2(_04996_),
    .B1(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__nand2_1 _05870_ (.A(_04991_),
    .B(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__nand2_1 _05871_ (.A(_04947_),
    .B(_04888_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _05872_ (.A(_04880_),
    .B(_04897_),
    .Y(_05001_));
 sky130_fd_sc_hd__inv_2 _05873_ (.A(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__nand2_1 _05874_ (.A(_04895_),
    .B(net40),
    .Y(_05003_));
 sky130_fd_sc_hd__inv_2 _05875_ (.A(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__nand2_1 _05876_ (.A(_05002_),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__nand2_1 _05877_ (.A(_05001_),
    .B(_05003_),
    .Y(_05006_));
 sky130_fd_sc_hd__nand3b_1 _05878_ (.A_N(_05000_),
    .B(_05005_),
    .C(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_1 _05879_ (.A(_05007_),
    .B(_05005_),
    .Y(_05008_));
 sky130_fd_sc_hd__nor2_1 _05880_ (.A(_04998_),
    .B(_04991_),
    .Y(_05009_));
 sky130_fd_sc_hd__a21oi_1 _05881_ (.A1(_04999_),
    .A2(_05008_),
    .B1(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__nand2_1 _05882_ (.A(_04988_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__nor2_1 _05883_ (.A(_05010_),
    .B(_04988_),
    .Y(_05012_));
 sky130_fd_sc_hd__a21oi_1 _05884_ (.A1(_04981_),
    .A2(_05011_),
    .B1(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__inv_2 _05885_ (.A(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__nand2_1 _05886_ (.A(_04973_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__nand3_1 _05887_ (.A(_04971_),
    .B(_04972_),
    .C(_05013_),
    .Y(_05016_));
 sky130_fd_sc_hd__nand2_1 _05888_ (.A(_05015_),
    .B(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__inv_2 _05889_ (.A(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__nor2_1 _05890_ (.A(_04796_),
    .B(_03534_),
    .Y(_05019_));
 sky130_fd_sc_hd__a21o_1 _05891_ (.A1(_04805_),
    .A2(_05018_),
    .B1(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__nor2_1 _05892_ (.A(_02467_),
    .B(_02456_),
    .Y(_05021_));
 sky130_fd_sc_hd__a21oi_2 _05893_ (.A1(_02478_),
    .A2(_03479_),
    .B1(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__nor2_1 _05894_ (.A(_02093_),
    .B(_02049_),
    .Y(_05023_));
 sky130_fd_sc_hd__a21oi_2 _05895_ (.A1(_02390_),
    .A2(_02379_),
    .B1(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__inv_2 _05896_ (.A(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__nand2_1 _05897_ (.A(_01796_),
    .B(_01818_),
    .Y(_05026_));
 sky130_fd_sc_hd__nor2_1 _05898_ (.A(_01818_),
    .B(_01796_),
    .Y(_05027_));
 sky130_fd_sc_hd__a21oi_2 _05899_ (.A1(_05026_),
    .A2(_02016_),
    .B1(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__inv_2 _05900_ (.A(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__nand2_1 _05901_ (.A(net55),
    .B(_00685_),
    .Y(_05030_));
 sky130_fd_sc_hd__inv_2 _05902_ (.A(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_1 _05903_ (.A(_00300_),
    .B(_00421_),
    .Y(_05032_));
 sky130_fd_sc_hd__inv_2 _05904_ (.A(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__nand2_1 _05905_ (.A(_05031_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_1 _05906_ (.A(_05030_),
    .B(_05032_),
    .Y(_05035_));
 sky130_fd_sc_hd__nand2_1 _05907_ (.A(_05034_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_1 _05908_ (.A(_00410_),
    .B(_01895_),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _05909_ (.A(_05036_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__inv_2 _05910_ (.A(_05037_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand3_1 _05911_ (.A(_05034_),
    .B(_05039_),
    .C(_05035_),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_1 _05912_ (.A(_05038_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__nor2_1 _05913_ (.A(_01686_),
    .B(_01664_),
    .Y(_05042_));
 sky130_fd_sc_hd__a21oi_2 _05914_ (.A1(_01774_),
    .A2(_01763_),
    .B1(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__inv_2 _05915_ (.A(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__nand2_1 _05916_ (.A(_05041_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand3_1 _05917_ (.A(_05038_),
    .B(_05043_),
    .C(_05040_),
    .Y(_05046_));
 sky130_fd_sc_hd__nand2_1 _05918_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_1 _05919_ (.A(_00641_),
    .B(_00355_),
    .Y(_05048_));
 sky130_fd_sc_hd__buf_4 _05920_ (.A(net15),
    .X(_05049_));
 sky130_fd_sc_hd__nand2_1 _05921_ (.A(_00674_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__nor2_1 _05922_ (.A(_05048_),
    .B(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__inv_2 _05923_ (.A(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__nand2_1 _05924_ (.A(_05048_),
    .B(_05050_),
    .Y(_05053_));
 sky130_fd_sc_hd__nand2_1 _05925_ (.A(_05052_),
    .B(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__nand2_1 _05926_ (.A(_00751_),
    .B(_00311_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_1 _05927_ (.A(_05054_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__inv_2 _05928_ (.A(_05055_),
    .Y(_05057_));
 sky130_fd_sc_hd__nand3_1 _05929_ (.A(_05052_),
    .B(_05053_),
    .C(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand2_1 _05930_ (.A(_05056_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__inv_2 _05931_ (.A(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_1 _05932_ (.A(_05047_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__nand3_1 _05933_ (.A(_05045_),
    .B(_05046_),
    .C(_05059_),
    .Y(_05062_));
 sky130_fd_sc_hd__nand2_1 _05934_ (.A(_05061_),
    .B(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _05935_ (.A(_05029_),
    .B(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand3_1 _05936_ (.A(_05028_),
    .B(_05061_),
    .C(_05062_),
    .Y(_05065_));
 sky130_fd_sc_hd__nand2_1 _05937_ (.A(_05064_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__nand2_1 _05938_ (.A(_01224_),
    .B(_00960_),
    .Y(_05067_));
 sky130_fd_sc_hd__clkbuf_8 _05939_ (.A(_01257_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _05940_ (.A(_05068_),
    .B(_00520_),
    .Y(_05069_));
 sky130_fd_sc_hd__or2_1 _05941_ (.A(_05067_),
    .B(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__nand2_1 _05942_ (.A(_05067_),
    .B(_05069_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _05943_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_1 _05944_ (.A(_02203_),
    .B(_04128_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_1 _05945_ (.A(_05072_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand3b_1 _05946_ (.A_N(_05073_),
    .B(_05070_),
    .C(_05071_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand2_1 _05947_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__nor2_1 _05948_ (.A(_01873_),
    .B(_01906_),
    .Y(_05077_));
 sky130_fd_sc_hd__a21oi_2 _05949_ (.A1(_01939_),
    .A2(_01983_),
    .B1(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__inv_2 _05950_ (.A(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2_1 _05951_ (.A(_05076_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand3_1 _05952_ (.A(_05074_),
    .B(_05075_),
    .C(_05078_),
    .Y(_05081_));
 sky130_fd_sc_hd__nand2_1 _05953_ (.A(_05080_),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__nand2_1 _05954_ (.A(_02247_),
    .B(_02170_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _05955_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__inv_2 _05956_ (.A(_05083_),
    .Y(_05085_));
 sky130_fd_sc_hd__nand3_1 _05957_ (.A(_05080_),
    .B(_05081_),
    .C(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__nand2_1 _05958_ (.A(_05084_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__inv_2 _05959_ (.A(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand2_1 _05960_ (.A(_05066_),
    .B(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__nand3_1 _05961_ (.A(_05064_),
    .B(_05065_),
    .C(_05087_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2_1 _05962_ (.A(_05089_),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__nand2_1 _05963_ (.A(_05025_),
    .B(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__nand3_1 _05964_ (.A(_05024_),
    .B(_05089_),
    .C(_05090_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _05965_ (.A(_05092_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__nand2_1 _05966_ (.A(_03149_),
    .B(_03072_),
    .Y(_05095_));
 sky130_fd_sc_hd__clkbuf_8 _05967_ (.A(_02522_),
    .X(_05096_));
 sky130_fd_sc_hd__nand2_1 _05968_ (.A(_05096_),
    .B(_01334_),
    .Y(_05097_));
 sky130_fd_sc_hd__inv_2 _05969_ (.A(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__nand2_1 _05970_ (.A(_03039_),
    .B(_02214_),
    .Y(_05099_));
 sky130_fd_sc_hd__inv_2 _05971_ (.A(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _05972_ (.A(_05098_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__nand2_1 _05973_ (.A(_05097_),
    .B(_05099_),
    .Y(_05102_));
 sky130_fd_sc_hd__nand2_1 _05974_ (.A(_05101_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__nand2_1 _05975_ (.A(_01532_),
    .B(_02687_),
    .Y(_05104_));
 sky130_fd_sc_hd__nand2_1 _05976_ (.A(_05103_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__inv_2 _05977_ (.A(_05104_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand3_1 _05978_ (.A(_05101_),
    .B(_05106_),
    .C(_05102_),
    .Y(_05107_));
 sky130_fd_sc_hd__nand3_1 _05979_ (.A(_05095_),
    .B(_05105_),
    .C(_05107_),
    .Y(_05108_));
 sky130_fd_sc_hd__nand2_1 _05980_ (.A(_05105_),
    .B(_05107_),
    .Y(_05109_));
 sky130_fd_sc_hd__a21boi_1 _05981_ (.A1(_03138_),
    .A2(_03083_),
    .B1_N(_03072_),
    .Y(_05110_));
 sky130_fd_sc_hd__nand2_1 _05982_ (.A(_05109_),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__nand2_1 _05983_ (.A(_05108_),
    .B(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__clkbuf_8 _05984_ (.A(_02511_),
    .X(_05113_));
 sky130_fd_sc_hd__clkbuf_8 _05985_ (.A(net37),
    .X(_05114_));
 sky130_fd_sc_hd__nand2_1 _05986_ (.A(_05113_),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand2_1 _05987_ (.A(_03105_),
    .B(_03248_),
    .Y(_05116_));
 sky130_fd_sc_hd__nor2_1 _05988_ (.A(_05115_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__inv_2 _05989_ (.A(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__nand2_1 _05990_ (.A(_05115_),
    .B(_05116_),
    .Y(_05119_));
 sky130_fd_sc_hd__nand2_1 _05991_ (.A(_05118_),
    .B(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2_1 _05992_ (.A(_02555_),
    .B(_04645_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand2_1 _05993_ (.A(_05120_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__inv_2 _05994_ (.A(_05121_),
    .Y(_05123_));
 sky130_fd_sc_hd__nand3_1 _05995_ (.A(_05118_),
    .B(_05123_),
    .C(_05119_),
    .Y(_05124_));
 sky130_fd_sc_hd__nand2_1 _05996_ (.A(_05122_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__nand2_1 _05997_ (.A(_05112_),
    .B(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand3b_1 _05998_ (.A_N(_05125_),
    .B(_05108_),
    .C(_05111_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _05999_ (.A(_05126_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__nand2_1 _06000_ (.A(_02258_),
    .B(_02280_),
    .Y(_05129_));
 sky130_fd_sc_hd__nor2_1 _06001_ (.A(_02280_),
    .B(_02258_),
    .Y(_05130_));
 sky130_fd_sc_hd__a21oi_2 _06002_ (.A1(_05129_),
    .A2(_02335_),
    .B1(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__inv_2 _06003_ (.A(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand2_1 _06004_ (.A(_05128_),
    .B(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand3_1 _06005_ (.A(_05131_),
    .B(_05126_),
    .C(_05127_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_1 _06006_ (.A(_05133_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21ai_2 _06007_ (.A1(_03182_),
    .A2(_03160_),
    .B1(_03380_),
    .Y(_05136_));
 sky130_fd_sc_hd__nand2_1 _06008_ (.A(_05135_),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand3b_1 _06009_ (.A_N(_05136_),
    .B(_05133_),
    .C(_05134_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_1 _06010_ (.A(_05137_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__inv_2 _06011_ (.A(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__nand2_1 _06012_ (.A(_05094_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand3_1 _06013_ (.A(_05092_),
    .B(_05093_),
    .C(_05139_),
    .Y(_05142_));
 sky130_fd_sc_hd__nand3_1 _06014_ (.A(_05022_),
    .B(_05141_),
    .C(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__nand2_1 _06015_ (.A(_05141_),
    .B(_05142_),
    .Y(_05144_));
 sky130_fd_sc_hd__nand2_1 _06016_ (.A(_03490_),
    .B(_02445_),
    .Y(_05145_));
 sky130_fd_sc_hd__nand2_1 _06017_ (.A(_05144_),
    .B(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_1 _06018_ (.A(_05143_),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__o21ai_1 _06019_ (.A1(_04906_),
    .A2(_04930_),
    .B1(_04964_),
    .Y(_05148_));
 sky130_fd_sc_hd__nor2_1 _06020_ (.A(_04907_),
    .B(_04920_),
    .Y(_05149_));
 sky130_fd_sc_hd__a21oi_2 _06021_ (.A1(_04921_),
    .A2(_04922_),
    .B1(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__inv_2 _06022_ (.A(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__nand2_1 _06023_ (.A(_02874_),
    .B(_04899_),
    .Y(_05152_));
 sky130_fd_sc_hd__inv_2 _06024_ (.A(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__nand2_1 _06025_ (.A(_02797_),
    .B(_04897_),
    .Y(_05154_));
 sky130_fd_sc_hd__inv_2 _06026_ (.A(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_1 _06027_ (.A(_05153_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__nand2_1 _06028_ (.A(_05152_),
    .B(_05154_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2_1 _06029_ (.A(_05156_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__buf_8 _06030_ (.A(_04634_),
    .X(_05159_));
 sky130_fd_sc_hd__nand2_1 _06031_ (.A(_05159_),
    .B(_04888_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_1 _06032_ (.A(_05158_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__nand3b_1 _06033_ (.A_N(_05160_),
    .B(_05156_),
    .C(_05157_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_1 _06034_ (.A(_05161_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__a21oi_2 _06035_ (.A1(_03292_),
    .A2(_03336_),
    .B1(_03270_),
    .Y(_05164_));
 sky130_fd_sc_hd__inv_2 _06036_ (.A(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_1 _06037_ (.A(_05163_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand3_1 _06038_ (.A(_05161_),
    .B(_05162_),
    .C(_05164_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand2_1 _06039_ (.A(_05166_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand2_1 _06040_ (.A(_04916_),
    .B(_04914_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_1 _06041_ (.A(_05168_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__nand3b_1 _06042_ (.A_N(_05169_),
    .B(_05166_),
    .C(_05167_),
    .Y(_05171_));
 sky130_fd_sc_hd__nand2_1 _06043_ (.A(_05170_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__nand2_1 _06044_ (.A(_05151_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__nand3_1 _06045_ (.A(_05150_),
    .B(_05170_),
    .C(_05171_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_1 _06046_ (.A(_05173_),
    .B(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__nand2_1 _06047_ (.A(_04880_),
    .B(_04933_),
    .Y(_05176_));
 sky130_fd_sc_hd__nand3b_2 _06048_ (.A_N(_05176_),
    .B(_04814_),
    .C(_04936_),
    .Y(_05177_));
 sky130_fd_sc_hd__inv_2 _06049_ (.A(_04814_),
    .Y(_05178_));
 sky130_fd_sc_hd__inv_2 _06050_ (.A(_04936_),
    .Y(_05179_));
 sky130_fd_sc_hd__o21ai_1 _06051_ (.A1(_05178_),
    .A2(_05179_),
    .B1(_05176_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand2_1 _06052_ (.A(_05177_),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _06053_ (.A(_04895_),
    .B(_04941_),
    .Y(_05182_));
 sky130_fd_sc_hd__nand2_1 _06054_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__nand3b_2 _06055_ (.A_N(_05182_),
    .B(_05177_),
    .C(_05180_),
    .Y(_05184_));
 sky130_fd_sc_hd__nand2_1 _06056_ (.A(_05183_),
    .B(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__nand2_1 _06057_ (.A(_04945_),
    .B(_04939_),
    .Y(_05186_));
 sky130_fd_sc_hd__nand2_1 _06058_ (.A(_05185_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__inv_2 _06059_ (.A(_05186_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand3_1 _06060_ (.A(_05188_),
    .B(_05183_),
    .C(_05184_),
    .Y(_05189_));
 sky130_fd_sc_hd__nand2_1 _06061_ (.A(_05187_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__buf_4 _06062_ (.A(net47),
    .X(_05191_));
 sky130_fd_sc_hd__nand2_1 _06063_ (.A(_05191_),
    .B(net1),
    .Y(_05192_));
 sky130_fd_sc_hd__nand2_1 _06064_ (.A(net46),
    .B(_04947_),
    .Y(_05193_));
 sky130_fd_sc_hd__nor2_1 _06065_ (.A(_05192_),
    .B(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__inv_2 _06066_ (.A(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__nand2_1 _06067_ (.A(_05192_),
    .B(_05193_),
    .Y(_05196_));
 sky130_fd_sc_hd__nand2_1 _06068_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__inv_2 _06069_ (.A(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_1 _06070_ (.A(_05190_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__nand3_1 _06071_ (.A(_05187_),
    .B(_05189_),
    .C(_05197_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand2_1 _06072_ (.A(_05199_),
    .B(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__inv_2 _06073_ (.A(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__nand2_1 _06074_ (.A(_05175_),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__nand3_1 _06075_ (.A(_05173_),
    .B(_05174_),
    .C(_05201_),
    .Y(_05204_));
 sky130_fd_sc_hd__nand2_1 _06076_ (.A(_05203_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__nand2_1 _06077_ (.A(_03402_),
    .B(_02995_),
    .Y(_05206_));
 sky130_fd_sc_hd__nor2_1 _06078_ (.A(_02995_),
    .B(_03402_),
    .Y(_05207_));
 sky130_fd_sc_hd__a21oi_2 _06079_ (.A1(_05206_),
    .A2(_02962_),
    .B1(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__inv_2 _06080_ (.A(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__nand2_1 _06081_ (.A(_05205_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__nand3_1 _06082_ (.A(_05208_),
    .B(_05203_),
    .C(_05204_),
    .Y(_05211_));
 sky130_fd_sc_hd__nand3b_1 _06083_ (.A_N(_05148_),
    .B(_05210_),
    .C(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_1 _06084_ (.A(_05210_),
    .B(_05211_),
    .Y(_05213_));
 sky130_fd_sc_hd__nand2_1 _06085_ (.A(_05213_),
    .B(_05148_),
    .Y(_05214_));
 sky130_fd_sc_hd__nand2_1 _06086_ (.A(_05212_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__inv_2 _06087_ (.A(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_1 _06088_ (.A(_05147_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__nand3_1 _06089_ (.A(_05143_),
    .B(_05146_),
    .C(_05215_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand3_1 _06090_ (.A(_05020_),
    .B(_05217_),
    .C(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__and2_1 _06091_ (.A(_04961_),
    .B(_04956_),
    .X(_05220_));
 sky130_fd_sc_hd__o21a_1 _06092_ (.A1(_04966_),
    .A2(_04969_),
    .B1(_05015_),
    .X(_05221_));
 sky130_fd_sc_hd__nor2_1 _06093_ (.A(_05220_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__inv_2 _06094_ (.A(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__nand2_1 _06095_ (.A(_05221_),
    .B(_05220_),
    .Y(_05224_));
 sky130_fd_sc_hd__nand2_1 _06096_ (.A(_05223_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__inv_2 _06097_ (.A(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand2_1 _06098_ (.A(_05217_),
    .B(_05218_),
    .Y(_05227_));
 sky130_fd_sc_hd__a21oi_1 _06099_ (.A1(_04805_),
    .A2(_05018_),
    .B1(_05019_),
    .Y(_05228_));
 sky130_fd_sc_hd__nand2_1 _06100_ (.A(_05227_),
    .B(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__nand3_1 _06101_ (.A(_05219_),
    .B(_05226_),
    .C(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__nand2_1 _06102_ (.A(_05227_),
    .B(_05020_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand3_1 _06103_ (.A(_05228_),
    .B(_05217_),
    .C(_05218_),
    .Y(_05232_));
 sky130_fd_sc_hd__nand3_1 _06104_ (.A(_05231_),
    .B(_05232_),
    .C(_05225_),
    .Y(_05233_));
 sky130_fd_sc_hd__nand2_1 _06105_ (.A(_05230_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__nand3_1 _06106_ (.A(_04796_),
    .B(_03490_),
    .C(_03523_),
    .Y(_05235_));
 sky130_fd_sc_hd__a21o_1 _06107_ (.A1(_04315_),
    .A2(_04776_),
    .B1(_04785_),
    .X(_05236_));
 sky130_fd_sc_hd__nand2_1 _06108_ (.A(_03534_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__nand2_1 _06109_ (.A(_05235_),
    .B(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__nand2_1 _06110_ (.A(_05238_),
    .B(_05018_),
    .Y(_05239_));
 sky130_fd_sc_hd__nand3_1 _06111_ (.A(_05235_),
    .B(_05237_),
    .C(_05017_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2_1 _06112_ (.A(_05239_),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__nand3_1 _06113_ (.A(_05010_),
    .B(_04987_),
    .C(_04985_),
    .Y(_05242_));
 sky130_fd_sc_hd__a21o_1 _06114_ (.A1(_04999_),
    .A2(_05008_),
    .B1(_05009_),
    .X(_05243_));
 sky130_fd_sc_hd__nand2_1 _06115_ (.A(_05243_),
    .B(_04988_),
    .Y(_05244_));
 sky130_fd_sc_hd__nand2_1 _06116_ (.A(_05242_),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__nand2_1 _06117_ (.A(_05245_),
    .B(_04981_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand3_1 _06118_ (.A(_05242_),
    .B(_05244_),
    .C(_04980_),
    .Y(_05247_));
 sky130_fd_sc_hd__nand2_1 _06119_ (.A(_05246_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__nand2_1 _06120_ (.A(_04458_),
    .B(_04557_),
    .Y(_05249_));
 sky130_fd_sc_hd__nand3_1 _06121_ (.A(_04436_),
    .B(_04447_),
    .C(_04535_),
    .Y(_05250_));
 sky130_fd_sc_hd__nand3_1 _06122_ (.A(_05249_),
    .B(_05250_),
    .C(_04700_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_1 _06123_ (.A(_04722_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_1 _06124_ (.A(_03864_),
    .B(_03875_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2_1 _06125_ (.A(_05253_),
    .B(_03809_),
    .Y(_05254_));
 sky130_fd_sc_hd__nand2_1 _06126_ (.A(_05254_),
    .B(_03886_),
    .Y(_05255_));
 sky130_fd_sc_hd__nand2_1 _06127_ (.A(_00641_),
    .B(net5),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_1 _06128_ (.A(_00674_),
    .B(_00311_),
    .Y(_05257_));
 sky130_fd_sc_hd__nand2_1 _06129_ (.A(_05256_),
    .B(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__nand2_1 _06130_ (.A(_00751_),
    .B(net4),
    .Y(_05259_));
 sky130_fd_sc_hd__inv_2 _06131_ (.A(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__nor2_1 _06132_ (.A(_05256_),
    .B(_05257_),
    .Y(_05261_));
 sky130_fd_sc_hd__a21oi_2 _06133_ (.A1(_05258_),
    .A2(_05260_),
    .B1(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__nand2_1 _06134_ (.A(_05255_),
    .B(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__nand2_1 _06135_ (.A(_02489_),
    .B(_01224_),
    .Y(_05264_));
 sky130_fd_sc_hd__inv_2 _06136_ (.A(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_1 _06137_ (.A(_01521_),
    .B(_01257_),
    .Y(_05266_));
 sky130_fd_sc_hd__inv_2 _06138_ (.A(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand2_1 _06139_ (.A(_05265_),
    .B(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _06140_ (.A(_02511_),
    .B(_01323_),
    .Y(_05269_));
 sky130_fd_sc_hd__inv_2 _06141_ (.A(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_1 _06142_ (.A(_05264_),
    .B(_05266_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand3_1 _06143_ (.A(_05268_),
    .B(_05270_),
    .C(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand2_1 _06144_ (.A(_05272_),
    .B(_05268_),
    .Y(_05273_));
 sky130_fd_sc_hd__nor2_1 _06145_ (.A(_05262_),
    .B(_05255_),
    .Y(_05274_));
 sky130_fd_sc_hd__a21oi_2 _06146_ (.A1(_05263_),
    .A2(_05273_),
    .B1(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_1 _06147_ (.A(_05252_),
    .B(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_2 _06148_ (.A(_02797_),
    .B(_02522_),
    .Y(_05277_));
 sky130_fd_sc_hd__clkbuf_8 _06149_ (.A(_02555_),
    .X(_05278_));
 sky130_fd_sc_hd__nand2_2 _06150_ (.A(_05278_),
    .B(net64),
    .Y(_05279_));
 sky130_fd_sc_hd__nand2_1 _06151_ (.A(_05277_),
    .B(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__nand2_1 _06152_ (.A(_02874_),
    .B(net35),
    .Y(_05281_));
 sky130_fd_sc_hd__inv_2 _06153_ (.A(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__nor2_1 _06154_ (.A(_05277_),
    .B(_05279_),
    .Y(_05283_));
 sky130_fd_sc_hd__a21oi_2 _06155_ (.A1(_05280_),
    .A2(_05282_),
    .B1(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__inv_2 _06156_ (.A(_04480_),
    .Y(_05285_));
 sky130_fd_sc_hd__nand2_1 _06157_ (.A(_05285_),
    .B(_04469_),
    .Y(_05286_));
 sky130_fd_sc_hd__inv_2 _06158_ (.A(_04469_),
    .Y(_05287_));
 sky130_fd_sc_hd__nand2_1 _06159_ (.A(_05287_),
    .B(_04480_),
    .Y(_05288_));
 sky130_fd_sc_hd__nand3_1 _06160_ (.A(_05286_),
    .B(_05288_),
    .C(_04502_),
    .Y(_05289_));
 sky130_fd_sc_hd__nand2_1 _06161_ (.A(_05287_),
    .B(_05285_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand3_1 _06162_ (.A(_05290_),
    .B(_04513_),
    .C(_04491_),
    .Y(_05291_));
 sky130_fd_sc_hd__nand2_1 _06163_ (.A(_05289_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__inv_2 _06164_ (.A(_05284_),
    .Y(_05293_));
 sky130_fd_sc_hd__nand2_1 _06165_ (.A(_05292_),
    .B(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__nand3_1 _06166_ (.A(_05284_),
    .B(_05289_),
    .C(_05291_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_1 _06167_ (.A(_05294_),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__inv_2 _06168_ (.A(_04994_),
    .Y(_05297_));
 sky130_fd_sc_hd__o21ai_1 _06169_ (.A1(_04997_),
    .A2(_05297_),
    .B1(_04995_),
    .Y(_05298_));
 sky130_fd_sc_hd__nand3b_1 _06170_ (.A_N(_04997_),
    .B(_04996_),
    .C(_04994_),
    .Y(_05299_));
 sky130_fd_sc_hd__nand2_1 _06171_ (.A(_05298_),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__inv_2 _06172_ (.A(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__nand2_1 _06173_ (.A(_05296_),
    .B(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__o21ai_2 _06174_ (.A1(_05284_),
    .A2(_05292_),
    .B1(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__nor2_1 _06175_ (.A(_05275_),
    .B(_05252_),
    .Y(_05304_));
 sky130_fd_sc_hd__a21oi_2 _06176_ (.A1(_05276_),
    .A2(_05303_),
    .B1(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__inv_2 _06177_ (.A(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand2_1 _06178_ (.A(_05248_),
    .B(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__nand3_1 _06179_ (.A(_05305_),
    .B(_05246_),
    .C(_05247_),
    .Y(_05308_));
 sky130_fd_sc_hd__nand2_1 _06180_ (.A(_05307_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__buf_6 _06181_ (.A(_04947_),
    .X(_05310_));
 sky130_fd_sc_hd__a22o_1 _06182_ (.A1(_05310_),
    .A2(_04936_),
    .B1(_04958_),
    .B2(_04933_),
    .X(_05311_));
 sky130_fd_sc_hd__nand2_1 _06183_ (.A(_04975_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__inv_2 _06184_ (.A(_04998_),
    .Y(_05313_));
 sky130_fd_sc_hd__nand2_1 _06185_ (.A(_04991_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__nand3_1 _06186_ (.A(_04990_),
    .B(_04903_),
    .C(_04998_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_1 _06187_ (.A(_05314_),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_1 _06188_ (.A(_05316_),
    .B(_05008_),
    .Y(_05317_));
 sky130_fd_sc_hd__nand3b_1 _06189_ (.A_N(_05008_),
    .B(_05314_),
    .C(_05315_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand2_1 _06190_ (.A(_05317_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand2_1 _06191_ (.A(_04814_),
    .B(net37),
    .Y(_05320_));
 sky130_fd_sc_hd__nand2_1 _06192_ (.A(_04634_),
    .B(_03248_),
    .Y(_05321_));
 sky130_fd_sc_hd__nand2_1 _06193_ (.A(_05320_),
    .B(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand2_1 _06194_ (.A(_04880_),
    .B(net38),
    .Y(_05323_));
 sky130_fd_sc_hd__inv_2 _06195_ (.A(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__nor2_1 _06196_ (.A(_05320_),
    .B(_05321_),
    .Y(_05325_));
 sky130_fd_sc_hd__a21oi_1 _06197_ (.A1(_05322_),
    .A2(_05324_),
    .B1(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__inv_2 _06198_ (.A(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__nand2_1 _06199_ (.A(_05005_),
    .B(_05006_),
    .Y(_05328_));
 sky130_fd_sc_hd__nand2_1 _06200_ (.A(_05328_),
    .B(_05000_),
    .Y(_05329_));
 sky130_fd_sc_hd__nand3_1 _06201_ (.A(_05327_),
    .B(_05007_),
    .C(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _06202_ (.A(_05329_),
    .B(_05007_),
    .Y(_05331_));
 sky130_fd_sc_hd__nand2_1 _06203_ (.A(_05331_),
    .B(_05326_),
    .Y(_05332_));
 sky130_fd_sc_hd__nand2_1 _06204_ (.A(net1),
    .B(_04888_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand2_1 _06205_ (.A(_04947_),
    .B(_04899_),
    .Y(_05334_));
 sky130_fd_sc_hd__inv_2 _06206_ (.A(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand2_1 _06207_ (.A(_04895_),
    .B(_04897_),
    .Y(_05336_));
 sky130_fd_sc_hd__inv_2 _06208_ (.A(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__nand2_1 _06209_ (.A(_05335_),
    .B(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _06210_ (.A(_05334_),
    .B(_05336_),
    .Y(_00000_));
 sky130_fd_sc_hd__nand3b_1 _06211_ (.A_N(_05333_),
    .B(_05338_),
    .C(_00000_),
    .Y(_00001_));
 sky130_fd_sc_hd__nand2_1 _06212_ (.A(_00001_),
    .B(_05338_),
    .Y(_00002_));
 sky130_fd_sc_hd__nand3_1 _06213_ (.A(_05330_),
    .B(_05332_),
    .C(_00002_),
    .Y(_00003_));
 sky130_fd_sc_hd__nand2_1 _06214_ (.A(_00003_),
    .B(_05330_),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _06215_ (.A(_00004_),
    .Y(_00005_));
 sky130_fd_sc_hd__nand2_1 _06216_ (.A(_05319_),
    .B(_00005_),
    .Y(_00006_));
 sky130_fd_sc_hd__nand3_1 _06217_ (.A(_00004_),
    .B(_05317_),
    .C(_05318_),
    .Y(_00007_));
 sky130_fd_sc_hd__nand3b_1 _06218_ (.A_N(_05312_),
    .B(_00006_),
    .C(_00007_),
    .Y(_00008_));
 sky130_fd_sc_hd__nand2_1 _06219_ (.A(_00008_),
    .B(_00007_),
    .Y(_00009_));
 sky130_fd_sc_hd__nand2_1 _06220_ (.A(_05309_),
    .B(_00009_),
    .Y(_00010_));
 sky130_fd_sc_hd__nand3b_1 _06221_ (.A_N(_00009_),
    .B(_05307_),
    .C(_05308_),
    .Y(_00011_));
 sky130_fd_sc_hd__nand2_1 _06222_ (.A(_00010_),
    .B(_00011_),
    .Y(_00012_));
 sky130_fd_sc_hd__inv_2 _06223_ (.A(_00012_),
    .Y(_00013_));
 sky130_fd_sc_hd__inv_2 _06224_ (.A(_03611_),
    .Y(_00014_));
 sky130_fd_sc_hd__inv_2 _06225_ (.A(_04304_),
    .Y(_00015_));
 sky130_fd_sc_hd__nand2_1 _06226_ (.A(_00014_),
    .B(_00015_),
    .Y(_00016_));
 sky130_fd_sc_hd__nand3_1 _06227_ (.A(_00016_),
    .B(_04776_),
    .C(_04315_),
    .Y(_00017_));
 sky130_fd_sc_hd__nand2_1 _06228_ (.A(_00014_),
    .B(_04304_),
    .Y(_00018_));
 sky130_fd_sc_hd__nand2_1 _06229_ (.A(_00015_),
    .B(_03611_),
    .Y(_00019_));
 sky130_fd_sc_hd__nand3_1 _06230_ (.A(_00018_),
    .B(_04766_),
    .C(_00019_),
    .Y(_00020_));
 sky130_fd_sc_hd__nand2_1 _06231_ (.A(_00017_),
    .B(_00020_),
    .Y(_00021_));
 sky130_fd_sc_hd__inv_2 _06232_ (.A(_05275_),
    .Y(_00022_));
 sky130_fd_sc_hd__nand2_1 _06233_ (.A(_05252_),
    .B(_00022_),
    .Y(_00023_));
 sky130_fd_sc_hd__nand3_1 _06234_ (.A(_05275_),
    .B(_04722_),
    .C(_05251_),
    .Y(_00024_));
 sky130_fd_sc_hd__nand2_1 _06235_ (.A(_00023_),
    .B(_00024_),
    .Y(_00025_));
 sky130_fd_sc_hd__nand2_1 _06236_ (.A(_00025_),
    .B(_05303_),
    .Y(_00026_));
 sky130_fd_sc_hd__nand3b_1 _06237_ (.A_N(_05303_),
    .B(_00023_),
    .C(_00024_),
    .Y(_00027_));
 sky130_fd_sc_hd__nand2_1 _06238_ (.A(_00026_),
    .B(_00027_),
    .Y(_00028_));
 sky130_fd_sc_hd__inv_2 _06239_ (.A(_00028_),
    .Y(_00029_));
 sky130_fd_sc_hd__nand3_1 _06240_ (.A(_04271_),
    .B(_03996_),
    .C(_04007_),
    .Y(_00030_));
 sky130_fd_sc_hd__inv_2 _06241_ (.A(_04194_),
    .Y(_00031_));
 sky130_fd_sc_hd__nand3_1 _06242_ (.A(_00031_),
    .B(_04095_),
    .C(_04073_),
    .Y(_00032_));
 sky130_fd_sc_hd__nand3_2 _06243_ (.A(_00032_),
    .B(_04205_),
    .C(_04249_),
    .Y(_00033_));
 sky130_fd_sc_hd__nand2_1 _06244_ (.A(_00033_),
    .B(_00032_),
    .Y(_00034_));
 sky130_fd_sc_hd__nand2_1 _06245_ (.A(_04018_),
    .B(_00034_),
    .Y(_00035_));
 sky130_fd_sc_hd__nand2_1 _06246_ (.A(_00030_),
    .B(_00035_),
    .Y(_00036_));
 sky130_fd_sc_hd__nand2_1 _06247_ (.A(_00036_),
    .B(_03941_),
    .Y(_00037_));
 sky130_fd_sc_hd__nand3_1 _06248_ (.A(_00030_),
    .B(_00035_),
    .C(_03930_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _06249_ (.A(_00037_),
    .B(_00038_),
    .Y(_00039_));
 sky130_fd_sc_hd__inv_2 _06250_ (.A(_05262_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand3_1 _06251_ (.A(_00040_),
    .B(_03886_),
    .C(_05254_),
    .Y(_00041_));
 sky130_fd_sc_hd__nand2_1 _06252_ (.A(_00041_),
    .B(_05263_),
    .Y(_00042_));
 sky130_fd_sc_hd__and2_1 _06253_ (.A(_05272_),
    .B(_05268_),
    .X(_00043_));
 sky130_fd_sc_hd__nand2_1 _06254_ (.A(_00042_),
    .B(_00043_),
    .Y(_00044_));
 sky130_fd_sc_hd__nand3_1 _06255_ (.A(_00041_),
    .B(_05263_),
    .C(_05273_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand2_1 _06256_ (.A(_00044_),
    .B(_00045_),
    .Y(_00046_));
 sky130_fd_sc_hd__inv_2 _06257_ (.A(_00046_),
    .Y(_00047_));
 sky130_fd_sc_hd__nand2_1 _06258_ (.A(_04106_),
    .B(_00031_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand3_1 _06259_ (.A(_04194_),
    .B(_04073_),
    .C(_04095_),
    .Y(_00049_));
 sky130_fd_sc_hd__nand3_1 _06260_ (.A(_00048_),
    .B(_00049_),
    .C(_04238_),
    .Y(_00050_));
 sky130_fd_sc_hd__nand2_1 _06261_ (.A(_00033_),
    .B(_00050_),
    .Y(_00051_));
 sky130_fd_sc_hd__inv_2 _06262_ (.A(_04139_),
    .Y(_00052_));
 sky130_fd_sc_hd__nand2_1 _06263_ (.A(_00052_),
    .B(_04117_),
    .Y(_00053_));
 sky130_fd_sc_hd__inv_2 _06264_ (.A(_04117_),
    .Y(_00054_));
 sky130_fd_sc_hd__nand2_1 _06265_ (.A(_00054_),
    .B(_04139_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand3_1 _06266_ (.A(_00053_),
    .B(_00055_),
    .C(_04161_),
    .Y(_00056_));
 sky130_fd_sc_hd__nand2_1 _06267_ (.A(_00054_),
    .B(_00052_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand3_1 _06268_ (.A(_00057_),
    .B(_04172_),
    .C(_04150_),
    .Y(_00058_));
 sky130_fd_sc_hd__nand2_1 _06269_ (.A(_00056_),
    .B(_00058_),
    .Y(_00059_));
 sky130_fd_sc_hd__nand2_1 _06270_ (.A(_00344_),
    .B(_04128_),
    .Y(_00060_));
 sky130_fd_sc_hd__nand2_1 _06271_ (.A(_00300_),
    .B(_02214_),
    .Y(_00061_));
 sky130_fd_sc_hd__nand2_1 _06272_ (.A(_00060_),
    .B(_00061_),
    .Y(_00062_));
 sky130_fd_sc_hd__nand2_1 _06273_ (.A(_00410_),
    .B(_00960_),
    .Y(_00063_));
 sky130_fd_sc_hd__inv_2 _06274_ (.A(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__nor2_1 _06275_ (.A(_00060_),
    .B(_00061_),
    .Y(_00065_));
 sky130_fd_sc_hd__a21oi_2 _06276_ (.A1(_00062_),
    .A2(_00064_),
    .B1(_00065_),
    .Y(_00066_));
 sky130_fd_sc_hd__nand2_1 _06277_ (.A(_00059_),
    .B(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _06278_ (.A(_05257_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_1 _06279_ (.A(_00068_),
    .B(_05256_),
    .Y(_00069_));
 sky130_fd_sc_hd__inv_2 _06280_ (.A(_05256_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_1 _06281_ (.A(_00070_),
    .B(_05257_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand3_1 _06282_ (.A(_00069_),
    .B(_00071_),
    .C(_05259_),
    .Y(_00072_));
 sky130_fd_sc_hd__nand2_1 _06283_ (.A(_00070_),
    .B(_00068_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand3_1 _06284_ (.A(_00073_),
    .B(_05260_),
    .C(_05258_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_1 _06285_ (.A(_00072_),
    .B(_00074_),
    .Y(_00075_));
 sky130_fd_sc_hd__inv_2 _06286_ (.A(_00075_),
    .Y(_00076_));
 sky130_fd_sc_hd__nor2_1 _06287_ (.A(_00066_),
    .B(_00059_),
    .Y(_00077_));
 sky130_fd_sc_hd__a21oi_1 _06288_ (.A1(_00067_),
    .A2(_00076_),
    .B1(_00077_),
    .Y(_00078_));
 sky130_fd_sc_hd__nand2_1 _06289_ (.A(_00051_),
    .B(_00078_),
    .Y(_00079_));
 sky130_fd_sc_hd__nor2_1 _06290_ (.A(_00078_),
    .B(_00051_),
    .Y(_00080_));
 sky130_fd_sc_hd__a21oi_1 _06291_ (.A1(_00047_),
    .A2(_00079_),
    .B1(_00080_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _06292_ (.A(_00039_),
    .B(_00081_),
    .Y(_00082_));
 sky130_fd_sc_hd__nor2_1 _06293_ (.A(_00081_),
    .B(_00039_),
    .Y(_00083_));
 sky130_fd_sc_hd__a21oi_2 _06294_ (.A1(_00029_),
    .A2(_00082_),
    .B1(_00083_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _06295_ (.A(_00021_),
    .B(_00084_),
    .Y(_00085_));
 sky130_fd_sc_hd__nor2_1 _06296_ (.A(_00084_),
    .B(_00021_),
    .Y(_00086_));
 sky130_fd_sc_hd__a21oi_2 _06297_ (.A1(_00013_),
    .A2(_00085_),
    .B1(_00086_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand2_1 _06298_ (.A(_05241_),
    .B(_00087_),
    .Y(_00088_));
 sky130_fd_sc_hd__or2_1 _06299_ (.A(_05305_),
    .B(_05248_),
    .X(_00089_));
 sky130_fd_sc_hd__and2_1 _06300_ (.A(_00010_),
    .B(_00089_),
    .X(_00090_));
 sky130_fd_sc_hd__nor2_1 _06301_ (.A(_04978_),
    .B(_00090_),
    .Y(_00091_));
 sky130_fd_sc_hd__nand2_1 _06302_ (.A(_00090_),
    .B(_04978_),
    .Y(_00092_));
 sky130_fd_sc_hd__nor2b_1 _06303_ (.A(_00091_),
    .B_N(_00092_),
    .Y(_00093_));
 sky130_fd_sc_hd__nor2_1 _06304_ (.A(_00087_),
    .B(_05241_),
    .Y(_00094_));
 sky130_fd_sc_hd__a21o_1 _06305_ (.A1(_00088_),
    .A2(_00093_),
    .B1(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__nand2_1 _06306_ (.A(_05234_),
    .B(_00095_),
    .Y(_00096_));
 sky130_fd_sc_hd__a21oi_1 _06307_ (.A1(_00088_),
    .A2(_00093_),
    .B1(_00094_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand3_1 _06308_ (.A(_00097_),
    .B(_05230_),
    .C(_05233_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_1 _06309_ (.A(_00096_),
    .B(_00098_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand2_1 _06310_ (.A(_00099_),
    .B(_00091_),
    .Y(_00100_));
 sky130_fd_sc_hd__nand3b_2 _06311_ (.A_N(_00091_),
    .B(_00096_),
    .C(_00098_),
    .Y(_00101_));
 sky130_fd_sc_hd__nand2_1 _06312_ (.A(_00100_),
    .B(_00101_),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_2 _06313_ (.A(_00084_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_1 _06314_ (.A(_00021_),
    .B(_00103_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand3_1 _06315_ (.A(_00084_),
    .B(_00017_),
    .C(_00020_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_1 _06316_ (.A(_00104_),
    .B(_00105_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_1 _06317_ (.A(_00106_),
    .B(_00013_),
    .Y(_00107_));
 sky130_fd_sc_hd__nand3_1 _06318_ (.A(_00104_),
    .B(_00105_),
    .C(_00012_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_1 _06319_ (.A(_00107_),
    .B(_00108_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand3_1 _06320_ (.A(_05294_),
    .B(_05295_),
    .C(_05300_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_1 _06321_ (.A(_05302_),
    .B(_00110_),
    .Y(_00111_));
 sky130_fd_sc_hd__nand2_1 _06322_ (.A(_05267_),
    .B(_05264_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _06323_ (.A(_05265_),
    .B(_05266_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand3_1 _06324_ (.A(_00112_),
    .B(_00113_),
    .C(_05269_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _06325_ (.A(_00114_),
    .B(_05272_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_1 _06326_ (.A(_00641_),
    .B(_01334_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_1 _06327_ (.A(_00674_),
    .B(_00520_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_1 _06328_ (.A(_00116_),
    .B(_00117_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_1 _06329_ (.A(_01521_),
    .B(_00751_),
    .Y(_00119_));
 sky130_fd_sc_hd__inv_2 _06330_ (.A(_00119_),
    .Y(_00120_));
 sky130_fd_sc_hd__nor2_1 _06331_ (.A(_00116_),
    .B(_00117_),
    .Y(_00121_));
 sky130_fd_sc_hd__a21oi_2 _06332_ (.A1(_00118_),
    .A2(_00120_),
    .B1(_00121_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_1 _06333_ (.A(_00115_),
    .B(_00122_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _06334_ (.A(_02489_),
    .B(_01257_),
    .Y(_00124_));
 sky130_fd_sc_hd__inv_2 _06335_ (.A(_00124_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _06336_ (.A(_02511_),
    .B(_01224_),
    .Y(_00126_));
 sky130_fd_sc_hd__inv_2 _06337_ (.A(_00126_),
    .Y(_00127_));
 sky130_fd_sc_hd__nand2_1 _06338_ (.A(_00125_),
    .B(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _06339_ (.A(_05278_),
    .B(_01323_),
    .Y(_00129_));
 sky130_fd_sc_hd__inv_2 _06340_ (.A(_00129_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _06341_ (.A(_00124_),
    .B(_00126_),
    .Y(_00131_));
 sky130_fd_sc_hd__nand3_1 _06342_ (.A(_00128_),
    .B(_00130_),
    .C(_00131_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _06343_ (.A(_00132_),
    .B(_00128_),
    .Y(_00133_));
 sky130_fd_sc_hd__nor2_1 _06344_ (.A(_00122_),
    .B(_00115_),
    .Y(_00134_));
 sky130_fd_sc_hd__a21oi_1 _06345_ (.A1(_00123_),
    .A2(_00133_),
    .B1(_00134_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand2_1 _06346_ (.A(_00111_),
    .B(_00135_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand2_1 _06347_ (.A(_02874_),
    .B(_02522_),
    .Y(_00137_));
 sky130_fd_sc_hd__buf_8 _06348_ (.A(_02797_),
    .X(_00138_));
 sky130_fd_sc_hd__nand2_2 _06349_ (.A(_00138_),
    .B(net64),
    .Y(_00139_));
 sky130_fd_sc_hd__nand2_1 _06350_ (.A(_00137_),
    .B(_00139_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand2_1 _06351_ (.A(_04634_),
    .B(net35),
    .Y(_00141_));
 sky130_fd_sc_hd__inv_2 _06352_ (.A(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__nor2_1 _06353_ (.A(_00137_),
    .B(_00139_),
    .Y(_00143_));
 sky130_fd_sc_hd__a21oi_2 _06354_ (.A1(_00140_),
    .A2(_00142_),
    .B1(_00143_),
    .Y(_00144_));
 sky130_fd_sc_hd__inv_2 _06355_ (.A(_05279_),
    .Y(_00145_));
 sky130_fd_sc_hd__nand2_1 _06356_ (.A(_00145_),
    .B(_05277_),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_2 _06357_ (.A(_05277_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand2_1 _06358_ (.A(_00147_),
    .B(_05279_),
    .Y(_00148_));
 sky130_fd_sc_hd__nand3_1 _06359_ (.A(_00146_),
    .B(_00148_),
    .C(_05281_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand2_1 _06360_ (.A(_00147_),
    .B(_00145_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand3_1 _06361_ (.A(_00150_),
    .B(_05282_),
    .C(_05280_),
    .Y(_00151_));
 sky130_fd_sc_hd__nand2_1 _06362_ (.A(_00149_),
    .B(_00151_),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _06363_ (.A(_00144_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand2_1 _06364_ (.A(_00152_),
    .B(_00153_),
    .Y(_00154_));
 sky130_fd_sc_hd__nand3_1 _06365_ (.A(_00144_),
    .B(_00149_),
    .C(_00151_),
    .Y(_00155_));
 sky130_fd_sc_hd__nand2_1 _06366_ (.A(_00154_),
    .B(_00155_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _06367_ (.A(_05322_),
    .Y(_00157_));
 sky130_fd_sc_hd__o21ai_1 _06368_ (.A1(_05325_),
    .A2(_00157_),
    .B1(_05323_),
    .Y(_00158_));
 sky130_fd_sc_hd__nand3b_1 _06369_ (.A_N(_05325_),
    .B(_05324_),
    .C(_05322_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand2_1 _06370_ (.A(_00158_),
    .B(_00159_),
    .Y(_00160_));
 sky130_fd_sc_hd__inv_2 _06371_ (.A(_00160_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _06372_ (.A(_00156_),
    .B(_00161_),
    .Y(_00162_));
 sky130_fd_sc_hd__o21ai_1 _06373_ (.A1(_00144_),
    .A2(_00152_),
    .B1(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__nor2_1 _06374_ (.A(_00135_),
    .B(_00111_),
    .Y(_00164_));
 sky130_fd_sc_hd__a21oi_1 _06375_ (.A1(_00136_),
    .A2(_00163_),
    .B1(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _06376_ (.A(_00006_),
    .B(_00007_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand2_1 _06377_ (.A(_00166_),
    .B(_05312_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand3b_1 _06378_ (.A_N(_00165_),
    .B(_00008_),
    .C(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _06379_ (.A(_00167_),
    .B(_00008_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand2_1 _06380_ (.A(_00169_),
    .B(_00165_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_1 _06381_ (.A(_00168_),
    .B(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__nand2_1 _06382_ (.A(_05330_),
    .B(_05332_),
    .Y(_00172_));
 sky130_fd_sc_hd__inv_2 _06383_ (.A(_00002_),
    .Y(_00173_));
 sky130_fd_sc_hd__nand2_1 _06384_ (.A(_00172_),
    .B(_00173_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _06385_ (.A(_00174_),
    .B(_00003_),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _06386_ (.A(_05338_),
    .B(_00000_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand2_1 _06387_ (.A(_00176_),
    .B(_05333_),
    .Y(_00177_));
 sky130_fd_sc_hd__nand2_1 _06388_ (.A(_00177_),
    .B(_00001_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _06389_ (.A(_04880_),
    .B(net37),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _06390_ (.A(_04814_),
    .B(_03248_),
    .Y(_00180_));
 sky130_fd_sc_hd__nand2_1 _06391_ (.A(_00179_),
    .B(_00180_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _06392_ (.A(_04895_),
    .B(_04645_),
    .Y(_00182_));
 sky130_fd_sc_hd__inv_2 _06393_ (.A(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__nor2_1 _06394_ (.A(_00179_),
    .B(_00180_),
    .Y(_00184_));
 sky130_fd_sc_hd__a21oi_1 _06395_ (.A1(_00181_),
    .A2(_00183_),
    .B1(_00184_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_1 _06396_ (.A(_00178_),
    .B(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__clkinv_4 _06397_ (.A(_04947_),
    .Y(_00187_));
 sky130_fd_sc_hd__inv_2 _06398_ (.A(_04897_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _06399_ (.A(_04958_),
    .B(_04899_),
    .Y(_00189_));
 sky130_fd_sc_hd__nor3_2 _06400_ (.A(_00187_),
    .B(_00188_),
    .C(_00189_),
    .Y(_00190_));
 sky130_fd_sc_hd__nor2_1 _06401_ (.A(_00185_),
    .B(_00178_),
    .Y(_00191_));
 sky130_fd_sc_hd__a21oi_2 _06402_ (.A1(_00186_),
    .A2(_00190_),
    .B1(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _06403_ (.A(_00175_),
    .B(_00192_),
    .Y(_00193_));
 sky130_fd_sc_hd__buf_6 _06404_ (.A(_04958_),
    .X(_00194_));
 sky130_fd_sc_hd__nand2_1 _06405_ (.A(_00194_),
    .B(_04936_),
    .Y(_00195_));
 sky130_fd_sc_hd__inv_2 _06406_ (.A(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__nor2_1 _06407_ (.A(_00192_),
    .B(_00175_),
    .Y(_00197_));
 sky130_fd_sc_hd__a21oi_1 _06408_ (.A1(_00193_),
    .A2(_00196_),
    .B1(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _06409_ (.A(_00171_),
    .B(_00198_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand3b_1 _06410_ (.A_N(_00198_),
    .B(_00168_),
    .C(_00170_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _06411_ (.A(_00199_),
    .B(_00200_),
    .Y(_00201_));
 sky130_fd_sc_hd__inv_2 _06412_ (.A(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand3_1 _06413_ (.A(_00081_),
    .B(_00037_),
    .C(_00038_),
    .Y(_00203_));
 sky130_fd_sc_hd__a21o_1 _06414_ (.A1(_00047_),
    .A2(_00079_),
    .B1(_00080_),
    .X(_00204_));
 sky130_fd_sc_hd__nand2_1 _06415_ (.A(_00039_),
    .B(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _06416_ (.A(_00203_),
    .B(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _06417_ (.A(_00206_),
    .B(_00029_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand3_1 _06418_ (.A(_00203_),
    .B(_00205_),
    .C(_00028_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _06419_ (.A(_00207_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_2 _06420_ (.A(_00066_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand3_1 _06421_ (.A(_00210_),
    .B(_00058_),
    .C(_00056_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand3_1 _06422_ (.A(_00211_),
    .B(_00067_),
    .C(_00076_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _06423_ (.A(_00212_),
    .B(_00211_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _06424_ (.A(_00051_),
    .B(_00213_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand3_1 _06425_ (.A(_00078_),
    .B(_00033_),
    .C(_00050_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _06426_ (.A(_00214_),
    .B(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _06427_ (.A(_00216_),
    .B(_00047_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand3_1 _06428_ (.A(_00214_),
    .B(_00215_),
    .C(_00046_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _06429_ (.A(_00217_),
    .B(_00218_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _06430_ (.A(_00059_),
    .B(_00210_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand3_1 _06431_ (.A(_00066_),
    .B(_00056_),
    .C(_00058_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand3_1 _06432_ (.A(_00220_),
    .B(_00221_),
    .C(_00075_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _06433_ (.A(_00212_),
    .B(_00222_),
    .Y(_00223_));
 sky130_fd_sc_hd__inv_2 _06434_ (.A(_00061_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _06435_ (.A(_00224_),
    .B(_00060_),
    .Y(_00225_));
 sky130_fd_sc_hd__inv_2 _06436_ (.A(_00060_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _06437_ (.A(_00226_),
    .B(_00061_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand3_1 _06438_ (.A(_00225_),
    .B(_00227_),
    .C(_00063_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _06439_ (.A(_00226_),
    .B(_00224_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand3_1 _06440_ (.A(_00229_),
    .B(_00064_),
    .C(_00062_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _06441_ (.A(_00228_),
    .B(_00230_),
    .Y(_00231_));
 sky130_fd_sc_hd__buf_6 _06442_ (.A(_00344_),
    .X(_00232_));
 sky130_fd_sc_hd__nand2_1 _06443_ (.A(_00232_),
    .B(_02214_),
    .Y(_00233_));
 sky130_fd_sc_hd__buf_6 _06444_ (.A(_00300_),
    .X(_00234_));
 sky130_fd_sc_hd__nand2_1 _06445_ (.A(_00234_),
    .B(_01334_),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_1 _06446_ (.A(_00233_),
    .B(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _06447_ (.A(_00410_),
    .B(_04128_),
    .Y(_00237_));
 sky130_fd_sc_hd__inv_2 _06448_ (.A(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__nor2_1 _06449_ (.A(_00233_),
    .B(_00235_),
    .Y(_00239_));
 sky130_fd_sc_hd__a21oi_1 _06450_ (.A1(_00236_),
    .A2(_00238_),
    .B1(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _06451_ (.A(_00231_),
    .B(_00240_),
    .Y(_00241_));
 sky130_fd_sc_hd__inv_2 _06452_ (.A(_00117_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _06453_ (.A(_00242_),
    .B(_00116_),
    .Y(_00243_));
 sky130_fd_sc_hd__inv_2 _06454_ (.A(_00116_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _06455_ (.A(_00244_),
    .B(_00117_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand3_1 _06456_ (.A(_00243_),
    .B(_00245_),
    .C(_00119_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _06457_ (.A(_00244_),
    .B(_00242_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand3_1 _06458_ (.A(_00247_),
    .B(_00120_),
    .C(_00118_),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _06459_ (.A(_00246_),
    .B(_00248_),
    .Y(_00249_));
 sky130_fd_sc_hd__inv_2 _06460_ (.A(_00249_),
    .Y(_00250_));
 sky130_fd_sc_hd__nor2_1 _06461_ (.A(_00240_),
    .B(_00231_),
    .Y(_00251_));
 sky130_fd_sc_hd__a21oi_1 _06462_ (.A1(_00241_),
    .A2(_00250_),
    .B1(_00251_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _06463_ (.A(_00223_),
    .B(_00252_),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_2 _06464_ (.A(_00122_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _06465_ (.A(_00115_),
    .B(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand3_1 _06466_ (.A(_00122_),
    .B(_00114_),
    .C(_05272_),
    .Y(_00256_));
 sky130_fd_sc_hd__nand2_1 _06467_ (.A(_00255_),
    .B(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _06468_ (.A(_00257_),
    .B(_00133_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand3b_1 _06469_ (.A_N(_00133_),
    .B(_00255_),
    .C(_00256_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _06470_ (.A(_00258_),
    .B(_00259_),
    .Y(_00260_));
 sky130_fd_sc_hd__inv_2 _06471_ (.A(_00260_),
    .Y(_00261_));
 sky130_fd_sc_hd__nor2_1 _06472_ (.A(_00252_),
    .B(_00223_),
    .Y(_00262_));
 sky130_fd_sc_hd__a21oi_1 _06473_ (.A1(_00253_),
    .A2(_00261_),
    .B1(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _06474_ (.A(_00219_),
    .B(_00263_),
    .Y(_00264_));
 sky130_fd_sc_hd__a21o_1 _06475_ (.A1(_00123_),
    .A2(_00133_),
    .B1(_00134_),
    .X(_00265_));
 sky130_fd_sc_hd__nand2_1 _06476_ (.A(_00111_),
    .B(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand3_1 _06477_ (.A(_00135_),
    .B(_05302_),
    .C(_00110_),
    .Y(_00267_));
 sky130_fd_sc_hd__nand3b_1 _06478_ (.A_N(_00163_),
    .B(_00266_),
    .C(_00267_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _06479_ (.A(_00267_),
    .B(_00266_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _06480_ (.A(_00269_),
    .B(_00163_),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _06481_ (.A(_00268_),
    .B(_00270_),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _06482_ (.A(_00271_),
    .Y(_00272_));
 sky130_fd_sc_hd__nor2_1 _06483_ (.A(_00263_),
    .B(_00219_),
    .Y(_00273_));
 sky130_fd_sc_hd__a21oi_2 _06484_ (.A1(_00264_),
    .A2(_00272_),
    .B1(_00273_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _06485_ (.A(_00209_),
    .B(_00274_),
    .Y(_00275_));
 sky130_fd_sc_hd__nor2_1 _06486_ (.A(_00274_),
    .B(_00209_),
    .Y(_00276_));
 sky130_fd_sc_hd__a21oi_2 _06487_ (.A1(_00202_),
    .A2(_00275_),
    .B1(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _06488_ (.A(_00109_),
    .B(_00277_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _06489_ (.A(_00200_),
    .B(_00168_),
    .Y(_00279_));
 sky130_fd_sc_hd__nor2_1 _06490_ (.A(_00277_),
    .B(_00109_),
    .Y(_00280_));
 sky130_fd_sc_hd__a21oi_1 _06491_ (.A1(_00278_),
    .A2(_00279_),
    .B1(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _06492_ (.A(_00281_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand3_1 _06493_ (.A(_00087_),
    .B(_05239_),
    .C(_05240_),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _06494_ (.A(_00087_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _06495_ (.A(_00284_),
    .B(_05241_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _06496_ (.A(_00283_),
    .B(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _06497_ (.A(_00286_),
    .B(_00093_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand3b_1 _06498_ (.A_N(_00093_),
    .B(_00283_),
    .C(_00285_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand3_2 _06499_ (.A(_00282_),
    .B(_00287_),
    .C(_00288_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _06500_ (.A(_00102_),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__inv_2 _06501_ (.A(_00289_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand3_4 _06502_ (.A(_00100_),
    .B(_00101_),
    .C(_00291_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _06503_ (.A(_00290_),
    .B(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand3_1 _06504_ (.A(_00154_),
    .B(_00155_),
    .C(_00160_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _06505_ (.A(_00162_),
    .B(_00294_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _06506_ (.A(_00127_),
    .B(_00124_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _06507_ (.A(_00125_),
    .B(_00126_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand3_1 _06508_ (.A(_00296_),
    .B(_00297_),
    .C(_00129_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _06509_ (.A(_00298_),
    .B(_00132_),
    .Y(_00299_));
 sky130_fd_sc_hd__buf_6 _06510_ (.A(_00641_),
    .X(_00301_));
 sky130_fd_sc_hd__nand2_1 _06511_ (.A(_01532_),
    .B(_00301_),
    .Y(_00302_));
 sky130_fd_sc_hd__buf_6 _06512_ (.A(_00674_),
    .X(_00303_));
 sky130_fd_sc_hd__nand2_1 _06513_ (.A(_00303_),
    .B(_00960_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _06514_ (.A(_00302_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__clkbuf_8 _06515_ (.A(_00751_),
    .X(_00306_));
 sky130_fd_sc_hd__nand2_1 _06516_ (.A(_03105_),
    .B(_00306_),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _06517_ (.A(_00307_),
    .Y(_00308_));
 sky130_fd_sc_hd__nor2_1 _06518_ (.A(_00302_),
    .B(_00304_),
    .Y(_00309_));
 sky130_fd_sc_hd__a21oi_1 _06519_ (.A1(_00305_),
    .A2(_00308_),
    .B1(_00309_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _06520_ (.A(_00299_),
    .B(_00310_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _06521_ (.A(_05113_),
    .B(_05068_),
    .Y(_00313_));
 sky130_fd_sc_hd__inv_2 _06522_ (.A(_00313_),
    .Y(_00314_));
 sky130_fd_sc_hd__buf_6 _06523_ (.A(_01224_),
    .X(_00315_));
 sky130_fd_sc_hd__nand2_1 _06524_ (.A(_05278_),
    .B(_00315_),
    .Y(_00316_));
 sky130_fd_sc_hd__inv_2 _06525_ (.A(_00316_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _06526_ (.A(_00314_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_1 _06527_ (.A(_00138_),
    .B(_02203_),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _06528_ (.A(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _06529_ (.A(_00313_),
    .B(_00316_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand3_1 _06530_ (.A(_00318_),
    .B(_00320_),
    .C(_00321_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _06531_ (.A(_00323_),
    .B(_00318_),
    .Y(_00324_));
 sky130_fd_sc_hd__nor2_1 _06532_ (.A(_00310_),
    .B(_00299_),
    .Y(_00325_));
 sky130_fd_sc_hd__a21oi_1 _06533_ (.A1(_00312_),
    .A2(_00324_),
    .B1(_00325_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _06534_ (.A(_00295_),
    .B(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _06535_ (.A(_04634_),
    .B(_02522_),
    .Y(_00328_));
 sky130_fd_sc_hd__buf_8 _06536_ (.A(_02874_),
    .X(_00329_));
 sky130_fd_sc_hd__nand2_1 _06537_ (.A(_00329_),
    .B(_03039_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _06538_ (.A(_00328_),
    .B(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _06539_ (.A(_04814_),
    .B(net35),
    .Y(_00332_));
 sky130_fd_sc_hd__inv_2 _06540_ (.A(_00332_),
    .Y(_00334_));
 sky130_fd_sc_hd__nor2_1 _06541_ (.A(_00328_),
    .B(_00330_),
    .Y(_00335_));
 sky130_fd_sc_hd__a21oi_2 _06542_ (.A1(_00331_),
    .A2(_00334_),
    .B1(_00335_),
    .Y(_00336_));
 sky130_fd_sc_hd__inv_2 _06543_ (.A(_00137_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _06544_ (.A(_00337_),
    .B(_00139_),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_2 _06545_ (.A(_00139_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _06546_ (.A(_00339_),
    .B(_00137_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand3_1 _06547_ (.A(_00338_),
    .B(_00340_),
    .C(_00141_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _06548_ (.A(_00337_),
    .B(_00339_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand3_1 _06549_ (.A(_00342_),
    .B(_00142_),
    .C(_00140_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _06550_ (.A(_00341_),
    .B(_00343_),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_2 _06551_ (.A(_00336_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _06552_ (.A(_00345_),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand3_1 _06553_ (.A(_00336_),
    .B(_00341_),
    .C(_00343_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _06554_ (.A(_00347_),
    .B(_00348_),
    .Y(_00349_));
 sky130_fd_sc_hd__inv_2 _06555_ (.A(_00181_),
    .Y(_00350_));
 sky130_fd_sc_hd__o21ai_1 _06556_ (.A1(_00184_),
    .A2(_00350_),
    .B1(_00182_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand3b_1 _06557_ (.A_N(_00184_),
    .B(_00183_),
    .C(_00181_),
    .Y(_00352_));
 sky130_fd_sc_hd__nand2_1 _06558_ (.A(_00351_),
    .B(_00352_),
    .Y(_00353_));
 sky130_fd_sc_hd__inv_2 _06559_ (.A(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _06560_ (.A(_00349_),
    .B(_00354_),
    .Y(_00356_));
 sky130_fd_sc_hd__o21ai_2 _06561_ (.A1(_00336_),
    .A2(_00345_),
    .B1(_00356_),
    .Y(_00357_));
 sky130_fd_sc_hd__nor2_1 _06562_ (.A(_00326_),
    .B(_00295_),
    .Y(_00358_));
 sky130_fd_sc_hd__a21oi_1 _06563_ (.A1(_00327_),
    .A2(_00357_),
    .B1(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__inv_2 _06564_ (.A(_00359_),
    .Y(_00360_));
 sky130_fd_sc_hd__inv_2 _06565_ (.A(_00192_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_1 _06566_ (.A(_00175_),
    .B(_00361_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand3_1 _06567_ (.A(_00192_),
    .B(_00174_),
    .C(_00003_),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_1 _06568_ (.A(_00362_),
    .B(_00363_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand2_1 _06569_ (.A(_00364_),
    .B(_00196_),
    .Y(_00365_));
 sky130_fd_sc_hd__nand3_1 _06570_ (.A(_00362_),
    .B(_00363_),
    .C(_00195_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand3_1 _06571_ (.A(_00360_),
    .B(_00365_),
    .C(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__nand2_1 _06572_ (.A(_00365_),
    .B(_00367_),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _06573_ (.A(_00369_),
    .B(_00359_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand2_1 _06574_ (.A(_00368_),
    .B(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_2 _06575_ (.A(_00191_),
    .Y(_00372_));
 sky130_fd_sc_hd__nand2_1 _06576_ (.A(_00372_),
    .B(_00186_),
    .Y(_00373_));
 sky130_fd_sc_hd__inv_2 _06577_ (.A(_00190_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(_00373_),
    .B(_00374_),
    .Y(_00375_));
 sky130_fd_sc_hd__nand3_1 _06579_ (.A(_00372_),
    .B(_00190_),
    .C(_00186_),
    .Y(_00376_));
 sky130_fd_sc_hd__o21ai_1 _06580_ (.A1(_00187_),
    .A2(_00188_),
    .B1(_00189_),
    .Y(_00378_));
 sky130_fd_sc_hd__nand2_1 _06581_ (.A(_00374_),
    .B(_00378_),
    .Y(_00379_));
 sky130_fd_sc_hd__nand2_1 _06582_ (.A(_05310_),
    .B(_04645_),
    .Y(_00380_));
 sky130_fd_sc_hd__buf_8 _06583_ (.A(_04895_),
    .X(_00381_));
 sky130_fd_sc_hd__nand2_1 _06584_ (.A(_00381_),
    .B(_05114_),
    .Y(_00382_));
 sky130_fd_sc_hd__inv_2 _06585_ (.A(_00382_),
    .Y(_00383_));
 sky130_fd_sc_hd__buf_12 _06586_ (.A(_04880_),
    .X(_00384_));
 sky130_fd_sc_hd__nand2_1 _06587_ (.A(_00384_),
    .B(_03248_),
    .Y(_00385_));
 sky130_fd_sc_hd__inv_2 _06588_ (.A(_00385_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _06589_ (.A(_00383_),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _06590_ (.A(_00382_),
    .B(_00385_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand3b_1 _06591_ (.A_N(_00380_),
    .B(_00387_),
    .C(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__and2_1 _06592_ (.A(_00390_),
    .B(_00387_),
    .X(_00391_));
 sky130_fd_sc_hd__nor2_1 _06593_ (.A(_00379_),
    .B(_00391_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand3_1 _06594_ (.A(_00375_),
    .B(_00376_),
    .C(_00392_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _06595_ (.A(_00371_),
    .B(_00393_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand3b_1 _06596_ (.A_N(_00393_),
    .B(_00368_),
    .C(_00370_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _06597_ (.A(_00394_),
    .B(_00395_),
    .Y(_00396_));
 sky130_fd_sc_hd__a21o_1 _06598_ (.A1(_00253_),
    .A2(_00261_),
    .B1(_00262_),
    .X(_00397_));
 sky130_fd_sc_hd__nand3_1 _06599_ (.A(_00397_),
    .B(_00217_),
    .C(_00218_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand3_1 _06600_ (.A(_00398_),
    .B(_00272_),
    .C(_00264_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _06601_ (.A(_00219_),
    .B(_00397_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand3_1 _06602_ (.A(_00263_),
    .B(_00217_),
    .C(_00218_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand3_1 _06603_ (.A(_00401_),
    .B(_00402_),
    .C(_00271_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _06604_ (.A(_00400_),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__nand3_1 _06605_ (.A(_00252_),
    .B(_00212_),
    .C(_00222_),
    .Y(_00405_));
 sky130_fd_sc_hd__a21o_1 _06606_ (.A1(_00236_),
    .A2(_00238_),
    .B1(_00239_),
    .X(_00406_));
 sky130_fd_sc_hd__nand3_1 _06607_ (.A(_00406_),
    .B(_00230_),
    .C(_00228_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand3_1 _06608_ (.A(_00407_),
    .B(_00241_),
    .C(_00250_),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _06609_ (.A(_00408_),
    .B(_00407_),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _06610_ (.A(_00223_),
    .B(_00409_),
    .Y(_00411_));
 sky130_fd_sc_hd__nand2_1 _06611_ (.A(_00405_),
    .B(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _06612_ (.A(_00412_),
    .B(_00261_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand3_2 _06613_ (.A(_00405_),
    .B(_00411_),
    .C(_00260_),
    .Y(_00414_));
 sky130_fd_sc_hd__nand2_1 _06614_ (.A(_00413_),
    .B(_00414_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _06615_ (.A(_00231_),
    .B(_00406_),
    .Y(_00416_));
 sky130_fd_sc_hd__nand3_1 _06616_ (.A(_00240_),
    .B(_00228_),
    .C(_00230_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand3_1 _06617_ (.A(_00416_),
    .B(_00417_),
    .C(_00249_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _06618_ (.A(_00408_),
    .B(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__inv_2 _06619_ (.A(_00235_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _06620_ (.A(_00420_),
    .B(_00233_),
    .Y(_00422_));
 sky130_fd_sc_hd__inv_2 _06621_ (.A(_00233_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _06622_ (.A(_00423_),
    .B(_00235_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand3_1 _06623_ (.A(_00422_),
    .B(_00424_),
    .C(_00237_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _06624_ (.A(_00423_),
    .B(_00420_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand3_1 _06625_ (.A(_00426_),
    .B(_00238_),
    .C(_00236_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _06626_ (.A(_00425_),
    .B(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _06627_ (.A(_00344_),
    .B(_01334_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _06628_ (.A(_00300_),
    .B(_01532_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _06629_ (.A(_00429_),
    .B(_00430_),
    .Y(_00431_));
 sky130_fd_sc_hd__buf_6 _06630_ (.A(_00410_),
    .X(_00433_));
 sky130_fd_sc_hd__nand2_1 _06631_ (.A(_00433_),
    .B(_02214_),
    .Y(_00434_));
 sky130_fd_sc_hd__inv_2 _06632_ (.A(_00434_),
    .Y(_00435_));
 sky130_fd_sc_hd__nor2_1 _06633_ (.A(_00429_),
    .B(_00430_),
    .Y(_00436_));
 sky130_fd_sc_hd__a21oi_1 _06634_ (.A1(_00431_),
    .A2(_00435_),
    .B1(_00436_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _06635_ (.A(_00428_),
    .B(_00437_),
    .Y(_00438_));
 sky130_fd_sc_hd__inv_2 _06636_ (.A(_00304_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _06637_ (.A(_00439_),
    .B(_00302_),
    .Y(_00440_));
 sky130_fd_sc_hd__inv_2 _06638_ (.A(_00302_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _06639_ (.A(_00441_),
    .B(_00304_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand3_1 _06640_ (.A(_00440_),
    .B(_00442_),
    .C(_00307_),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _06641_ (.A(_00441_),
    .B(_00439_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand3_1 _06642_ (.A(_00445_),
    .B(_00308_),
    .C(_00305_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _06643_ (.A(_00444_),
    .B(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__inv_2 _06644_ (.A(_00447_),
    .Y(_00448_));
 sky130_fd_sc_hd__nor2_1 _06645_ (.A(_00437_),
    .B(_00428_),
    .Y(_00449_));
 sky130_fd_sc_hd__a21oi_1 _06646_ (.A1(_00438_),
    .A2(_00448_),
    .B1(_00449_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _06647_ (.A(_00419_),
    .B(_00450_),
    .Y(_00451_));
 sky130_fd_sc_hd__a21o_1 _06648_ (.A1(_00305_),
    .A2(_00308_),
    .B1(_00309_),
    .X(_00452_));
 sky130_fd_sc_hd__nand2_1 _06649_ (.A(_00299_),
    .B(_00452_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand3_1 _06650_ (.A(_00310_),
    .B(_00298_),
    .C(_00132_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand3b_1 _06651_ (.A_N(_00324_),
    .B(_00453_),
    .C(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand3_1 _06652_ (.A(_00452_),
    .B(_00132_),
    .C(_00298_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand3_1 _06653_ (.A(_00457_),
    .B(_00312_),
    .C(_00324_),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _06654_ (.A(_00456_),
    .B(_00458_),
    .Y(_00459_));
 sky130_fd_sc_hd__inv_2 _06655_ (.A(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__nor2_1 _06656_ (.A(_00450_),
    .B(_00419_),
    .Y(_00461_));
 sky130_fd_sc_hd__a21oi_1 _06657_ (.A1(_00451_),
    .A2(_00460_),
    .B1(_00461_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _06658_ (.A(_00415_),
    .B(_00462_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand3_1 _06659_ (.A(_00326_),
    .B(_00162_),
    .C(_00294_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _06660_ (.A(_00458_),
    .B(_00457_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _06661_ (.A(_00295_),
    .B(_00466_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _06662_ (.A(_00464_),
    .B(_00467_),
    .Y(_00468_));
 sky130_fd_sc_hd__nand2_1 _06663_ (.A(_00468_),
    .B(_00357_),
    .Y(_00469_));
 sky130_fd_sc_hd__inv_2 _06664_ (.A(_00357_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand3_1 _06665_ (.A(_00470_),
    .B(_00464_),
    .C(_00467_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _06666_ (.A(_00469_),
    .B(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__inv_2 _06667_ (.A(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2_1 _06668_ (.A(_00462_),
    .B(_00415_),
    .Y(_00474_));
 sky130_fd_sc_hd__a21oi_1 _06669_ (.A1(_00463_),
    .A2(_00473_),
    .B1(_00474_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _06670_ (.A(_00404_),
    .B(_00475_),
    .Y(_00477_));
 sky130_fd_sc_hd__inv_2 _06671_ (.A(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__nor2_1 _06672_ (.A(_00475_),
    .B(_00404_),
    .Y(_00479_));
 sky130_fd_sc_hd__o21bai_1 _06673_ (.A1(_00396_),
    .A2(_00478_),
    .B1_N(_00479_),
    .Y(_00480_));
 sky130_fd_sc_hd__inv_2 _06674_ (.A(_00274_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _06675_ (.A(_00209_),
    .B(_00481_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand3_1 _06676_ (.A(_00274_),
    .B(_00207_),
    .C(_00208_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _06677_ (.A(_00482_),
    .B(_00483_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _06678_ (.A(_00484_),
    .B(_00202_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand3_1 _06679_ (.A(_00482_),
    .B(_00483_),
    .C(_00201_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand3_1 _06680_ (.A(_00480_),
    .B(_00485_),
    .C(_00486_),
    .Y(_00488_));
 sky130_fd_sc_hd__nand2_1 _06681_ (.A(_00485_),
    .B(_00486_),
    .Y(_00489_));
 sky130_fd_sc_hd__inv_2 _06682_ (.A(_00396_),
    .Y(_00490_));
 sky130_fd_sc_hd__a21oi_1 _06683_ (.A1(_00490_),
    .A2(_00477_),
    .B1(_00479_),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _06684_ (.A(_00489_),
    .B(_00491_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _06685_ (.A(_00395_),
    .B(_00368_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand3_1 _06686_ (.A(_00488_),
    .B(_00492_),
    .C(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _06687_ (.A(_00494_),
    .B(_00488_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand3_1 _06688_ (.A(_00277_),
    .B(_00107_),
    .C(_00108_),
    .Y(_00496_));
 sky130_fd_sc_hd__inv_2 _06689_ (.A(_00277_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _06690_ (.A(_00497_),
    .B(_00109_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _06691_ (.A(_00496_),
    .B(_00499_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _06692_ (.A(_00500_),
    .B(_00279_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand3b_1 _06693_ (.A_N(_00279_),
    .B(_00496_),
    .C(_00499_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand3_2 _06694_ (.A(_00495_),
    .B(_00501_),
    .C(_00502_),
    .Y(_00503_));
 sky130_fd_sc_hd__inv_2 _06695_ (.A(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _06696_ (.A(_00287_),
    .B(_00288_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _06697_ (.A(_00505_),
    .B(_00281_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand3_1 _06698_ (.A(_00504_),
    .B(_00289_),
    .C(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(_00293_),
    .B(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__inv_2 _06700_ (.A(_00507_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand3_2 _06701_ (.A(_00290_),
    .B(_00292_),
    .C(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _06702_ (.A(_00508_),
    .B(_00511_),
    .Y(_00512_));
 sky130_fd_sc_hd__inv_2 _06703_ (.A(_00512_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(_05234_),
    .B(_00097_),
    .Y(_00514_));
 sky130_fd_sc_hd__nor2_1 _06705_ (.A(_00097_),
    .B(_05234_),
    .Y(_00515_));
 sky130_fd_sc_hd__a21o_1 _06706_ (.A1(_00514_),
    .A2(_00091_),
    .B1(_00515_),
    .X(_00516_));
 sky130_fd_sc_hd__nand2_1 _06707_ (.A(_05063_),
    .B(_05028_),
    .Y(_00517_));
 sky130_fd_sc_hd__nor2_1 _06708_ (.A(_05028_),
    .B(_05063_),
    .Y(_00518_));
 sky130_fd_sc_hd__a21o_1 _06709_ (.A1(_05088_),
    .A2(_00517_),
    .B1(_00518_),
    .X(_00519_));
 sky130_fd_sc_hd__nand2_1 _06710_ (.A(_05041_),
    .B(_05043_),
    .Y(_00521_));
 sky130_fd_sc_hd__nor2_1 _06711_ (.A(_05043_),
    .B(_05041_),
    .Y(_00522_));
 sky130_fd_sc_hd__a21oi_1 _06712_ (.A1(_05060_),
    .A2(_00521_),
    .B1(_00522_),
    .Y(_00523_));
 sky130_fd_sc_hd__inv_2 _06713_ (.A(_00523_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(_00641_),
    .B(_00421_),
    .Y(_00525_));
 sky130_fd_sc_hd__clkbuf_4 _06715_ (.A(net16),
    .X(_00526_));
 sky130_fd_sc_hd__nand2_1 _06716_ (.A(_00303_),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__or2_1 _06717_ (.A(_00525_),
    .B(_00527_),
    .X(_00528_));
 sky130_fd_sc_hd__nand2_1 _06718_ (.A(_00525_),
    .B(_00527_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _06719_ (.A(_00528_),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _06720_ (.A(_00306_),
    .B(_00355_),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _06721_ (.A(_00530_),
    .B(_00532_),
    .Y(_00533_));
 sky130_fd_sc_hd__inv_2 _06722_ (.A(_00532_),
    .Y(_00534_));
 sky130_fd_sc_hd__nand3_1 _06723_ (.A(_00528_),
    .B(_00534_),
    .C(_00529_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _06724_ (.A(_00533_),
    .B(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _06725_ (.A(_00344_),
    .B(_01895_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _06726_ (.A(_00234_),
    .B(_00685_),
    .Y(_00538_));
 sky130_fd_sc_hd__or2_1 _06727_ (.A(_00537_),
    .B(_00538_),
    .X(_00539_));
 sky130_fd_sc_hd__nand2_1 _06728_ (.A(_00537_),
    .B(_00538_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _06729_ (.A(_00539_),
    .B(_00540_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _06730_ (.A(_00433_),
    .B(_05049_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _06731_ (.A(_00541_),
    .B(_00543_),
    .Y(_00544_));
 sky130_fd_sc_hd__nand3b_2 _06732_ (.A_N(_00543_),
    .B(_00539_),
    .C(_00540_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _06733_ (.A(_00544_),
    .B(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _06734_ (.A(_05040_),
    .B(_05034_),
    .Y(_00547_));
 sky130_fd_sc_hd__inv_2 _06735_ (.A(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _06736_ (.A(_00546_),
    .B(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand3_2 _06737_ (.A(_00547_),
    .B(_00544_),
    .C(_00545_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand3b_2 _06738_ (.A_N(_00536_),
    .B(_00549_),
    .C(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _06739_ (.A(_00549_),
    .B(_00550_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _06740_ (.A(_00552_),
    .B(_00536_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand3_1 _06741_ (.A(_00524_),
    .B(_00551_),
    .C(_00554_),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _06742_ (.A(_00554_),
    .B(_00551_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand2_1 _06743_ (.A(_00556_),
    .B(_00523_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _06744_ (.A(_00315_),
    .B(_00520_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand3b_1 _06745_ (.A_N(_00558_),
    .B(_05068_),
    .C(_00311_),
    .Y(_00559_));
 sky130_fd_sc_hd__inv_2 _06746_ (.A(_01257_),
    .Y(_00560_));
 sky130_fd_sc_hd__inv_2 _06747_ (.A(_00311_),
    .Y(_00561_));
 sky130_fd_sc_hd__o21ai_1 _06748_ (.A1(_00560_),
    .A2(_00561_),
    .B1(_00558_),
    .Y(_00562_));
 sky130_fd_sc_hd__nand2_1 _06749_ (.A(_00559_),
    .B(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _06750_ (.A(_02203_),
    .B(_00960_),
    .Y(_00565_));
 sky130_fd_sc_hd__nand2_1 _06751_ (.A(_00563_),
    .B(_00565_),
    .Y(_00566_));
 sky130_fd_sc_hd__inv_2 _06752_ (.A(_00565_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand3_1 _06753_ (.A(_00559_),
    .B(_00562_),
    .C(_00567_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _06754_ (.A(_00566_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _06755_ (.A(_05058_),
    .B(_05052_),
    .Y(_00570_));
 sky130_fd_sc_hd__inv_2 _06756_ (.A(_00570_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _06757_ (.A(_00569_),
    .B(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand3_1 _06758_ (.A(_00570_),
    .B(_00566_),
    .C(_00568_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _06759_ (.A(_00572_),
    .B(_00573_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _06760_ (.A(_05075_),
    .B(_05070_),
    .Y(_00576_));
 sky130_fd_sc_hd__inv_2 _06761_ (.A(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _06762_ (.A(_00574_),
    .B(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand3_1 _06763_ (.A(_00572_),
    .B(_00573_),
    .C(_00576_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _06764_ (.A(_00578_),
    .B(_00579_),
    .Y(_00580_));
 sky130_fd_sc_hd__inv_2 _06765_ (.A(_00580_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand3_2 _06766_ (.A(_00555_),
    .B(_00557_),
    .C(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _06767_ (.A(_00556_),
    .B(_00524_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand3_1 _06768_ (.A(_00523_),
    .B(_00554_),
    .C(_00551_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand3_1 _06769_ (.A(_00583_),
    .B(_00584_),
    .C(_00580_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand3_1 _06770_ (.A(_00519_),
    .B(_00582_),
    .C(_00585_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_1 _06771_ (.A(_00582_),
    .B(_00585_),
    .Y(_00588_));
 sky130_fd_sc_hd__a21oi_1 _06772_ (.A1(_05088_),
    .A2(_00517_),
    .B1(_00518_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _06773_ (.A(_00588_),
    .B(_00589_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(_03105_),
    .B(_05114_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand2_1 _06775_ (.A(_01532_),
    .B(_03248_),
    .Y(_00592_));
 sky130_fd_sc_hd__or2_1 _06776_ (.A(_00591_),
    .B(_00592_),
    .X(_00593_));
 sky130_fd_sc_hd__nand2_1 _06777_ (.A(_00591_),
    .B(_00592_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _06778_ (.A(_00593_),
    .B(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _06779_ (.A(_05113_),
    .B(_04645_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _06780_ (.A(_00595_),
    .B(_00596_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand3b_1 _06781_ (.A_N(_00596_),
    .B(_00593_),
    .C(_00594_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _06782_ (.A(_00598_),
    .B(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(_05096_),
    .B(_02214_),
    .Y(_00601_));
 sky130_fd_sc_hd__inv_2 _06784_ (.A(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _06785_ (.A(_03039_),
    .B(_04128_),
    .Y(_00603_));
 sky130_fd_sc_hd__inv_2 _06786_ (.A(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _06787_ (.A(_00602_),
    .B(_00604_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _06788_ (.A(_00601_),
    .B(_00603_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _06789_ (.A(_02687_),
    .B(_01334_),
    .Y(_00607_));
 sky130_fd_sc_hd__inv_2 _06790_ (.A(_00607_),
    .Y(_00609_));
 sky130_fd_sc_hd__a21o_1 _06791_ (.A1(_00605_),
    .A2(_00606_),
    .B1(_00609_),
    .X(_00610_));
 sky130_fd_sc_hd__nand3_2 _06792_ (.A(_00605_),
    .B(_00609_),
    .C(_00606_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(_00610_),
    .B(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__a21boi_1 _06794_ (.A1(_05106_),
    .A2(_05102_),
    .B1_N(_05101_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(_00612_),
    .B(_00613_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _06796_ (.A(_05107_),
    .B(_05101_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand3_1 _06797_ (.A(_00610_),
    .B(_00615_),
    .C(_00611_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand3b_1 _06798_ (.A_N(_00600_),
    .B(_00614_),
    .C(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _06799_ (.A(_00612_),
    .B(_00615_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand3_1 _06800_ (.A(_00610_),
    .B(_00613_),
    .C(_00611_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand3_1 _06801_ (.A(_00618_),
    .B(_00620_),
    .C(_00600_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _06802_ (.A(_00617_),
    .B(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _06803_ (.A(_05076_),
    .B(_05078_),
    .Y(_00623_));
 sky130_fd_sc_hd__nor2_1 _06804_ (.A(_05078_),
    .B(_05076_),
    .Y(_00624_));
 sky130_fd_sc_hd__a21oi_2 _06805_ (.A1(_00623_),
    .A2(_05083_),
    .B1(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__inv_2 _06806_ (.A(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _06807_ (.A(_00622_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand3_1 _06808_ (.A(_00625_),
    .B(_00617_),
    .C(_00621_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _06809_ (.A(_00627_),
    .B(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _06810_ (.A(_05127_),
    .B(_05108_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(_00629_),
    .B(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand3b_1 _06812_ (.A_N(_00631_),
    .B(_00627_),
    .C(_00628_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _06813_ (.A(_00632_),
    .B(_00633_),
    .Y(_00634_));
 sky130_fd_sc_hd__inv_2 _06814_ (.A(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand3_2 _06815_ (.A(_00587_),
    .B(_00590_),
    .C(_00635_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _06816_ (.A(_00588_),
    .B(_00519_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand3_1 _06817_ (.A(_00589_),
    .B(_00582_),
    .C(_00585_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand3_1 _06818_ (.A(_00637_),
    .B(_00638_),
    .C(_00634_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2_1 _06819_ (.A(_00636_),
    .B(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _06820_ (.A(_05091_),
    .B(_05024_),
    .Y(_00642_));
 sky130_fd_sc_hd__nor2_1 _06821_ (.A(_05024_),
    .B(_05091_),
    .Y(_00643_));
 sky130_fd_sc_hd__a21o_1 _06822_ (.A1(_00642_),
    .A2(_05140_),
    .B1(_00643_),
    .X(_00644_));
 sky130_fd_sc_hd__nand2_1 _06823_ (.A(_00640_),
    .B(_00644_),
    .Y(_00645_));
 sky130_fd_sc_hd__a21oi_1 _06824_ (.A1(_00642_),
    .A2(_05140_),
    .B1(_00643_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand3_1 _06825_ (.A(_00646_),
    .B(_00636_),
    .C(_00639_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_1 _06826_ (.A(_00645_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _06827_ (.A(_00138_),
    .B(_04899_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_1 _06828_ (.A(_05278_),
    .B(_04897_),
    .Y(_00650_));
 sky130_fd_sc_hd__or2_1 _06829_ (.A(_00649_),
    .B(_00650_),
    .X(_00651_));
 sky130_fd_sc_hd__nand2_1 _06830_ (.A(_00649_),
    .B(_00650_),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _06831_ (.A(_00651_),
    .B(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _06832_ (.A(_00329_),
    .B(_04888_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand2_1 _06833_ (.A(_00654_),
    .B(_00655_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand3b_1 _06834_ (.A_N(_00655_),
    .B(_00651_),
    .C(_00653_),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_00656_),
    .B(_00657_),
    .Y(_00658_));
 sky130_fd_sc_hd__a21oi_2 _06836_ (.A1(_05119_),
    .A2(_05123_),
    .B1(_05117_),
    .Y(_00659_));
 sky130_fd_sc_hd__inv_2 _06837_ (.A(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_00658_),
    .B(_00660_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand3_1 _06839_ (.A(_00656_),
    .B(_00657_),
    .C(_00659_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(_00661_),
    .B(_00662_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand2_1 _06841_ (.A(_05162_),
    .B(_05156_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _06842_ (.A(_00664_),
    .B(_00665_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand3b_1 _06843_ (.A_N(_00665_),
    .B(_00661_),
    .C(_00662_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _06844_ (.A(_00666_),
    .B(_00667_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand2_1 _06845_ (.A(_05163_),
    .B(_05164_),
    .Y(_00669_));
 sky130_fd_sc_hd__nor2_1 _06846_ (.A(_05164_),
    .B(_05163_),
    .Y(_00670_));
 sky130_fd_sc_hd__a21oi_2 _06847_ (.A1(_00669_),
    .A2(_05169_),
    .B1(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__inv_2 _06848_ (.A(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(_00668_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand3_1 _06850_ (.A(_00666_),
    .B(_00667_),
    .C(_00671_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_1 _06851_ (.A(_00673_),
    .B(_00675_),
    .Y(_00676_));
 sky130_fd_sc_hd__nand2_1 _06852_ (.A(_05191_),
    .B(_04947_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(net46),
    .B(_04895_),
    .Y(_00678_));
 sky130_fd_sc_hd__or2_1 _06854_ (.A(_00677_),
    .B(_00678_),
    .X(_00679_));
 sky130_fd_sc_hd__nand2_1 _06855_ (.A(_00677_),
    .B(_00678_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _06856_ (.A(_00679_),
    .B(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__buf_4 _06857_ (.A(net48),
    .X(_00682_));
 sky130_fd_sc_hd__nand3b_1 _06858_ (.A_N(_00681_),
    .B(_00682_),
    .C(_04958_),
    .Y(_00683_));
 sky130_fd_sc_hd__nand2_1 _06859_ (.A(_00682_),
    .B(_04958_),
    .Y(_00684_));
 sky130_fd_sc_hd__nand2_1 _06860_ (.A(_00681_),
    .B(_00684_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand2_1 _06861_ (.A(_00683_),
    .B(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(_00384_),
    .B(_04941_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _06863_ (.A(_04814_),
    .B(_04933_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(_04634_),
    .B(_04936_),
    .Y(_00690_));
 sky130_fd_sc_hd__or2_1 _06865_ (.A(_00689_),
    .B(_00690_),
    .X(_00691_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(_00689_),
    .B(_00690_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _06867_ (.A(_00691_),
    .B(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__or2_1 _06868_ (.A(_00688_),
    .B(_00693_),
    .X(_00694_));
 sky130_fd_sc_hd__nand2_1 _06869_ (.A(_05184_),
    .B(_05177_),
    .Y(_00695_));
 sky130_fd_sc_hd__nand2_1 _06870_ (.A(_00693_),
    .B(_00688_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand3_1 _06871_ (.A(_00694_),
    .B(_00695_),
    .C(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _06872_ (.A(_00694_),
    .B(_00697_),
    .Y(_00699_));
 sky130_fd_sc_hd__inv_2 _06873_ (.A(_00695_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2_1 _06874_ (.A(_00699_),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand3b_1 _06875_ (.A_N(_00687_),
    .B(_00698_),
    .C(_00701_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand2_1 _06876_ (.A(_00701_),
    .B(_00698_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(_00703_),
    .B(_00687_),
    .Y(_00704_));
 sky130_fd_sc_hd__nand2_1 _06878_ (.A(_00702_),
    .B(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__inv_2 _06879_ (.A(_00705_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(_00676_),
    .B(_00706_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand3_1 _06881_ (.A(_00705_),
    .B(_00673_),
    .C(_00675_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _06882_ (.A(_00708_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand2_1 _06883_ (.A(_05128_),
    .B(_05131_),
    .Y(_00711_));
 sky130_fd_sc_hd__nor2_1 _06884_ (.A(_05131_),
    .B(_05128_),
    .Y(_00712_));
 sky130_fd_sc_hd__a21oi_2 _06885_ (.A1(_00711_),
    .A2(_05136_),
    .B1(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__inv_2 _06886_ (.A(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _06887_ (.A(_00710_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand3_1 _06888_ (.A(_00708_),
    .B(_00709_),
    .C(_00713_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2_1 _06889_ (.A(_00715_),
    .B(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__nor2_1 _06890_ (.A(_05150_),
    .B(_05172_),
    .Y(_00719_));
 sky130_fd_sc_hd__inv_2 _06891_ (.A(_05203_),
    .Y(_00720_));
 sky130_fd_sc_hd__nor2_1 _06892_ (.A(_00719_),
    .B(_00720_),
    .Y(_00721_));
 sky130_fd_sc_hd__inv_2 _06893_ (.A(_00721_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand2_1 _06894_ (.A(_00717_),
    .B(_00722_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand3_1 _06895_ (.A(_00715_),
    .B(_00716_),
    .C(_00721_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _06896_ (.A(_00723_),
    .B(_00724_),
    .Y(_00725_));
 sky130_fd_sc_hd__inv_2 _06897_ (.A(_00725_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand2_1 _06898_ (.A(_00648_),
    .B(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand3_1 _06899_ (.A(_00645_),
    .B(_00647_),
    .C(_00725_),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_1 _06900_ (.A(_00727_),
    .B(_00728_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _06901_ (.A(_05144_),
    .B(_05022_),
    .Y(_00731_));
 sky130_fd_sc_hd__nor2_1 _06902_ (.A(_05022_),
    .B(_05144_),
    .Y(_00732_));
 sky130_fd_sc_hd__a21oi_2 _06903_ (.A1(_00731_),
    .A2(_05216_),
    .B1(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hd__inv_2 _06904_ (.A(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _06905_ (.A(_00730_),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand3_1 _06906_ (.A(_00733_),
    .B(_00727_),
    .C(_00728_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand2_1 _06907_ (.A(_00735_),
    .B(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__o21a_1 _06908_ (.A1(_05188_),
    .A2(_05185_),
    .B1(_05199_),
    .X(_00738_));
 sky130_fd_sc_hd__or2_1 _06909_ (.A(_05195_),
    .B(_00738_),
    .X(_00739_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(_00738_),
    .B(_05195_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand2_1 _06911_ (.A(_00739_),
    .B(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__o21a_1 _06912_ (.A1(_05205_),
    .A2(_05208_),
    .B1(_05214_),
    .X(_00743_));
 sky130_fd_sc_hd__nor2_1 _06913_ (.A(_00742_),
    .B(_00743_),
    .Y(_00744_));
 sky130_fd_sc_hd__inv_2 _06914_ (.A(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand2_1 _06915_ (.A(_00743_),
    .B(_00742_),
    .Y(_00746_));
 sky130_fd_sc_hd__nand2_1 _06916_ (.A(_00745_),
    .B(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hd__inv_2 _06917_ (.A(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__nand2_1 _06918_ (.A(_00737_),
    .B(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand3_1 _06919_ (.A(_00735_),
    .B(_00736_),
    .C(_00747_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand2_1 _06920_ (.A(_00749_),
    .B(_00750_),
    .Y(_00752_));
 sky130_fd_sc_hd__nor2_1 _06921_ (.A(_05228_),
    .B(_05227_),
    .Y(_00753_));
 sky130_fd_sc_hd__a21oi_2 _06922_ (.A1(_05229_),
    .A2(_05226_),
    .B1(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__inv_2 _06923_ (.A(_00754_),
    .Y(_00755_));
 sky130_fd_sc_hd__nand2_1 _06924_ (.A(_00752_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__nand3_1 _06925_ (.A(_00754_),
    .B(_00749_),
    .C(_00750_),
    .Y(_00757_));
 sky130_fd_sc_hd__nand2_1 _06926_ (.A(_00756_),
    .B(_00757_),
    .Y(_00758_));
 sky130_fd_sc_hd__nand2_1 _06927_ (.A(_00758_),
    .B(_05222_),
    .Y(_00759_));
 sky130_fd_sc_hd__nand3_1 _06928_ (.A(_00756_),
    .B(_00757_),
    .C(_05223_),
    .Y(_00760_));
 sky130_fd_sc_hd__nand3_2 _06929_ (.A(_00516_),
    .B(_00759_),
    .C(_00760_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2_1 _06930_ (.A(_00759_),
    .B(_00760_),
    .Y(_00763_));
 sky130_fd_sc_hd__a21oi_1 _06931_ (.A1(_00514_),
    .A2(_00091_),
    .B1(_00515_),
    .Y(_00764_));
 sky130_fd_sc_hd__nand2_1 _06932_ (.A(_00763_),
    .B(_00764_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand2_1 _06933_ (.A(_00761_),
    .B(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hd__inv_2 _06934_ (.A(_00292_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand2_1 _06935_ (.A(_00766_),
    .B(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand3_1 _06936_ (.A(_00761_),
    .B(_00765_),
    .C(_00292_),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2_2 _06937_ (.A(_00768_),
    .B(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hd__nand3_1 _06938_ (.A(_00491_),
    .B(_00485_),
    .C(_00486_),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_1 _06939_ (.A(_00489_),
    .B(_00480_),
    .Y(_00772_));
 sky130_fd_sc_hd__inv_2 _06940_ (.A(_00493_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand3_1 _06941_ (.A(_00771_),
    .B(_00772_),
    .C(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand2_1 _06942_ (.A(_00494_),
    .B(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand3_1 _06943_ (.A(_00475_),
    .B(_00400_),
    .C(_00403_),
    .Y(_00777_));
 sky130_fd_sc_hd__a21o_1 _06944_ (.A1(_00463_),
    .A2(_00473_),
    .B1(_00474_),
    .X(_00778_));
 sky130_fd_sc_hd__nand2_1 _06945_ (.A(_00404_),
    .B(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hd__nand2_1 _06946_ (.A(_00777_),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(_00780_),
    .B(_00490_),
    .Y(_00781_));
 sky130_fd_sc_hd__nand3_1 _06948_ (.A(_00777_),
    .B(_00779_),
    .C(_00396_),
    .Y(_00782_));
 sky130_fd_sc_hd__nand2_1 _06949_ (.A(_00781_),
    .B(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__a21o_1 _06950_ (.A1(_00451_),
    .A2(_00460_),
    .B1(_00461_),
    .X(_00785_));
 sky130_fd_sc_hd__nand3_1 _06951_ (.A(_00785_),
    .B(_00413_),
    .C(_00414_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand3_1 _06952_ (.A(_00786_),
    .B(_00473_),
    .C(_00463_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand2_1 _06953_ (.A(_00415_),
    .B(_00785_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand3_1 _06954_ (.A(_00462_),
    .B(_00413_),
    .C(_00414_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand3_1 _06955_ (.A(_00788_),
    .B(_00789_),
    .C(_00472_),
    .Y(_00790_));
 sky130_fd_sc_hd__nand2_1 _06956_ (.A(_00787_),
    .B(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__nand3_1 _06957_ (.A(_00450_),
    .B(_00408_),
    .C(_00418_),
    .Y(_00792_));
 sky130_fd_sc_hd__a21o_1 _06958_ (.A1(_00431_),
    .A2(_00435_),
    .B1(_00436_),
    .X(_00793_));
 sky130_fd_sc_hd__nand3_1 _06959_ (.A(_00793_),
    .B(_00427_),
    .C(_00425_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand3_1 _06960_ (.A(_00794_),
    .B(_00438_),
    .C(_00448_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand2_1 _06961_ (.A(_00796_),
    .B(_00794_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _06962_ (.A(_00419_),
    .B(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__nand2_1 _06963_ (.A(_00792_),
    .B(_00798_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_1 _06964_ (.A(_00799_),
    .B(_00460_),
    .Y(_00800_));
 sky130_fd_sc_hd__nand3_2 _06965_ (.A(_00792_),
    .B(_00798_),
    .C(_00459_),
    .Y(_00801_));
 sky130_fd_sc_hd__nand2_1 _06966_ (.A(_00800_),
    .B(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__nand2_1 _06967_ (.A(_00428_),
    .B(_00793_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand3_1 _06968_ (.A(_00437_),
    .B(_00425_),
    .C(_00427_),
    .Y(_00804_));
 sky130_fd_sc_hd__nand3_1 _06969_ (.A(_00803_),
    .B(_00804_),
    .C(_00447_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand2_1 _06970_ (.A(_00796_),
    .B(_00805_),
    .Y(_00807_));
 sky130_fd_sc_hd__inv_2 _06971_ (.A(_00430_),
    .Y(_00808_));
 sky130_fd_sc_hd__nand2_1 _06972_ (.A(_00808_),
    .B(_00429_),
    .Y(_00809_));
 sky130_fd_sc_hd__inv_2 _06973_ (.A(_00429_),
    .Y(_00810_));
 sky130_fd_sc_hd__nand2_1 _06974_ (.A(_00810_),
    .B(_00430_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand3_1 _06975_ (.A(_00809_),
    .B(_00811_),
    .C(_00434_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _06976_ (.A(_00810_),
    .B(_00808_),
    .Y(_00813_));
 sky130_fd_sc_hd__nand3_1 _06977_ (.A(_00813_),
    .B(_00435_),
    .C(_00431_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(_00812_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _06979_ (.A(_00232_),
    .B(_01532_),
    .Y(_00816_));
 sky130_fd_sc_hd__nand2_1 _06980_ (.A(_03105_),
    .B(_00234_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _06981_ (.A(_00816_),
    .B(_00818_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _06982_ (.A(_00433_),
    .B(_01334_),
    .Y(_00820_));
 sky130_fd_sc_hd__inv_2 _06983_ (.A(_00820_),
    .Y(_00821_));
 sky130_fd_sc_hd__nor2_1 _06984_ (.A(_00816_),
    .B(_00818_),
    .Y(_00822_));
 sky130_fd_sc_hd__a21oi_1 _06985_ (.A1(_00819_),
    .A2(_00821_),
    .B1(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__nand2_1 _06986_ (.A(_00815_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_1 _06987_ (.A(_00674_),
    .B(_04128_),
    .Y(_00825_));
 sky130_fd_sc_hd__inv_2 _06988_ (.A(_00825_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _06989_ (.A(_03105_),
    .B(_00641_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_1 _06990_ (.A(_00826_),
    .B(_00827_),
    .Y(_00829_));
 sky130_fd_sc_hd__inv_2 _06991_ (.A(_00827_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_1 _06992_ (.A(_00830_),
    .B(_00825_),
    .Y(_00831_));
 sky130_fd_sc_hd__nand2_1 _06993_ (.A(_05113_),
    .B(_00306_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand3_1 _06994_ (.A(_00829_),
    .B(_00831_),
    .C(_00832_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand2_1 _06995_ (.A(_00830_),
    .B(_00826_),
    .Y(_00834_));
 sky130_fd_sc_hd__inv_2 _06996_ (.A(_00832_),
    .Y(_00835_));
 sky130_fd_sc_hd__nand2_1 _06997_ (.A(_00827_),
    .B(_00825_),
    .Y(_00836_));
 sky130_fd_sc_hd__nand3_1 _06998_ (.A(_00834_),
    .B(_00835_),
    .C(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__nand2_1 _06999_ (.A(_00833_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__inv_2 _07000_ (.A(_00838_),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2_1 _07001_ (.A(_00823_),
    .B(_00815_),
    .Y(_00841_));
 sky130_fd_sc_hd__a21oi_1 _07002_ (.A1(_00824_),
    .A2(_00840_),
    .B1(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__nand2_1 _07003_ (.A(_00807_),
    .B(_00842_),
    .Y(_00843_));
 sky130_fd_sc_hd__nand2_1 _07004_ (.A(_00317_),
    .B(_00313_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(_00314_),
    .B(_00316_),
    .Y(_00845_));
 sky130_fd_sc_hd__nand3_1 _07006_ (.A(_00844_),
    .B(_00845_),
    .C(_00319_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _07007_ (.A(_00846_),
    .B(_00323_),
    .Y(_00847_));
 sky130_fd_sc_hd__nor2_1 _07008_ (.A(_00827_),
    .B(_00825_),
    .Y(_00848_));
 sky130_fd_sc_hd__a21oi_2 _07009_ (.A1(_00836_),
    .A2(_00835_),
    .B1(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__inv_2 _07010_ (.A(_00849_),
    .Y(_00851_));
 sky130_fd_sc_hd__nand2_1 _07011_ (.A(_00847_),
    .B(_00851_),
    .Y(_00852_));
 sky130_fd_sc_hd__nand3_1 _07012_ (.A(_00849_),
    .B(_00846_),
    .C(_00323_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_1 _07013_ (.A(_00852_),
    .B(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__nand2_1 _07014_ (.A(_05278_),
    .B(_05068_),
    .Y(_00855_));
 sky130_fd_sc_hd__inv_2 _07015_ (.A(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand2_1 _07016_ (.A(_00138_),
    .B(_01224_),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _07017_ (.A(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__nand2_1 _07018_ (.A(_00856_),
    .B(_00858_),
    .Y(_00859_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(_00329_),
    .B(_02203_),
    .Y(_00860_));
 sky130_fd_sc_hd__inv_2 _07020_ (.A(_00860_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _07021_ (.A(_00855_),
    .B(_00857_),
    .Y(_00863_));
 sky130_fd_sc_hd__nand3_2 _07022_ (.A(_00859_),
    .B(_00862_),
    .C(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2_1 _07023_ (.A(_00864_),
    .B(_00859_),
    .Y(_00865_));
 sky130_fd_sc_hd__nand2_1 _07024_ (.A(_00854_),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__nand3b_1 _07025_ (.A_N(_00865_),
    .B(_00852_),
    .C(_00853_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2_1 _07026_ (.A(_00866_),
    .B(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__inv_2 _07027_ (.A(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__nor2_1 _07028_ (.A(_00842_),
    .B(_00807_),
    .Y(_00870_));
 sky130_fd_sc_hd__a21oi_2 _07029_ (.A1(_00843_),
    .A2(_00869_),
    .B1(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(_00802_),
    .B(_00871_),
    .Y(_00873_));
 sky130_fd_sc_hd__nand2_1 _07031_ (.A(_00847_),
    .B(_00849_),
    .Y(_00874_));
 sky130_fd_sc_hd__nor2_1 _07032_ (.A(_00849_),
    .B(_00847_),
    .Y(_00875_));
 sky130_fd_sc_hd__a21oi_1 _07033_ (.A1(_00874_),
    .A2(_00865_),
    .B1(_00875_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand3_1 _07034_ (.A(_00347_),
    .B(_00348_),
    .C(_00353_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand3_1 _07035_ (.A(_00876_),
    .B(_00356_),
    .C(_00877_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand2_1 _07036_ (.A(_00356_),
    .B(_00877_),
    .Y(_00879_));
 sky130_fd_sc_hd__a21o_1 _07037_ (.A1(_00874_),
    .A2(_00865_),
    .B1(_00875_),
    .X(_00880_));
 sky130_fd_sc_hd__nand2_1 _07038_ (.A(_00879_),
    .B(_00880_),
    .Y(_00881_));
 sky130_fd_sc_hd__nand2_1 _07039_ (.A(_00878_),
    .B(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__inv_2 _07040_ (.A(_00328_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _07041_ (.A(_00884_),
    .B(_00330_),
    .Y(_00885_));
 sky130_fd_sc_hd__inv_2 _07042_ (.A(_00330_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand2_1 _07043_ (.A(_00886_),
    .B(_00328_),
    .Y(_00887_));
 sky130_fd_sc_hd__nand3_1 _07044_ (.A(_00885_),
    .B(_00887_),
    .C(_00332_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_1 _07045_ (.A(_00884_),
    .B(_00886_),
    .Y(_00889_));
 sky130_fd_sc_hd__nand3_1 _07046_ (.A(_00889_),
    .B(_00334_),
    .C(_00331_),
    .Y(_00890_));
 sky130_fd_sc_hd__nand2_1 _07047_ (.A(_00888_),
    .B(_00890_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_1 _07048_ (.A(_05159_),
    .B(_03039_),
    .Y(_00892_));
 sky130_fd_sc_hd__buf_8 _07049_ (.A(_04814_),
    .X(_00893_));
 sky130_fd_sc_hd__nand2_2 _07050_ (.A(_00893_),
    .B(_05096_),
    .Y(_00895_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(_00892_),
    .B(_00895_),
    .Y(_00896_));
 sky130_fd_sc_hd__nand2_1 _07052_ (.A(_00384_),
    .B(_02687_),
    .Y(_00897_));
 sky130_fd_sc_hd__inv_2 _07053_ (.A(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__nor2_1 _07054_ (.A(_00892_),
    .B(_00895_),
    .Y(_00899_));
 sky130_fd_sc_hd__a21oi_1 _07055_ (.A1(_00896_),
    .A2(_00898_),
    .B1(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hd__inv_2 _07056_ (.A(_00900_),
    .Y(_00901_));
 sky130_fd_sc_hd__nand2_1 _07057_ (.A(_00891_),
    .B(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand3_1 _07058_ (.A(_00900_),
    .B(_00888_),
    .C(_00890_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand2_1 _07059_ (.A(_00902_),
    .B(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_1 _07060_ (.A(_00387_),
    .B(_00389_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand2_1 _07061_ (.A(_00906_),
    .B(_00380_),
    .Y(_00907_));
 sky130_fd_sc_hd__nand2_1 _07062_ (.A(_00907_),
    .B(_00390_),
    .Y(_00908_));
 sky130_fd_sc_hd__inv_2 _07063_ (.A(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand2_1 _07064_ (.A(_00904_),
    .B(_00909_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand3_1 _07065_ (.A(_00901_),
    .B(_00890_),
    .C(_00888_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _07066_ (.A(_00910_),
    .B(_00911_),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_1 _07067_ (.A(_00882_),
    .B(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand3b_1 _07068_ (.A_N(_00912_),
    .B(_00878_),
    .C(_00881_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _07069_ (.A(_00913_),
    .B(_00914_),
    .Y(_00915_));
 sky130_fd_sc_hd__inv_2 _07070_ (.A(_00915_),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2_1 _07071_ (.A(_00871_),
    .B(_00802_),
    .Y(_00918_));
 sky130_fd_sc_hd__a21oi_1 _07072_ (.A1(_00873_),
    .A2(_00917_),
    .B1(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand2_1 _07073_ (.A(_00791_),
    .B(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand2_1 _07074_ (.A(_00879_),
    .B(_00876_),
    .Y(_00921_));
 sky130_fd_sc_hd__nor2_1 _07075_ (.A(_00876_),
    .B(_00879_),
    .Y(_00922_));
 sky130_fd_sc_hd__a21oi_1 _07076_ (.A1(_00921_),
    .A2(_00912_),
    .B1(_00922_),
    .Y(_00923_));
 sky130_fd_sc_hd__inv_2 _07077_ (.A(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand2_1 _07078_ (.A(_00375_),
    .B(_00376_),
    .Y(_00925_));
 sky130_fd_sc_hd__inv_2 _07079_ (.A(_00392_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_1 _07080_ (.A(_00925_),
    .B(_00926_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _07081_ (.A(_00928_),
    .B(_00393_),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _07082_ (.A(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _07083_ (.A(_00924_),
    .B(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _07084_ (.A(_00923_),
    .B(_00929_),
    .Y(_00932_));
 sky130_fd_sc_hd__nand2_1 _07085_ (.A(_00931_),
    .B(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_1 _07086_ (.A(_00194_),
    .B(_04897_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand2_1 _07087_ (.A(_04958_),
    .B(_04645_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand2_1 _07088_ (.A(_04947_),
    .B(_05114_),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _07089_ (.A(_00381_),
    .B(_03248_),
    .Y(_00937_));
 sky130_fd_sc_hd__or2_1 _07090_ (.A(_00936_),
    .B(_00937_),
    .X(_00939_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(_00936_),
    .B(_00937_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand3b_1 _07092_ (.A_N(_00935_),
    .B(_00939_),
    .C(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__and2_1 _07093_ (.A(_00941_),
    .B(_00939_),
    .X(_00942_));
 sky130_fd_sc_hd__nor2_1 _07094_ (.A(_00934_),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__inv_2 _07095_ (.A(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__nand2_1 _07096_ (.A(_00391_),
    .B(_00379_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _07097_ (.A(_00926_),
    .B(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__or2_1 _07098_ (.A(_00944_),
    .B(_00946_),
    .X(_00947_));
 sky130_fd_sc_hd__nand2_1 _07099_ (.A(_00933_),
    .B(_00947_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand3b_1 _07100_ (.A_N(_00947_),
    .B(_00931_),
    .C(_00932_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand2_1 _07101_ (.A(_00948_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__inv_2 _07102_ (.A(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__nor2_1 _07103_ (.A(_00919_),
    .B(_00791_),
    .Y(_00953_));
 sky130_fd_sc_hd__a21oi_2 _07104_ (.A1(_00920_),
    .A2(_00952_),
    .B1(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__nand2_1 _07105_ (.A(_00783_),
    .B(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_2 _07106_ (.A(_00950_),
    .B(_00931_),
    .Y(_00956_));
 sky130_fd_sc_hd__nor2_1 _07107_ (.A(_00954_),
    .B(_00783_),
    .Y(_00957_));
 sky130_fd_sc_hd__a21oi_2 _07108_ (.A1(_00955_),
    .A2(_00956_),
    .B1(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__inv_2 _07109_ (.A(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(_00776_),
    .B(_00959_),
    .Y(_00961_));
 sky130_fd_sc_hd__nand3_1 _07111_ (.A(_00958_),
    .B(_00494_),
    .C(_00775_),
    .Y(_00962_));
 sky130_fd_sc_hd__nand2_1 _07112_ (.A(_00961_),
    .B(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand3_1 _07113_ (.A(_00919_),
    .B(_00787_),
    .C(_00790_),
    .Y(_00964_));
 sky130_fd_sc_hd__a21o_1 _07114_ (.A1(_00873_),
    .A2(_00917_),
    .B1(_00918_),
    .X(_00965_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(_00791_),
    .B(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__nand2_1 _07116_ (.A(_00964_),
    .B(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand2_1 _07117_ (.A(_00967_),
    .B(_00952_),
    .Y(_00968_));
 sky130_fd_sc_hd__nand3_1 _07118_ (.A(_00964_),
    .B(_00966_),
    .C(_00951_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_1 _07119_ (.A(_00968_),
    .B(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__a21o_1 _07120_ (.A1(_00843_),
    .A2(_00869_),
    .B1(_00870_),
    .X(_00972_));
 sky130_fd_sc_hd__nand3_1 _07121_ (.A(_00972_),
    .B(_00800_),
    .C(_00801_),
    .Y(_00973_));
 sky130_fd_sc_hd__nand3_1 _07122_ (.A(_00973_),
    .B(_00917_),
    .C(_00873_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand2_1 _07123_ (.A(_00802_),
    .B(_00972_),
    .Y(_00975_));
 sky130_fd_sc_hd__nand3_1 _07124_ (.A(_00871_),
    .B(_00800_),
    .C(_00801_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand3_1 _07125_ (.A(_00975_),
    .B(_00976_),
    .C(_00915_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_1 _07126_ (.A(_00974_),
    .B(_00977_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand3_1 _07127_ (.A(_00842_),
    .B(_00796_),
    .C(_00805_),
    .Y(_00979_));
 sky130_fd_sc_hd__a21o_1 _07128_ (.A1(_00819_),
    .A2(_00821_),
    .B1(_00822_),
    .X(_00980_));
 sky130_fd_sc_hd__nand3_1 _07129_ (.A(_00980_),
    .B(_00814_),
    .C(_00812_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand3_1 _07130_ (.A(_00981_),
    .B(_00824_),
    .C(_00840_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_1 _07131_ (.A(_00983_),
    .B(_00981_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _07132_ (.A(_00807_),
    .B(_00984_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _07133_ (.A(_00979_),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _07134_ (.A(_00986_),
    .B(_00869_),
    .Y(_00987_));
 sky130_fd_sc_hd__nand3_1 _07135_ (.A(_00979_),
    .B(_00985_),
    .C(_00868_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _07136_ (.A(_00987_),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _07137_ (.A(_00815_),
    .B(_00980_),
    .Y(_00990_));
 sky130_fd_sc_hd__nand3_1 _07138_ (.A(_00823_),
    .B(_00812_),
    .C(_00814_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand3_1 _07139_ (.A(_00990_),
    .B(_00991_),
    .C(_00838_),
    .Y(_00992_));
 sky130_fd_sc_hd__nand2_1 _07140_ (.A(_00983_),
    .B(_00992_),
    .Y(_00994_));
 sky130_fd_sc_hd__inv_2 _07141_ (.A(_00818_),
    .Y(_00995_));
 sky130_fd_sc_hd__nand2_1 _07142_ (.A(_00995_),
    .B(_00816_),
    .Y(_00996_));
 sky130_fd_sc_hd__inv_2 _07143_ (.A(_00816_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_1 _07144_ (.A(_00997_),
    .B(_00818_),
    .Y(_00998_));
 sky130_fd_sc_hd__nand3_1 _07145_ (.A(_00996_),
    .B(_00998_),
    .C(_00820_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _07146_ (.A(_00997_),
    .B(_00995_),
    .Y(_01000_));
 sky130_fd_sc_hd__nand3_1 _07147_ (.A(_01000_),
    .B(_00821_),
    .C(_00819_),
    .Y(_01001_));
 sky130_fd_sc_hd__nand2_1 _07148_ (.A(_00999_),
    .B(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__nand2_2 _07149_ (.A(_03105_),
    .B(_00232_),
    .Y(_01003_));
 sky130_fd_sc_hd__nand2_1 _07150_ (.A(_05113_),
    .B(_00234_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _07151_ (.A(_01003_),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand2_1 _07152_ (.A(_00410_),
    .B(_01532_),
    .Y(_01007_));
 sky130_fd_sc_hd__inv_2 _07153_ (.A(_01007_),
    .Y(_01008_));
 sky130_fd_sc_hd__nor2_1 _07154_ (.A(_01003_),
    .B(_01005_),
    .Y(_01009_));
 sky130_fd_sc_hd__a21oi_2 _07155_ (.A1(_01006_),
    .A2(_01008_),
    .B1(_01009_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_1 _07156_ (.A(_01002_),
    .B(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(_05113_),
    .B(_00301_),
    .Y(_01012_));
 sky130_fd_sc_hd__inv_2 _07158_ (.A(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _07159_ (.A(_00303_),
    .B(_02214_),
    .Y(_01014_));
 sky130_fd_sc_hd__inv_2 _07160_ (.A(_01014_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _07161_ (.A(_01013_),
    .B(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _07162_ (.A(_01012_),
    .B(_01014_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _07163_ (.A(_01017_),
    .B(_01018_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2_1 _07164_ (.A(_05278_),
    .B(_00306_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_1 _07165_ (.A(_01019_),
    .B(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hd__inv_2 _07166_ (.A(_01020_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand3_1 _07167_ (.A(_01017_),
    .B(_01022_),
    .C(_01018_),
    .Y(_01023_));
 sky130_fd_sc_hd__nand2_1 _07168_ (.A(_01021_),
    .B(_01023_),
    .Y(_01024_));
 sky130_fd_sc_hd__inv_2 _07169_ (.A(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__nor2_1 _07170_ (.A(_01010_),
    .B(_01002_),
    .Y(_01027_));
 sky130_fd_sc_hd__a21oi_1 _07171_ (.A1(_01011_),
    .A2(_01025_),
    .B1(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand2_1 _07172_ (.A(_00994_),
    .B(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _07173_ (.A(_00138_),
    .B(_05068_),
    .Y(_01030_));
 sky130_fd_sc_hd__inv_2 _07174_ (.A(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _07175_ (.A(_00329_),
    .B(_00315_),
    .Y(_01032_));
 sky130_fd_sc_hd__inv_2 _07176_ (.A(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__nand2_1 _07177_ (.A(_01031_),
    .B(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__nand2_1 _07178_ (.A(_05159_),
    .B(_02203_),
    .Y(_01035_));
 sky130_fd_sc_hd__inv_2 _07179_ (.A(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__nand2_1 _07180_ (.A(_01030_),
    .B(_01032_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand3_1 _07181_ (.A(_01034_),
    .B(_01036_),
    .C(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__nand2_1 _07182_ (.A(_01039_),
    .B(_01034_),
    .Y(_01040_));
 sky130_fd_sc_hd__nand2_1 _07183_ (.A(_00858_),
    .B(_00855_),
    .Y(_01041_));
 sky130_fd_sc_hd__nand2_1 _07184_ (.A(_00856_),
    .B(_00857_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand3_1 _07185_ (.A(_01041_),
    .B(_01042_),
    .C(_00860_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand2_1 _07186_ (.A(_01043_),
    .B(_00864_),
    .Y(_01044_));
 sky130_fd_sc_hd__nor2_1 _07187_ (.A(_01012_),
    .B(_01014_),
    .Y(_01045_));
 sky130_fd_sc_hd__a21o_1 _07188_ (.A1(_01018_),
    .A2(_01022_),
    .B1(_01045_),
    .X(_01046_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(_01044_),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__a21oi_2 _07190_ (.A1(_01018_),
    .A2(_01022_),
    .B1(_01045_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand3_1 _07191_ (.A(_01049_),
    .B(_01043_),
    .C(_00864_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand3b_1 _07192_ (.A_N(_01040_),
    .B(_01047_),
    .C(_01050_),
    .Y(_01051_));
 sky130_fd_sc_hd__nand3_1 _07193_ (.A(_01046_),
    .B(_00864_),
    .C(_01043_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand2_1 _07194_ (.A(_01044_),
    .B(_01049_),
    .Y(_01053_));
 sky130_fd_sc_hd__nand3_1 _07195_ (.A(_01052_),
    .B(_01053_),
    .C(_01040_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _07196_ (.A(_01051_),
    .B(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__inv_2 _07197_ (.A(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__nor2_1 _07198_ (.A(_01028_),
    .B(_00994_),
    .Y(_01057_));
 sky130_fd_sc_hd__a21oi_2 _07199_ (.A1(_01029_),
    .A2(_01056_),
    .B1(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__nand2_1 _07200_ (.A(_00989_),
    .B(_01058_),
    .Y(_01060_));
 sky130_fd_sc_hd__nor2_1 _07201_ (.A(_01049_),
    .B(_01044_),
    .Y(_01061_));
 sky130_fd_sc_hd__a21oi_1 _07202_ (.A1(_01053_),
    .A2(_01040_),
    .B1(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__nand3_1 _07203_ (.A(_00902_),
    .B(_00903_),
    .C(_00908_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand3_1 _07204_ (.A(_01062_),
    .B(_00910_),
    .C(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _07205_ (.A(_00910_),
    .B(_01063_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand2_1 _07206_ (.A(_01054_),
    .B(_01052_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_1 _07207_ (.A(_01065_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _07208_ (.A(_01064_),
    .B(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__inv_2 _07209_ (.A(_00895_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_1 _07210_ (.A(_01069_),
    .B(_00892_),
    .Y(_01071_));
 sky130_fd_sc_hd__inv_2 _07211_ (.A(_00892_),
    .Y(_01072_));
 sky130_fd_sc_hd__nand2_1 _07212_ (.A(_01072_),
    .B(_00895_),
    .Y(_01073_));
 sky130_fd_sc_hd__nand3_1 _07213_ (.A(_01071_),
    .B(_01073_),
    .C(_00897_),
    .Y(_01074_));
 sky130_fd_sc_hd__nand2_1 _07214_ (.A(_01072_),
    .B(_01069_),
    .Y(_01075_));
 sky130_fd_sc_hd__nand3_1 _07215_ (.A(_01075_),
    .B(_00898_),
    .C(_00896_),
    .Y(_01076_));
 sky130_fd_sc_hd__nand2_1 _07216_ (.A(_01074_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand2_1 _07217_ (.A(_00384_),
    .B(_05096_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand2_1 _07218_ (.A(_00893_),
    .B(_03039_),
    .Y(_01079_));
 sky130_fd_sc_hd__nand2_1 _07219_ (.A(_01078_),
    .B(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_1 _07220_ (.A(_00381_),
    .B(_02687_),
    .Y(_01082_));
 sky130_fd_sc_hd__inv_2 _07221_ (.A(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__nor2_1 _07222_ (.A(_01078_),
    .B(_01079_),
    .Y(_01084_));
 sky130_fd_sc_hd__a21oi_1 _07223_ (.A1(_01080_),
    .A2(_01083_),
    .B1(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__inv_2 _07224_ (.A(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__nand2_1 _07225_ (.A(_01077_),
    .B(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__nand3_1 _07226_ (.A(_01085_),
    .B(_01074_),
    .C(_01076_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2_1 _07227_ (.A(_01087_),
    .B(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _07228_ (.A(_00939_),
    .B(_00940_),
    .Y(_01090_));
 sky130_fd_sc_hd__nand2_1 _07229_ (.A(_01090_),
    .B(_00935_),
    .Y(_01091_));
 sky130_fd_sc_hd__nand2_1 _07230_ (.A(_01091_),
    .B(_00941_),
    .Y(_01093_));
 sky130_fd_sc_hd__inv_2 _07231_ (.A(_01093_),
    .Y(_01094_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(_01089_),
    .B(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__or2_1 _07233_ (.A(_01085_),
    .B(_01077_),
    .X(_01096_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(_01095_),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_1 _07235_ (.A(_01068_),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand3b_1 _07236_ (.A_N(_01097_),
    .B(_01064_),
    .C(_01067_),
    .Y(_01099_));
 sky130_fd_sc_hd__nand2_1 _07237_ (.A(_01098_),
    .B(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__inv_2 _07238_ (.A(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hd__nor2_1 _07239_ (.A(_01058_),
    .B(_00989_),
    .Y(_01102_));
 sky130_fd_sc_hd__a21oi_1 _07240_ (.A1(_01060_),
    .A2(_01101_),
    .B1(_01102_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _07241_ (.A(_00978_),
    .B(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(_00946_),
    .B(_00944_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand2_1 _07243_ (.A(_00947_),
    .B(_01106_),
    .Y(_01107_));
 sky130_fd_sc_hd__o21a_1 _07244_ (.A1(_01065_),
    .A2(_01062_),
    .B1(_01098_),
    .X(_01108_));
 sky130_fd_sc_hd__nor2_2 _07245_ (.A(_01107_),
    .B(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_1 _07246_ (.A(_01108_),
    .B(_01107_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2b_1 _07247_ (.A(_01109_),
    .B_N(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_1 _07248_ (.A(_01104_),
    .B(_00978_),
    .Y(_01112_));
 sky130_fd_sc_hd__a21oi_2 _07249_ (.A1(_01105_),
    .A2(_01111_),
    .B1(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _07250_ (.A(_00970_),
    .B(_01113_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _07251_ (.A(_01113_),
    .B(_00970_),
    .Y(_01116_));
 sky130_fd_sc_hd__a21oi_1 _07252_ (.A1(_01115_),
    .A2(_01109_),
    .B1(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__inv_2 _07253_ (.A(_00954_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand2_1 _07254_ (.A(_00783_),
    .B(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand3_1 _07255_ (.A(_00954_),
    .B(_00781_),
    .C(_00782_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _07256_ (.A(_01119_),
    .B(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_1 _07257_ (.A(_01121_),
    .B(_00956_),
    .Y(_01122_));
 sky130_fd_sc_hd__inv_2 _07258_ (.A(_00956_),
    .Y(_01123_));
 sky130_fd_sc_hd__nand3_1 _07259_ (.A(_01119_),
    .B(_01120_),
    .C(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(_01122_),
    .B(_01124_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_1 _07261_ (.A(_01117_),
    .B(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(_00963_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__nand2_1 _07263_ (.A(_00501_),
    .B(_00502_),
    .Y(_01129_));
 sky130_fd_sc_hd__inv_2 _07264_ (.A(_00495_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _07265_ (.A(_01129_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand2_1 _07266_ (.A(_01131_),
    .B(_00503_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_1 _07267_ (.A(_00958_),
    .B(_00776_),
    .Y(_01133_));
 sky130_fd_sc_hd__inv_2 _07268_ (.A(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hd__nand2_1 _07269_ (.A(_01132_),
    .B(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand3_2 _07270_ (.A(_01131_),
    .B(_00503_),
    .C(_01133_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand3b_2 _07271_ (.A_N(_01128_),
    .B(_01135_),
    .C(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand2_1 _07272_ (.A(_00289_),
    .B(_00506_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _07273_ (.A(_01139_),
    .B(_00504_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand3_1 _07274_ (.A(_00289_),
    .B(_00506_),
    .C(_00503_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand3_1 _07275_ (.A(_01140_),
    .B(_01141_),
    .C(_01137_),
    .Y(_01142_));
 sky130_fd_sc_hd__inv_2 _07276_ (.A(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(_01140_),
    .B(_01141_),
    .Y(_01144_));
 sky130_fd_sc_hd__inv_2 _07278_ (.A(_01137_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand2_1 _07279_ (.A(_01144_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__o21ai_1 _07280_ (.A1(_01138_),
    .A2(_01143_),
    .B1(_01146_),
    .Y(_01148_));
 sky130_fd_sc_hd__nand3_1 _07281_ (.A(_00513_),
    .B(_00770_),
    .C(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(_00766_),
    .B(_00292_),
    .Y(_01150_));
 sky130_fd_sc_hd__inv_2 _07283_ (.A(_00511_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _07284_ (.A(_00292_),
    .B(_00766_),
    .Y(_01152_));
 sky130_fd_sc_hd__a21oi_1 _07285_ (.A1(_01150_),
    .A2(_01151_),
    .B1(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__nand2_1 _07286_ (.A(_01149_),
    .B(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand3_1 _07287_ (.A(_01104_),
    .B(_00974_),
    .C(_00977_),
    .Y(_01155_));
 sky130_fd_sc_hd__a21o_1 _07288_ (.A1(_01060_),
    .A2(_01101_),
    .B1(_01102_),
    .X(_01156_));
 sky130_fd_sc_hd__nand2_1 _07289_ (.A(_00978_),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand2_1 _07290_ (.A(_01155_),
    .B(_01157_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _07291_ (.A(_01159_),
    .B(_01111_),
    .Y(_01160_));
 sky130_fd_sc_hd__inv_2 _07292_ (.A(_01109_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2_1 _07293_ (.A(_01161_),
    .B(_01110_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand3_1 _07294_ (.A(_01155_),
    .B(_01157_),
    .C(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _07295_ (.A(_01160_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__inv_2 _07296_ (.A(_01058_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand2_1 _07297_ (.A(_00989_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand3_1 _07298_ (.A(_01058_),
    .B(_00987_),
    .C(_00988_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand2_1 _07299_ (.A(_01166_),
    .B(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hd__nand2_1 _07300_ (.A(_01168_),
    .B(_01101_),
    .Y(_01170_));
 sky130_fd_sc_hd__nand3_1 _07301_ (.A(_01166_),
    .B(_01167_),
    .C(_01100_),
    .Y(_01171_));
 sky130_fd_sc_hd__nand2_1 _07302_ (.A(_01170_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand3_1 _07303_ (.A(_01028_),
    .B(_00983_),
    .C(_00992_),
    .Y(_01173_));
 sky130_fd_sc_hd__a21o_1 _07304_ (.A1(_01011_),
    .A2(_01025_),
    .B1(_01027_),
    .X(_01174_));
 sky130_fd_sc_hd__nand2_1 _07305_ (.A(_01174_),
    .B(_00994_),
    .Y(_01175_));
 sky130_fd_sc_hd__nand2_1 _07306_ (.A(_01173_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_1 _07307_ (.A(_01176_),
    .B(_01056_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand3_1 _07308_ (.A(_01173_),
    .B(_01175_),
    .C(_01055_),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_1 _07309_ (.A(_01177_),
    .B(_01178_),
    .Y(_01179_));
 sky130_fd_sc_hd__inv_2 _07310_ (.A(_01010_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand2_1 _07311_ (.A(_01002_),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__nand3_1 _07312_ (.A(_01010_),
    .B(_00999_),
    .C(_01001_),
    .Y(_01183_));
 sky130_fd_sc_hd__nand2_1 _07313_ (.A(_01182_),
    .B(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _07314_ (.A(_01184_),
    .B(_01025_),
    .Y(_01185_));
 sky130_fd_sc_hd__nand3_1 _07315_ (.A(_01182_),
    .B(_01183_),
    .C(_01024_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _07316_ (.A(_01185_),
    .B(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__inv_2 _07317_ (.A(_01005_),
    .Y(_01188_));
 sky130_fd_sc_hd__nand2_1 _07318_ (.A(_01188_),
    .B(_01003_),
    .Y(_01189_));
 sky130_fd_sc_hd__inv_2 _07319_ (.A(_01003_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _07320_ (.A(_01190_),
    .B(_01005_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand3_1 _07321_ (.A(_01189_),
    .B(_01192_),
    .C(_01007_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_1 _07322_ (.A(_01190_),
    .B(_01188_),
    .Y(_01194_));
 sky130_fd_sc_hd__nand3_1 _07323_ (.A(_01194_),
    .B(_01008_),
    .C(_01006_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _07324_ (.A(_01193_),
    .B(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_1 _07325_ (.A(_02511_),
    .B(net55),
    .Y(_01197_));
 sky130_fd_sc_hd__nand2_1 _07326_ (.A(_02555_),
    .B(net58),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_1 _07327_ (.A(_01197_),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _07328_ (.A(_02489_),
    .B(_00410_),
    .Y(_01200_));
 sky130_fd_sc_hd__inv_2 _07329_ (.A(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _07330_ (.A(_01197_),
    .B(_01198_),
    .Y(_01203_));
 sky130_fd_sc_hd__a21oi_4 _07331_ (.A1(_01199_),
    .A2(_01201_),
    .B1(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _07332_ (.A(_01196_),
    .B(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _07333_ (.A(_05278_),
    .B(_00301_),
    .Y(_01206_));
 sky130_fd_sc_hd__inv_2 _07334_ (.A(_01206_),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _07335_ (.A(_00303_),
    .B(_01334_),
    .Y(_01208_));
 sky130_fd_sc_hd__inv_2 _07336_ (.A(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_1 _07337_ (.A(_01207_),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_1 _07338_ (.A(_01206_),
    .B(_01208_),
    .Y(_01211_));
 sky130_fd_sc_hd__nand2_1 _07339_ (.A(_01210_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__nand2_1 _07340_ (.A(_00138_),
    .B(_00306_),
    .Y(_01214_));
 sky130_fd_sc_hd__nand2_1 _07341_ (.A(_01212_),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__inv_2 _07342_ (.A(_01214_),
    .Y(_01216_));
 sky130_fd_sc_hd__nand3_1 _07343_ (.A(_01210_),
    .B(_01216_),
    .C(_01211_),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_1 _07344_ (.A(_01215_),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__inv_2 _07345_ (.A(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_1 _07346_ (.A(_01204_),
    .B(_01196_),
    .Y(_01220_));
 sky130_fd_sc_hd__a21oi_1 _07347_ (.A1(_01205_),
    .A2(_01219_),
    .B1(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_1 _07348_ (.A(_01187_),
    .B(_01221_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand2_1 _07349_ (.A(_01033_),
    .B(_01030_),
    .Y(_01223_));
 sky130_fd_sc_hd__nand2_1 _07350_ (.A(_01031_),
    .B(_01032_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand3_1 _07351_ (.A(_01223_),
    .B(_01225_),
    .C(_01035_),
    .Y(_01226_));
 sky130_fd_sc_hd__nand2_1 _07352_ (.A(_01226_),
    .B(_01039_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor2_1 _07353_ (.A(_01206_),
    .B(_01208_),
    .Y(_01228_));
 sky130_fd_sc_hd__a21oi_2 _07354_ (.A1(_01211_),
    .A2(_01216_),
    .B1(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__inv_2 _07355_ (.A(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(_01227_),
    .B(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand3_1 _07357_ (.A(_01229_),
    .B(_01226_),
    .C(_01039_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_1 _07358_ (.A(_01231_),
    .B(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _07359_ (.A(_00893_),
    .B(_02203_),
    .Y(_01234_));
 sky130_fd_sc_hd__nand2_1 _07360_ (.A(_05159_),
    .B(_00315_),
    .Y(_01236_));
 sky130_fd_sc_hd__inv_2 _07361_ (.A(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_1 _07362_ (.A(_00329_),
    .B(_05068_),
    .Y(_01238_));
 sky130_fd_sc_hd__inv_2 _07363_ (.A(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__nand2_1 _07364_ (.A(_01237_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__nand2_1 _07365_ (.A(_01236_),
    .B(_01238_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand3b_2 _07366_ (.A_N(_01234_),
    .B(_01240_),
    .C(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand2_1 _07367_ (.A(_01242_),
    .B(_01240_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(_01233_),
    .B(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand3b_1 _07369_ (.A_N(_01243_),
    .B(_01231_),
    .C(_01232_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand2_1 _07370_ (.A(_01244_),
    .B(_01245_),
    .Y(_01247_));
 sky130_fd_sc_hd__inv_2 _07371_ (.A(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _07372_ (.A(_01221_),
    .B(_01187_),
    .Y(_01249_));
 sky130_fd_sc_hd__a21oi_2 _07373_ (.A1(_01222_),
    .A2(_01248_),
    .B1(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__nand2_1 _07374_ (.A(_01179_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__inv_2 _07375_ (.A(_01080_),
    .Y(_01252_));
 sky130_fd_sc_hd__o21ai_2 _07376_ (.A1(_01084_),
    .A2(_01252_),
    .B1(_01082_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand3b_1 _07377_ (.A_N(_01084_),
    .B(_01083_),
    .C(_01080_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand2_1 _07378_ (.A(_01253_),
    .B(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2_1 _07379_ (.A(_00381_),
    .B(_05096_),
    .Y(_01256_));
 sky130_fd_sc_hd__nand2_1 _07380_ (.A(_00384_),
    .B(_03039_),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _07381_ (.A(_01256_),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand2_1 _07382_ (.A(_05310_),
    .B(_02687_),
    .Y(_01260_));
 sky130_fd_sc_hd__inv_2 _07383_ (.A(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_1 _07384_ (.A(_01256_),
    .B(_01258_),
    .Y(_01262_));
 sky130_fd_sc_hd__a21oi_2 _07385_ (.A1(_01259_),
    .A2(_01261_),
    .B1(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__nand2_1 _07386_ (.A(_01255_),
    .B(_01263_),
    .Y(_01264_));
 sky130_fd_sc_hd__inv_2 _07387_ (.A(_01263_),
    .Y(_01265_));
 sky130_fd_sc_hd__nand3_1 _07388_ (.A(_01253_),
    .B(_01254_),
    .C(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__clkinv_4 _07389_ (.A(net36),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_1 _07390_ (.A(_04958_),
    .B(_05114_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor3_1 _07391_ (.A(_00187_),
    .B(_01267_),
    .C(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__inv_2 _07392_ (.A(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__o21ai_1 _07393_ (.A1(_00187_),
    .A2(_01267_),
    .B1(_01269_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _07394_ (.A(_01271_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__inv_2 _07395_ (.A(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand3_1 _07396_ (.A(_01264_),
    .B(_01266_),
    .C(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(_01275_),
    .B(_01266_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand3_1 _07398_ (.A(_01087_),
    .B(_01093_),
    .C(_01088_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_1 _07399_ (.A(_01095_),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2_1 _07400_ (.A(_01227_),
    .B(_01229_),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_1 _07401_ (.A(_01229_),
    .B(_01227_),
    .Y(_01281_));
 sky130_fd_sc_hd__a21o_1 _07402_ (.A1(_01280_),
    .A2(_01243_),
    .B1(_01281_),
    .X(_01282_));
 sky130_fd_sc_hd__nand2_1 _07403_ (.A(_01278_),
    .B(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__a21oi_1 _07404_ (.A1(_01280_),
    .A2(_01243_),
    .B1(_01281_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand3_1 _07405_ (.A(_01284_),
    .B(_01095_),
    .C(_01277_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand3b_1 _07406_ (.A_N(_01276_),
    .B(_01283_),
    .C(_01285_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _07407_ (.A(_01285_),
    .B(_01283_),
    .Y(_01287_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(_01287_),
    .B(_01276_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_1 _07409_ (.A(_01286_),
    .B(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__inv_2 _07410_ (.A(_01289_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_1 _07411_ (.A(_01250_),
    .B(_01179_),
    .Y(_01292_));
 sky130_fd_sc_hd__a21oi_1 _07412_ (.A1(_01251_),
    .A2(_01291_),
    .B1(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_1 _07413_ (.A(_01172_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(_00942_),
    .B(_00934_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _07415_ (.A(_00944_),
    .B(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__o21a_1 _07416_ (.A1(_01278_),
    .A2(_01284_),
    .B1(_01288_),
    .X(_01297_));
 sky130_fd_sc_hd__nor2_2 _07417_ (.A(_01296_),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _07418_ (.A(_01297_),
    .B(_01296_),
    .Y(_01299_));
 sky130_fd_sc_hd__nor2b_1 _07419_ (.A(_01298_),
    .B_N(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _07420_ (.A(_01293_),
    .B(_01172_),
    .Y(_01302_));
 sky130_fd_sc_hd__a21oi_2 _07421_ (.A1(_01294_),
    .A2(_01300_),
    .B1(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__nand2_1 _07422_ (.A(_01164_),
    .B(_01303_),
    .Y(_01304_));
 sky130_fd_sc_hd__nor2_1 _07423_ (.A(_01303_),
    .B(_01164_),
    .Y(_01305_));
 sky130_fd_sc_hd__a21o_1 _07424_ (.A1(_01304_),
    .A2(_01298_),
    .B1(_01305_),
    .X(_01306_));
 sky130_fd_sc_hd__inv_2 _07425_ (.A(_01113_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(_00970_),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand3_1 _07427_ (.A(_01113_),
    .B(_00968_),
    .C(_00969_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _07428_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand2_1 _07429_ (.A(_01310_),
    .B(_01109_),
    .Y(_01311_));
 sky130_fd_sc_hd__nand3_1 _07430_ (.A(_01308_),
    .B(_01309_),
    .C(_01161_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand3_2 _07431_ (.A(_01306_),
    .B(_01311_),
    .C(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__nand3_1 _07432_ (.A(_01293_),
    .B(_01170_),
    .C(_01171_),
    .Y(_01315_));
 sky130_fd_sc_hd__a21o_1 _07433_ (.A1(_01222_),
    .A2(_01248_),
    .B1(_01249_),
    .X(_01316_));
 sky130_fd_sc_hd__nand3_1 _07434_ (.A(_01316_),
    .B(_01177_),
    .C(_01178_),
    .Y(_01317_));
 sky130_fd_sc_hd__nand3_1 _07435_ (.A(_01317_),
    .B(_01291_),
    .C(_01251_),
    .Y(_01318_));
 sky130_fd_sc_hd__nand2_1 _07436_ (.A(_01318_),
    .B(_01317_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand2_1 _07437_ (.A(_01319_),
    .B(_01172_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand2_1 _07438_ (.A(_01315_),
    .B(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_1 _07439_ (.A(_01321_),
    .B(_01300_),
    .Y(_01322_));
 sky130_fd_sc_hd__inv_2 _07440_ (.A(_01298_),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2_1 _07441_ (.A(_01324_),
    .B(_01299_),
    .Y(_01325_));
 sky130_fd_sc_hd__nand3_1 _07442_ (.A(_01315_),
    .B(_01320_),
    .C(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_1 _07443_ (.A(_01322_),
    .B(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__nand2_1 _07444_ (.A(_01179_),
    .B(_01316_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand3_1 _07445_ (.A(_01250_),
    .B(_01177_),
    .C(_01178_),
    .Y(_01329_));
 sky130_fd_sc_hd__nand3_1 _07446_ (.A(_01328_),
    .B(_01329_),
    .C(_01289_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _07447_ (.A(_01318_),
    .B(_01330_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _07448_ (.A(_01255_),
    .B(_01265_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand3_1 _07449_ (.A(_01253_),
    .B(_01254_),
    .C(_01263_),
    .Y(_01333_));
 sky130_fd_sc_hd__nand3_1 _07450_ (.A(_01332_),
    .B(_01333_),
    .C(_01273_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(_01275_),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__nand2_1 _07452_ (.A(_01240_),
    .B(_01241_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _07453_ (.A(_01337_),
    .B(_01234_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2_1 _07454_ (.A(_01338_),
    .B(_01242_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand2_1 _07455_ (.A(_02797_),
    .B(_00641_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _07456_ (.A(_00674_),
    .B(_01521_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand2_1 _07457_ (.A(_01340_),
    .B(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__nand2_1 _07458_ (.A(_02874_),
    .B(_00751_),
    .Y(_01343_));
 sky130_fd_sc_hd__inv_2 _07459_ (.A(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _07460_ (.A(_01340_),
    .B(_01341_),
    .Y(_01346_));
 sky130_fd_sc_hd__a21oi_2 _07461_ (.A1(_01342_),
    .A2(_01344_),
    .B1(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_1 _07462_ (.A(_01339_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__nand2_1 _07463_ (.A(_04814_),
    .B(_01224_),
    .Y(_01349_));
 sky130_fd_sc_hd__inv_2 _07464_ (.A(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(_04634_),
    .B(_01257_),
    .Y(_01351_));
 sky130_fd_sc_hd__inv_2 _07466_ (.A(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_1 _07467_ (.A(_01350_),
    .B(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_1 _07468_ (.A(_04880_),
    .B(_01323_),
    .Y(_01354_));
 sky130_fd_sc_hd__inv_2 _07469_ (.A(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__nand2_1 _07470_ (.A(_01349_),
    .B(_01351_),
    .Y(_01357_));
 sky130_fd_sc_hd__nand3_1 _07471_ (.A(_01353_),
    .B(_01355_),
    .C(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__nand2_2 _07472_ (.A(_01358_),
    .B(_01353_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _07473_ (.A(_01347_),
    .B(_01339_),
    .Y(_01360_));
 sky130_fd_sc_hd__a21oi_2 _07474_ (.A1(_01348_),
    .A2(_01359_),
    .B1(_01360_),
    .Y(_01361_));
 sky130_fd_sc_hd__inv_2 _07475_ (.A(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__nand2_1 _07476_ (.A(_01336_),
    .B(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__nand3_1 _07477_ (.A(_01361_),
    .B(_01275_),
    .C(_01335_),
    .Y(_01364_));
 sky130_fd_sc_hd__nand2_1 _07478_ (.A(_01363_),
    .B(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_1 _07479_ (.A(_00194_),
    .B(_03248_),
    .Y(_01366_));
 sky130_fd_sc_hd__inv_2 _07480_ (.A(_01259_),
    .Y(_01368_));
 sky130_fd_sc_hd__o21ai_1 _07481_ (.A1(_01262_),
    .A2(_01368_),
    .B1(_01260_),
    .Y(_01369_));
 sky130_fd_sc_hd__nand3b_1 _07482_ (.A_N(_01262_),
    .B(_01261_),
    .C(_01259_),
    .Y(_01370_));
 sky130_fd_sc_hd__nand2_1 _07483_ (.A(_01369_),
    .B(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__nand2_1 _07484_ (.A(net12),
    .B(_02522_),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_1 _07485_ (.A(_04895_),
    .B(net64),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _07486_ (.A(_01372_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _07487_ (.A(_04958_),
    .B(_02687_),
    .Y(_01375_));
 sky130_fd_sc_hd__inv_2 _07488_ (.A(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _07489_ (.A(_01372_),
    .B(_01373_),
    .Y(_01377_));
 sky130_fd_sc_hd__a21oi_1 _07490_ (.A1(_01374_),
    .A2(_01376_),
    .B1(_01377_),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_1 _07491_ (.A(_01371_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__inv_2 _07492_ (.A(_01379_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand3_1 _07493_ (.A(_01369_),
    .B(_01370_),
    .C(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand3b_2 _07494_ (.A_N(_01366_),
    .B(_01380_),
    .C(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__nand2_1 _07495_ (.A(_01383_),
    .B(_01382_),
    .Y(_01384_));
 sky130_fd_sc_hd__nand2_1 _07496_ (.A(_01365_),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand3b_1 _07497_ (.A_N(_01384_),
    .B(_01363_),
    .C(_01364_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(_01385_),
    .B(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__inv_2 _07499_ (.A(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__nand3_1 _07500_ (.A(_01221_),
    .B(_01185_),
    .C(_01186_),
    .Y(_01390_));
 sky130_fd_sc_hd__a21o_1 _07501_ (.A1(_01205_),
    .A2(_01219_),
    .B1(_01220_),
    .X(_01391_));
 sky130_fd_sc_hd__nand2_1 _07502_ (.A(_01391_),
    .B(_01187_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand2_1 _07503_ (.A(_01390_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand2_1 _07504_ (.A(_01393_),
    .B(_01248_),
    .Y(_01394_));
 sky130_fd_sc_hd__nand3_1 _07505_ (.A(_01390_),
    .B(_01392_),
    .C(_01247_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _07506_ (.A(_01394_),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__inv_2 _07507_ (.A(_01204_),
    .Y(_01397_));
 sky130_fd_sc_hd__nand2_1 _07508_ (.A(_01196_),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand3_1 _07509_ (.A(_01204_),
    .B(_01193_),
    .C(_01195_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2_1 _07510_ (.A(_01398_),
    .B(_01399_),
    .Y(_01401_));
 sky130_fd_sc_hd__nand2_1 _07511_ (.A(_01401_),
    .B(_01219_),
    .Y(_01402_));
 sky130_fd_sc_hd__nand3_1 _07512_ (.A(_01398_),
    .B(_01399_),
    .C(_01218_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand2_1 _07513_ (.A(_01402_),
    .B(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__inv_2 _07514_ (.A(_01198_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand2_1 _07515_ (.A(_01405_),
    .B(_01197_),
    .Y(_01406_));
 sky130_fd_sc_hd__inv_2 _07516_ (.A(_01197_),
    .Y(_01407_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_01407_),
    .B(_01198_),
    .Y(_01408_));
 sky130_fd_sc_hd__nand3_2 _07518_ (.A(_01406_),
    .B(_01408_),
    .C(_01200_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2_1 _07519_ (.A(_01407_),
    .B(_01405_),
    .Y(_01410_));
 sky130_fd_sc_hd__nand3_2 _07520_ (.A(_01410_),
    .B(_01201_),
    .C(_01199_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _07521_ (.A(_01409_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__nand2_1 _07522_ (.A(_02797_),
    .B(net58),
    .Y(_01414_));
 sky130_fd_sc_hd__nand2_1 _07523_ (.A(_02555_),
    .B(net55),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2_1 _07524_ (.A(_01414_),
    .B(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__nand2_1 _07525_ (.A(_02511_),
    .B(net44),
    .Y(_01417_));
 sky130_fd_sc_hd__inv_2 _07526_ (.A(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _07527_ (.A(_01414_),
    .B(_01415_),
    .Y(_01419_));
 sky130_fd_sc_hd__a21oi_2 _07528_ (.A1(_01416_),
    .A2(_01418_),
    .B1(_01419_),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _07529_ (.A(_01413_),
    .B(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__inv_2 _07530_ (.A(_01340_),
    .Y(_01423_));
 sky130_fd_sc_hd__inv_2 _07531_ (.A(_01341_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand2_1 _07532_ (.A(_01423_),
    .B(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(_01425_),
    .B(_01342_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _07534_ (.A(_01426_),
    .B(_01343_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand3_1 _07535_ (.A(_01425_),
    .B(_01344_),
    .C(_01342_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _07536_ (.A(_01427_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__inv_2 _07537_ (.A(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__nor2_1 _07538_ (.A(_01420_),
    .B(_01413_),
    .Y(_01431_));
 sky130_fd_sc_hd__a21oi_2 _07539_ (.A1(_01421_),
    .A2(_01430_),
    .B1(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _07540_ (.A(_01404_),
    .B(_01432_),
    .Y(_01434_));
 sky130_fd_sc_hd__inv_2 _07541_ (.A(_01347_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand3_1 _07542_ (.A(_01435_),
    .B(_01242_),
    .C(_01338_),
    .Y(_01436_));
 sky130_fd_sc_hd__nand3_1 _07543_ (.A(_01436_),
    .B(_01348_),
    .C(_01359_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _07544_ (.A(_01339_),
    .B(_01435_),
    .Y(_01438_));
 sky130_fd_sc_hd__nand3_1 _07545_ (.A(_01338_),
    .B(_01242_),
    .C(_01347_),
    .Y(_01439_));
 sky130_fd_sc_hd__inv_2 _07546_ (.A(_01359_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand3_1 _07547_ (.A(_01438_),
    .B(_01439_),
    .C(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _07548_ (.A(_01437_),
    .B(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__inv_2 _07549_ (.A(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2_1 _07550_ (.A(_01432_),
    .B(_01404_),
    .Y(_01445_));
 sky130_fd_sc_hd__a21oi_2 _07551_ (.A1(_01434_),
    .A2(_01443_),
    .B1(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand2_1 _07552_ (.A(_01396_),
    .B(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__nor2_1 _07553_ (.A(_01446_),
    .B(_01396_),
    .Y(_01448_));
 sky130_fd_sc_hd__a21oi_2 _07554_ (.A1(_01388_),
    .A2(_01447_),
    .B1(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_1 _07555_ (.A(_01331_),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__o21a_1 _07556_ (.A1(_01336_),
    .A2(_01361_),
    .B1(_01385_),
    .X(_01451_));
 sky130_fd_sc_hd__xor2_2 _07557_ (.A(_01271_),
    .B(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__nor2_1 _07558_ (.A(_01449_),
    .B(_01331_),
    .Y(_01453_));
 sky130_fd_sc_hd__a21oi_2 _07559_ (.A1(_01450_),
    .A2(_01452_),
    .B1(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_1 _07560_ (.A(_01327_),
    .B(_01454_),
    .Y(_01456_));
 sky130_fd_sc_hd__nor2_1 _07561_ (.A(_01271_),
    .B(_01451_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor2_1 _07562_ (.A(_01454_),
    .B(_01327_),
    .Y(_01458_));
 sky130_fd_sc_hd__a21oi_1 _07563_ (.A1(_01456_),
    .A2(_01457_),
    .B1(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__inv_2 _07564_ (.A(_01303_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _07565_ (.A(_01164_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand3_1 _07566_ (.A(_01303_),
    .B(_01160_),
    .C(_01163_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _07567_ (.A(_01461_),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__nand2_1 _07568_ (.A(_01463_),
    .B(_01298_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand3_1 _07569_ (.A(_01461_),
    .B(_01462_),
    .C(_01324_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _07570_ (.A(_01464_),
    .B(_01465_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _07571_ (.A(_01459_),
    .B(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _07572_ (.A(_01311_),
    .B(_01313_),
    .Y(_01469_));
 sky130_fd_sc_hd__a21oi_1 _07573_ (.A1(_01304_),
    .A2(_01298_),
    .B1(_01305_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _07574_ (.A(_01469_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand3_1 _07575_ (.A(_01314_),
    .B(_01468_),
    .C(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__inv_2 _07576_ (.A(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_1 _07577_ (.A(_01470_),
    .B(_01469_),
    .Y(_01474_));
 sky130_fd_sc_hd__nand2_1 _07578_ (.A(_01121_),
    .B(_01123_),
    .Y(_01475_));
 sky130_fd_sc_hd__nand3_1 _07579_ (.A(_01119_),
    .B(_01120_),
    .C(_00956_),
    .Y(_01476_));
 sky130_fd_sc_hd__nand2_1 _07580_ (.A(_01475_),
    .B(_01476_),
    .Y(_01478_));
 sky130_fd_sc_hd__a21o_1 _07581_ (.A1(_01115_),
    .A2(_01109_),
    .B1(_01116_),
    .X(_01479_));
 sky130_fd_sc_hd__nand2_1 _07582_ (.A(_01478_),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2_1 _07583_ (.A(_01126_),
    .B(_01117_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand3_2 _07584_ (.A(_01474_),
    .B(_01480_),
    .C(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _07585_ (.A(_01480_),
    .B(_01481_),
    .Y(_01483_));
 sky130_fd_sc_hd__nand2_1 _07586_ (.A(_01483_),
    .B(_01314_),
    .Y(_01484_));
 sky130_fd_sc_hd__nand3_2 _07587_ (.A(_01473_),
    .B(_01482_),
    .C(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__nand3_1 _07588_ (.A(_00961_),
    .B(_00962_),
    .C(_01480_),
    .Y(_01486_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(_01128_),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__and2_1 _07590_ (.A(_01487_),
    .B(_01482_),
    .X(_01489_));
 sky130_fd_sc_hd__or2_1 _07591_ (.A(_01482_),
    .B(_01487_),
    .X(_01490_));
 sky130_fd_sc_hd__o21ai_1 _07592_ (.A1(_01485_),
    .A2(_01489_),
    .B1(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__nor2_1 _07593_ (.A(_01314_),
    .B(_01483_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _07594_ (.A(_00963_),
    .B(_01480_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand3_1 _07595_ (.A(_01127_),
    .B(_00961_),
    .C(_00962_),
    .Y(_01494_));
 sky130_fd_sc_hd__nand3_1 _07596_ (.A(_01492_),
    .B(_01493_),
    .C(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__nand3_1 _07597_ (.A(_01128_),
    .B(_01486_),
    .C(_01482_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(_01495_),
    .B(_01496_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand2_1 _07599_ (.A(_01484_),
    .B(_01482_),
    .Y(_01498_));
 sky130_fd_sc_hd__nand2_1 _07600_ (.A(_01498_),
    .B(_01472_),
    .Y(_01500_));
 sky130_fd_sc_hd__nand3_1 _07601_ (.A(_01497_),
    .B(_01500_),
    .C(_01485_),
    .Y(_01501_));
 sky130_fd_sc_hd__inv_2 _07602_ (.A(_01454_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand2_1 _07603_ (.A(_01327_),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__nand3_1 _07604_ (.A(_01454_),
    .B(_01322_),
    .C(_01326_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _07605_ (.A(_01503_),
    .B(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__nand2_1 _07606_ (.A(_01505_),
    .B(_01457_),
    .Y(_01506_));
 sky130_fd_sc_hd__inv_2 _07607_ (.A(_01457_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand3_1 _07608_ (.A(_01503_),
    .B(_01504_),
    .C(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__nand2_1 _07609_ (.A(_01506_),
    .B(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__a21o_1 _07610_ (.A1(_01434_),
    .A2(_01443_),
    .B1(_01445_),
    .X(_01511_));
 sky130_fd_sc_hd__nand3_1 _07611_ (.A(_01511_),
    .B(_01394_),
    .C(_01395_),
    .Y(_01512_));
 sky130_fd_sc_hd__nand3_1 _07612_ (.A(_01512_),
    .B(_01388_),
    .C(_01447_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_1 _07613_ (.A(_01396_),
    .B(_01511_),
    .Y(_01514_));
 sky130_fd_sc_hd__nand3_1 _07614_ (.A(_01446_),
    .B(_01394_),
    .C(_01395_),
    .Y(_01515_));
 sky130_fd_sc_hd__nand3_1 _07615_ (.A(_01514_),
    .B(_01515_),
    .C(_01387_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand2_1 _07616_ (.A(_01513_),
    .B(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _07617_ (.A(_01380_),
    .B(_01382_),
    .Y(_01518_));
 sky130_fd_sc_hd__nand2_1 _07618_ (.A(_01518_),
    .B(_01366_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _07619_ (.A(_01519_),
    .B(_01383_),
    .Y(_01520_));
 sky130_fd_sc_hd__nand2_1 _07620_ (.A(_01352_),
    .B(_01349_),
    .Y(_01522_));
 sky130_fd_sc_hd__nand2_1 _07621_ (.A(_01350_),
    .B(_01351_),
    .Y(_01523_));
 sky130_fd_sc_hd__nand3_1 _07622_ (.A(_01522_),
    .B(_01523_),
    .C(_01354_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand2_1 _07623_ (.A(_01524_),
    .B(_01358_),
    .Y(_01525_));
 sky130_fd_sc_hd__nand2_1 _07624_ (.A(_02874_),
    .B(_00641_),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(_02489_),
    .B(_00674_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand2_1 _07626_ (.A(_01526_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__nand2_1 _07627_ (.A(_04634_),
    .B(_00751_),
    .Y(_01529_));
 sky130_fd_sc_hd__inv_2 _07628_ (.A(_01529_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _07629_ (.A(_01526_),
    .B(_01527_),
    .Y(_01531_));
 sky130_fd_sc_hd__a21oi_2 _07630_ (.A1(_01528_),
    .A2(_01530_),
    .B1(_01531_),
    .Y(_01533_));
 sky130_fd_sc_hd__nand2_1 _07631_ (.A(_01525_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__nand2_1 _07632_ (.A(_00893_),
    .B(_05068_),
    .Y(_01535_));
 sky130_fd_sc_hd__nand2_1 _07633_ (.A(_00384_),
    .B(_00315_),
    .Y(_01536_));
 sky130_fd_sc_hd__or2_1 _07634_ (.A(_01535_),
    .B(_01536_),
    .X(_01537_));
 sky130_fd_sc_hd__nand2_1 _07635_ (.A(_04895_),
    .B(_01323_),
    .Y(_01538_));
 sky130_fd_sc_hd__inv_2 _07636_ (.A(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__nand2_1 _07637_ (.A(_01535_),
    .B(_01536_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand3_1 _07638_ (.A(_01537_),
    .B(_01539_),
    .C(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__nand2_1 _07639_ (.A(_01541_),
    .B(_01537_),
    .Y(_01542_));
 sky130_fd_sc_hd__nor2_1 _07640_ (.A(_01533_),
    .B(_01525_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21oi_2 _07641_ (.A1(_01534_),
    .A2(_01542_),
    .B1(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_1 _07642_ (.A(_01520_),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__inv_2 _07643_ (.A(_01545_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand3_2 _07644_ (.A(_01547_),
    .B(_01519_),
    .C(_01383_),
    .Y(_01548_));
 sky130_fd_sc_hd__nand2_1 _07645_ (.A(_01546_),
    .B(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__and4_1 _07646_ (.A(_04947_),
    .B(net1),
    .C(_03039_),
    .D(_02522_),
    .X(_01550_));
 sky130_fd_sc_hd__inv_2 _07647_ (.A(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__nor2b_1 _07648_ (.A(_01377_),
    .B_N(_01374_),
    .Y(_01552_));
 sky130_fd_sc_hd__xor2_1 _07649_ (.A(_01375_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__nor2_1 _07650_ (.A(_01551_),
    .B(_01553_),
    .Y(_01555_));
 sky130_fd_sc_hd__inv_2 _07651_ (.A(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__nand2_1 _07652_ (.A(_01549_),
    .B(_01556_),
    .Y(_01557_));
 sky130_fd_sc_hd__nand3_1 _07653_ (.A(_01546_),
    .B(_01548_),
    .C(_01555_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_1 _07654_ (.A(_01557_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__inv_2 _07655_ (.A(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__nand3_1 _07656_ (.A(_01432_),
    .B(_01402_),
    .C(_01403_),
    .Y(_01561_));
 sky130_fd_sc_hd__inv_2 _07657_ (.A(_01420_),
    .Y(_01562_));
 sky130_fd_sc_hd__nand3_1 _07658_ (.A(_01562_),
    .B(_01412_),
    .C(_01409_),
    .Y(_01563_));
 sky130_fd_sc_hd__nand3_1 _07659_ (.A(_01563_),
    .B(_01421_),
    .C(_01430_),
    .Y(_01564_));
 sky130_fd_sc_hd__nand2_1 _07660_ (.A(_01564_),
    .B(_01563_),
    .Y(_01566_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(_01404_),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__nand2_1 _07662_ (.A(_01561_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand2_1 _07663_ (.A(_01568_),
    .B(_01443_),
    .Y(_01569_));
 sky130_fd_sc_hd__nand3_1 _07664_ (.A(_01561_),
    .B(_01567_),
    .C(_01442_),
    .Y(_01570_));
 sky130_fd_sc_hd__nand2_1 _07665_ (.A(_01569_),
    .B(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__nand2_1 _07666_ (.A(_01413_),
    .B(_01562_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand3_1 _07667_ (.A(_01420_),
    .B(_01409_),
    .C(_01412_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand3_1 _07668_ (.A(_01572_),
    .B(_01573_),
    .C(_01429_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _07669_ (.A(_01564_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__inv_2 _07670_ (.A(_01414_),
    .Y(_01577_));
 sky130_fd_sc_hd__inv_2 _07671_ (.A(_01415_),
    .Y(_01578_));
 sky130_fd_sc_hd__nand2_1 _07672_ (.A(_01577_),
    .B(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(_01579_),
    .B(_01416_),
    .Y(_01580_));
 sky130_fd_sc_hd__nand2_1 _07674_ (.A(_01580_),
    .B(_01418_),
    .Y(_01581_));
 sky130_fd_sc_hd__nand2_1 _07675_ (.A(_02874_),
    .B(_00300_),
    .Y(_01582_));
 sky130_fd_sc_hd__nand2_1 _07676_ (.A(_00138_),
    .B(net55),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _07677_ (.A(_01582_),
    .B(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _07678_ (.A(_02555_),
    .B(_00410_),
    .Y(_01585_));
 sky130_fd_sc_hd__inv_2 _07679_ (.A(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor2_1 _07680_ (.A(_01582_),
    .B(_01583_),
    .Y(_01588_));
 sky130_fd_sc_hd__a21oi_2 _07681_ (.A1(_01584_),
    .A2(_01586_),
    .B1(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__nand3_1 _07682_ (.A(_01579_),
    .B(_01417_),
    .C(_01416_),
    .Y(_01590_));
 sky130_fd_sc_hd__nand3_2 _07683_ (.A(_01581_),
    .B(_01589_),
    .C(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__inv_2 _07684_ (.A(_01531_),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_1 _07685_ (.A(_01592_),
    .B(_01528_),
    .Y(_01593_));
 sky130_fd_sc_hd__nand2_1 _07686_ (.A(_01593_),
    .B(_01530_),
    .Y(_01594_));
 sky130_fd_sc_hd__nand3_1 _07687_ (.A(_01592_),
    .B(_01529_),
    .C(_01528_),
    .Y(_01595_));
 sky130_fd_sc_hd__nand2_2 _07688_ (.A(_01594_),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__nand2_1 _07689_ (.A(_01581_),
    .B(_01590_),
    .Y(_01597_));
 sky130_fd_sc_hd__inv_2 _07690_ (.A(_01589_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand2_2 _07691_ (.A(_01597_),
    .B(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__inv_2 _07692_ (.A(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__a21oi_1 _07693_ (.A1(_01591_),
    .A2(_01596_),
    .B1(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(_01575_),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__inv_2 _07695_ (.A(_01533_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _07696_ (.A(_01525_),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__nand3_1 _07697_ (.A(_01533_),
    .B(_01524_),
    .C(_01358_),
    .Y(_01606_));
 sky130_fd_sc_hd__nand2_1 _07698_ (.A(_01605_),
    .B(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__nand2_1 _07699_ (.A(_01607_),
    .B(_01542_),
    .Y(_01608_));
 sky130_fd_sc_hd__a21boi_1 _07700_ (.A1(_01539_),
    .A2(_01540_),
    .B1_N(_01537_),
    .Y(_01610_));
 sky130_fd_sc_hd__nand3_1 _07701_ (.A(_01605_),
    .B(_01606_),
    .C(_01610_),
    .Y(_01611_));
 sky130_fd_sc_hd__nand2_1 _07702_ (.A(_01608_),
    .B(_01611_),
    .Y(_01612_));
 sky130_fd_sc_hd__inv_2 _07703_ (.A(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hd__nor2_1 _07704_ (.A(_01602_),
    .B(_01575_),
    .Y(_01614_));
 sky130_fd_sc_hd__a21oi_4 _07705_ (.A1(_01603_),
    .A2(_01613_),
    .B1(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__nand2_1 _07706_ (.A(_01571_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__nor2_1 _07707_ (.A(_01615_),
    .B(_01571_),
    .Y(_01617_));
 sky130_fd_sc_hd__a21oi_2 _07708_ (.A1(_01560_),
    .A2(_01616_),
    .B1(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _07709_ (.A(_01517_),
    .B(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__nand2_2 _07710_ (.A(_01558_),
    .B(_01548_),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_1 _07711_ (.A(_01618_),
    .B(_01517_),
    .Y(_01622_));
 sky130_fd_sc_hd__a21o_1 _07712_ (.A1(_01619_),
    .A2(_01621_),
    .B1(_01622_),
    .X(_01623_));
 sky130_fd_sc_hd__nand3_1 _07713_ (.A(_01449_),
    .B(_01318_),
    .C(_01330_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_1 _07714_ (.A(_01513_),
    .B(_01512_),
    .Y(_01625_));
 sky130_fd_sc_hd__nand2_1 _07715_ (.A(_01625_),
    .B(_01331_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _07716_ (.A(_01624_),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__nand2_1 _07717_ (.A(_01627_),
    .B(_01452_),
    .Y(_01628_));
 sky130_fd_sc_hd__nand3b_2 _07718_ (.A_N(_01452_),
    .B(_01624_),
    .C(_01626_),
    .Y(_01629_));
 sky130_fd_sc_hd__nand3_4 _07719_ (.A(_01623_),
    .B(_01628_),
    .C(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__nand2_1 _07720_ (.A(_01509_),
    .B(_01630_),
    .Y(_01632_));
 sky130_fd_sc_hd__nand3b_2 _07721_ (.A_N(_01630_),
    .B(_01506_),
    .C(_01508_),
    .Y(_01633_));
 sky130_fd_sc_hd__inv_2 _07722_ (.A(_01615_),
    .Y(_01634_));
 sky130_fd_sc_hd__nand2_1 _07723_ (.A(_01571_),
    .B(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__nand3_1 _07724_ (.A(_01615_),
    .B(_01569_),
    .C(_01570_),
    .Y(_01636_));
 sky130_fd_sc_hd__nand2_1 _07725_ (.A(_01635_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2_1 _07726_ (.A(_01637_),
    .B(_01560_),
    .Y(_01638_));
 sky130_fd_sc_hd__nand3_1 _07727_ (.A(_01635_),
    .B(_01636_),
    .C(_01559_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_1 _07728_ (.A(_01638_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__inv_2 _07729_ (.A(_01575_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand3_1 _07730_ (.A(_01600_),
    .B(_01591_),
    .C(_01596_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand2_1 _07731_ (.A(_01643_),
    .B(_01600_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _07732_ (.A(_01641_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__nand3_1 _07733_ (.A(_01645_),
    .B(_01613_),
    .C(_01603_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _07734_ (.A(_01641_),
    .B(_01602_),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _07735_ (.A(_01575_),
    .B(_01644_),
    .Y(_01648_));
 sky130_fd_sc_hd__nand3_1 _07736_ (.A(_01647_),
    .B(_01612_),
    .C(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_2 _07737_ (.A(_01646_),
    .B(_01649_),
    .Y(_01650_));
 sky130_fd_sc_hd__inv_2 _07738_ (.A(_01584_),
    .Y(_01651_));
 sky130_fd_sc_hd__nor2_1 _07739_ (.A(_01588_),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _07740_ (.A(_01652_),
    .B(_01585_),
    .Y(_01654_));
 sky130_fd_sc_hd__inv_2 _07741_ (.A(_01582_),
    .Y(_01655_));
 sky130_fd_sc_hd__inv_2 _07742_ (.A(_01583_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _07743_ (.A(_01655_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _07744_ (.A(_01657_),
    .B(_01584_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_1 _07745_ (.A(_01658_),
    .B(_01586_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _07746_ (.A(_05159_),
    .B(_00300_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_00329_),
    .B(_00344_),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _07748_ (.A(_01660_),
    .B(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_1 _07749_ (.A(_02797_),
    .B(_00410_),
    .Y(_01663_));
 sky130_fd_sc_hd__inv_2 _07750_ (.A(_01663_),
    .Y(_01665_));
 sky130_fd_sc_hd__nor2_1 _07751_ (.A(_01660_),
    .B(_01661_),
    .Y(_01666_));
 sky130_fd_sc_hd__a21oi_1 _07752_ (.A1(_01662_),
    .A2(_01665_),
    .B1(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand3_2 _07753_ (.A(_01654_),
    .B(_01659_),
    .C(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__nand2_1 _07754_ (.A(_04634_),
    .B(_00641_),
    .Y(_01669_));
 sky130_fd_sc_hd__inv_2 _07755_ (.A(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _07756_ (.A(_02511_),
    .B(_00674_),
    .Y(_01671_));
 sky130_fd_sc_hd__inv_2 _07757_ (.A(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand2_1 _07758_ (.A(_01670_),
    .B(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__nand2_1 _07759_ (.A(_01669_),
    .B(_01671_),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_1 _07760_ (.A(_01673_),
    .B(_01674_),
    .Y(_01676_));
 sky130_fd_sc_hd__nand2_1 _07761_ (.A(_04814_),
    .B(_00751_),
    .Y(_01677_));
 sky130_fd_sc_hd__nand2_1 _07762_ (.A(_01676_),
    .B(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__inv_2 _07763_ (.A(_01677_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand3_1 _07764_ (.A(_01673_),
    .B(_01679_),
    .C(_01674_),
    .Y(_01680_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(_01678_),
    .B(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hd__inv_2 _07766_ (.A(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__inv_2 _07767_ (.A(_01667_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand2_1 _07768_ (.A(_01652_),
    .B(_01586_),
    .Y(_01684_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(_01658_),
    .B(_01585_),
    .Y(_01685_));
 sky130_fd_sc_hd__nand3_2 _07770_ (.A(_01683_),
    .B(_01684_),
    .C(_01685_),
    .Y(_01687_));
 sky130_fd_sc_hd__a21boi_1 _07771_ (.A1(_01668_),
    .A2(_01682_),
    .B1_N(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__nand2_1 _07772_ (.A(_01600_),
    .B(_01591_),
    .Y(_01689_));
 sky130_fd_sc_hd__inv_2 _07773_ (.A(_01596_),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _07774_ (.A(_01689_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _07775_ (.A(_01691_),
    .B(_01643_),
    .Y(_01692_));
 sky130_fd_sc_hd__nand2_2 _07776_ (.A(_01688_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__nand2_1 _07777_ (.A(_01537_),
    .B(_01540_),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _07778_ (.A(_01694_),
    .B(_01538_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _07779_ (.A(_01695_),
    .B(_01541_),
    .Y(_01696_));
 sky130_fd_sc_hd__a21boi_1 _07780_ (.A1(_01679_),
    .A2(_01674_),
    .B1_N(_01673_),
    .Y(_01698_));
 sky130_fd_sc_hd__nand2_1 _07781_ (.A(_01696_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _07782_ (.A(_01680_),
    .B(_01673_),
    .Y(_01700_));
 sky130_fd_sc_hd__nand3_1 _07783_ (.A(_01695_),
    .B(_01700_),
    .C(_01541_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_1 _07784_ (.A(_01699_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_1 _07785_ (.A(_04880_),
    .B(_01257_),
    .Y(_01703_));
 sky130_fd_sc_hd__inv_2 _07786_ (.A(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _07787_ (.A(_04895_),
    .B(_01224_),
    .Y(_01705_));
 sky130_fd_sc_hd__inv_2 _07788_ (.A(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__nand2_1 _07789_ (.A(_01704_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _07790_ (.A(_04947_),
    .B(_01323_),
    .Y(_01709_));
 sky130_fd_sc_hd__inv_2 _07791_ (.A(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand2_1 _07792_ (.A(_01703_),
    .B(_01705_),
    .Y(_01711_));
 sky130_fd_sc_hd__nand3_1 _07793_ (.A(_01707_),
    .B(_01710_),
    .C(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__nand2_1 _07794_ (.A(_01712_),
    .B(_01707_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2_1 _07795_ (.A(_01702_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__inv_2 _07796_ (.A(_01713_),
    .Y(_01715_));
 sky130_fd_sc_hd__nand3_1 _07797_ (.A(_01699_),
    .B(_01701_),
    .C(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__nand2_2 _07798_ (.A(_01714_),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(_01689_),
    .B(_01596_),
    .Y(_01718_));
 sky130_fd_sc_hd__nand3_1 _07800_ (.A(_01690_),
    .B(_01600_),
    .C(_01591_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _07801_ (.A(_01718_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__nand3_1 _07802_ (.A(_01687_),
    .B(_01668_),
    .C(_01682_),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(_01722_),
    .B(_01687_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_1 _07804_ (.A(_01721_),
    .B(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__a21boi_4 _07805_ (.A1(_01693_),
    .A2(_01717_),
    .B1_N(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(_01650_),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21boi_2 _07807_ (.A1(_01699_),
    .A2(_01713_),
    .B1_N(_01701_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand2_1 _07808_ (.A(_01553_),
    .B(_01551_),
    .Y(_01728_));
 sky130_fd_sc_hd__nand2_1 _07809_ (.A(_01556_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__nor2_1 _07810_ (.A(_01727_),
    .B(_01729_),
    .Y(_01731_));
 sky130_fd_sc_hd__nand2_1 _07811_ (.A(_01729_),
    .B(_01727_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2b_1 _07812_ (.A(_01731_),
    .B_N(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__nor2_1 _07813_ (.A(_01725_),
    .B(_01650_),
    .Y(_01734_));
 sky130_fd_sc_hd__a21oi_2 _07814_ (.A1(_01726_),
    .A2(_01733_),
    .B1(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(_01640_),
    .B(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__nor2_1 _07816_ (.A(_01735_),
    .B(_01640_),
    .Y(_01737_));
 sky130_fd_sc_hd__a21oi_1 _07817_ (.A1(_01736_),
    .A2(_01731_),
    .B1(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__inv_2 _07818_ (.A(_01517_),
    .Y(_01739_));
 sky130_fd_sc_hd__inv_2 _07819_ (.A(_01618_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _07820_ (.A(_01739_),
    .B(_01740_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand3_1 _07821_ (.A(_01742_),
    .B(_01621_),
    .C(_01619_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _07822_ (.A(_01739_),
    .B(_01618_),
    .Y(_01744_));
 sky130_fd_sc_hd__nand2_1 _07823_ (.A(_01740_),
    .B(_01517_),
    .Y(_01745_));
 sky130_fd_sc_hd__inv_2 _07824_ (.A(_01621_),
    .Y(_01746_));
 sky130_fd_sc_hd__nand3_1 _07825_ (.A(_01744_),
    .B(_01745_),
    .C(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_1 _07826_ (.A(_01743_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _07827_ (.A(_01738_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_1 _07828_ (.A(_01629_),
    .B(_01628_),
    .Y(_01750_));
 sky130_fd_sc_hd__a21oi_1 _07829_ (.A1(_01619_),
    .A2(_01621_),
    .B1(_01622_),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_1 _07830_ (.A(_01750_),
    .B(_01751_),
    .Y(_01753_));
 sky130_fd_sc_hd__nand3_4 _07831_ (.A(_01749_),
    .B(_01630_),
    .C(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__inv_2 _07832_ (.A(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__nand3_1 _07833_ (.A(_01632_),
    .B(_01633_),
    .C(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__nand2_1 _07834_ (.A(_01463_),
    .B(_01324_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand3_1 _07835_ (.A(_01461_),
    .B(_01462_),
    .C(_01298_),
    .Y(_01758_));
 sky130_fd_sc_hd__nand2_1 _07836_ (.A(_01757_),
    .B(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__a21o_1 _07837_ (.A1(_01456_),
    .A2(_01457_),
    .B1(_01458_),
    .X(_01760_));
 sky130_fd_sc_hd__nand2_1 _07838_ (.A(_01759_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_1 _07839_ (.A(_01467_),
    .B(_01459_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2_1 _07840_ (.A(_01761_),
    .B(_01762_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_1 _07841_ (.A(_01764_),
    .B(_01633_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_1 _07842_ (.A(_01630_),
    .B(_01509_),
    .Y(_01766_));
 sky130_fd_sc_hd__nand3_1 _07843_ (.A(_01766_),
    .B(_01761_),
    .C(_01762_),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _07844_ (.A(_01765_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _07845_ (.A(_01756_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand2_1 _07846_ (.A(_01314_),
    .B(_01471_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _07847_ (.A(_01770_),
    .B(_01468_),
    .Y(_01771_));
 sky130_fd_sc_hd__nand3_1 _07848_ (.A(_01314_),
    .B(_01761_),
    .C(_01471_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand3_1 _07849_ (.A(_01771_),
    .B(_01767_),
    .C(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__nand2_1 _07850_ (.A(_01770_),
    .B(_01761_),
    .Y(_01775_));
 sky130_fd_sc_hd__nand2_1 _07851_ (.A(_01775_),
    .B(_01472_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor2_1 _07852_ (.A(_01767_),
    .B(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__a21oi_1 _07853_ (.A1(_01769_),
    .A2(_01773_),
    .B1(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _07854_ (.A(_01501_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__nor2_1 _07855_ (.A(_01491_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _07856_ (.A(_01135_),
    .B(_01137_),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _07857_ (.A(_01781_),
    .B(_01128_),
    .Y(_01782_));
 sky130_fd_sc_hd__nand2_1 _07858_ (.A(_01138_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__nand2_1 _07859_ (.A(_01146_),
    .B(_01142_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _07860_ (.A(_01783_),
    .B(_01784_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand3_1 _07861_ (.A(_00513_),
    .B(_00770_),
    .C(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(_01780_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__nor2_1 _07863_ (.A(_01154_),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__inv_2 _07864_ (.A(_01787_),
    .Y(_01790_));
 sky130_fd_sc_hd__inv_2 _07865_ (.A(_01650_),
    .Y(_01791_));
 sky130_fd_sc_hd__nand2_1 _07866_ (.A(_01791_),
    .B(_01725_),
    .Y(_01792_));
 sky130_fd_sc_hd__inv_2 _07867_ (.A(_01725_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _07868_ (.A(_01793_),
    .B(_01650_),
    .Y(_01794_));
 sky130_fd_sc_hd__inv_2 _07869_ (.A(_01733_),
    .Y(_01795_));
 sky130_fd_sc_hd__nand3_1 _07870_ (.A(_01792_),
    .B(_01794_),
    .C(_01795_),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_1 _07871_ (.A(_01791_),
    .B(_01793_),
    .Y(_01798_));
 sky130_fd_sc_hd__nand3_1 _07872_ (.A(_01798_),
    .B(_01733_),
    .C(_01726_),
    .Y(_01799_));
 sky130_fd_sc_hd__nand2_2 _07873_ (.A(_01797_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__a22o_1 _07874_ (.A1(_05310_),
    .A2(_03039_),
    .B1(_04958_),
    .B2(_05096_),
    .X(_01801_));
 sky130_fd_sc_hd__nand2_1 _07875_ (.A(_01551_),
    .B(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__a21o_1 _07876_ (.A1(_01707_),
    .A2(_01711_),
    .B1(_01710_),
    .X(_01803_));
 sky130_fd_sc_hd__nand2_1 _07877_ (.A(_01803_),
    .B(_01712_),
    .Y(_01804_));
 sky130_fd_sc_hd__nand2_1 _07878_ (.A(_04880_),
    .B(_00751_),
    .Y(_01805_));
 sky130_fd_sc_hd__inv_2 _07879_ (.A(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _07880_ (.A(_04814_),
    .B(net59),
    .Y(_01808_));
 sky130_fd_sc_hd__nand2_1 _07881_ (.A(_02555_),
    .B(net33),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_1 _07882_ (.A(_01808_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__inv_2 _07883_ (.A(_01808_),
    .Y(_01811_));
 sky130_fd_sc_hd__inv_2 _07884_ (.A(_01809_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _07885_ (.A(_01811_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__a21boi_2 _07886_ (.A1(_01806_),
    .A2(_01810_),
    .B1_N(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__inv_2 _07887_ (.A(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__nand2_1 _07888_ (.A(_01804_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand3_1 _07889_ (.A(_01803_),
    .B(_01814_),
    .C(_01712_),
    .Y(_01817_));
 sky130_fd_sc_hd__nand2_1 _07890_ (.A(_01816_),
    .B(_01817_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _07891_ (.A(_04947_),
    .B(_01224_),
    .Y(_01820_));
 sky130_fd_sc_hd__inv_2 _07892_ (.A(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _07893_ (.A(_04895_),
    .B(_05068_),
    .Y(_01822_));
 sky130_fd_sc_hd__inv_2 _07894_ (.A(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__nand2_1 _07895_ (.A(_01821_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand2_1 _07896_ (.A(_01820_),
    .B(_01822_),
    .Y(_01825_));
 sky130_fd_sc_hd__nand2_1 _07897_ (.A(_04958_),
    .B(_01323_),
    .Y(_01826_));
 sky130_fd_sc_hd__inv_2 _07898_ (.A(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__nand3_1 _07899_ (.A(_01824_),
    .B(_01825_),
    .C(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__nand2_1 _07900_ (.A(_01828_),
    .B(_01824_),
    .Y(_01830_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(_01819_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__or2_1 _07902_ (.A(_01814_),
    .B(_01804_),
    .X(_01832_));
 sky130_fd_sc_hd__and2_1 _07903_ (.A(_01831_),
    .B(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__or2_2 _07904_ (.A(_01802_),
    .B(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__nand2_1 _07905_ (.A(_01833_),
    .B(_01802_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2_1 _07906_ (.A(_01834_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__inv_2 _07907_ (.A(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__nand2_1 _07908_ (.A(_01687_),
    .B(_01668_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _07909_ (.A(_01838_),
    .B(_01681_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _07910_ (.A(_01839_),
    .B(_01722_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _07911_ (.A(_01813_),
    .B(_01810_),
    .Y(_01842_));
 sky130_fd_sc_hd__nand2_1 _07912_ (.A(_01842_),
    .B(_01805_),
    .Y(_01843_));
 sky130_fd_sc_hd__nand3_1 _07913_ (.A(_01813_),
    .B(_01806_),
    .C(_01810_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_1 _07914_ (.A(_01843_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__inv_2 _07915_ (.A(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__inv_2 _07916_ (.A(_01660_),
    .Y(_01847_));
 sky130_fd_sc_hd__inv_2 _07917_ (.A(_01661_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _07918_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__nand2_1 _07919_ (.A(_01849_),
    .B(_01662_),
    .Y(_01850_));
 sky130_fd_sc_hd__inv_2 _07920_ (.A(_01850_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _07921_ (.A(_01852_),
    .B(_01663_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_1 _07922_ (.A(_01850_),
    .B(_01665_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand2_1 _07923_ (.A(_05159_),
    .B(_00344_),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _07924_ (.A(_00893_),
    .B(_00300_),
    .Y(_01856_));
 sky130_fd_sc_hd__nand2_1 _07925_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__nand2_1 _07926_ (.A(_00329_),
    .B(_00410_),
    .Y(_01858_));
 sky130_fd_sc_hd__inv_2 _07927_ (.A(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _07928_ (.A(_01855_),
    .B(_01856_),
    .Y(_01860_));
 sky130_fd_sc_hd__a21oi_1 _07929_ (.A1(_01857_),
    .A2(_01859_),
    .B1(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__nand3_1 _07930_ (.A(_01853_),
    .B(_01854_),
    .C(_01861_),
    .Y(_01863_));
 sky130_fd_sc_hd__a21oi_1 _07931_ (.A1(_01853_),
    .A2(_01854_),
    .B1(_01861_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21oi_1 _07932_ (.A1(_01846_),
    .A2(_01863_),
    .B1(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _07933_ (.A(_01841_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__inv_2 _07934_ (.A(_01830_),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _07935_ (.A(_01819_),
    .B(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__nand3_1 _07936_ (.A(_01816_),
    .B(_01817_),
    .C(_01830_),
    .Y(_01869_));
 sky130_fd_sc_hd__nand2_1 _07937_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _07938_ (.A(_01865_),
    .B(_01841_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21oi_1 _07939_ (.A1(_01866_),
    .A2(_01870_),
    .B1(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_1 _07940_ (.A(_01693_),
    .B(_01724_),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2_1 _07941_ (.A(_01874_),
    .B(_01717_),
    .Y(_01875_));
 sky130_fd_sc_hd__inv_2 _07942_ (.A(_01717_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand3_1 _07943_ (.A(_01876_),
    .B(_01693_),
    .C(_01724_),
    .Y(_01877_));
 sky130_fd_sc_hd__nand3_2 _07944_ (.A(_01872_),
    .B(_01875_),
    .C(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _07945_ (.A(_01852_),
    .B(_01665_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand2_1 _07946_ (.A(_01850_),
    .B(_01663_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand3b_2 _07947_ (.A_N(_01861_),
    .B(_01879_),
    .C(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand3_1 _07948_ (.A(_01881_),
    .B(_01863_),
    .C(_01846_),
    .Y(_01882_));
 sky130_fd_sc_hd__nand2_1 _07949_ (.A(_01882_),
    .B(_01881_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand2_1 _07950_ (.A(_01838_),
    .B(_01682_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand3_1 _07951_ (.A(_01687_),
    .B(_01668_),
    .C(_01681_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _07952_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_1 _07953_ (.A(_01883_),
    .B(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand3_1 _07954_ (.A(_01888_),
    .B(_01866_),
    .C(_01870_),
    .Y(_01889_));
 sky130_fd_sc_hd__nand2_1 _07955_ (.A(_01889_),
    .B(_01888_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _07956_ (.A(_01875_),
    .B(_01877_),
    .Y(_01891_));
 sky130_fd_sc_hd__nand2_1 _07957_ (.A(_01890_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__a21boi_4 _07958_ (.A1(_01837_),
    .A2(_01878_),
    .B1_N(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(_01800_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__inv_2 _07960_ (.A(_01834_),
    .Y(_01896_));
 sky130_fd_sc_hd__nor2_1 _07961_ (.A(_01893_),
    .B(_01800_),
    .Y(_01897_));
 sky130_fd_sc_hd__a21oi_1 _07962_ (.A1(_01894_),
    .A2(_01896_),
    .B1(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__nand3_1 _07963_ (.A(_01735_),
    .B(_01638_),
    .C(_01639_),
    .Y(_01899_));
 sky130_fd_sc_hd__inv_2 _07964_ (.A(_01735_),
    .Y(_01900_));
 sky130_fd_sc_hd__nand2_1 _07965_ (.A(_01900_),
    .B(_01640_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _07966_ (.A(_01899_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__nand2_1 _07967_ (.A(_01902_),
    .B(_01731_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand3b_1 _07968_ (.A_N(_01731_),
    .B(_01899_),
    .C(_01901_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand3_1 _07969_ (.A(_01898_),
    .B(_01903_),
    .C(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__a21o_1 _07970_ (.A1(_01894_),
    .A2(_01896_),
    .B1(_01897_),
    .X(_01907_));
 sky130_fd_sc_hd__nand2_1 _07971_ (.A(_01903_),
    .B(_01904_),
    .Y(_01908_));
 sky130_fd_sc_hd__nand2_1 _07972_ (.A(_01907_),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__nand2_1 _07973_ (.A(_01905_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(_01888_),
    .B(_01866_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand3_1 _07975_ (.A(_01816_),
    .B(_01817_),
    .C(_01867_),
    .Y(_01912_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(_01831_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2_1 _07977_ (.A(_01911_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__nand2_1 _07978_ (.A(_01914_),
    .B(_01889_),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _07979_ (.A(_01881_),
    .B(_01863_),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_1 _07980_ (.A(_01916_),
    .B(_01845_),
    .Y(_01918_));
 sky130_fd_sc_hd__nand2_1 _07981_ (.A(_01918_),
    .B(_01882_),
    .Y(_01919_));
 sky130_fd_sc_hd__nand2_1 _07982_ (.A(_04880_),
    .B(_00641_),
    .Y(_01920_));
 sky130_fd_sc_hd__nand2_1 _07983_ (.A(_00138_),
    .B(_00674_),
    .Y(_01921_));
 sky130_fd_sc_hd__nor2_1 _07984_ (.A(_01920_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__inv_2 _07985_ (.A(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand2_1 _07986_ (.A(_01920_),
    .B(_01921_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _07987_ (.A(_01923_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(_04895_),
    .B(_00751_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _07989_ (.A(_01925_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__inv_2 _07990_ (.A(_01926_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand3_1 _07991_ (.A(_01923_),
    .B(_01929_),
    .C(_01924_),
    .Y(_01930_));
 sky130_fd_sc_hd__nand2_1 _07992_ (.A(_01927_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__inv_2 _07993_ (.A(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__inv_2 _07994_ (.A(_01855_),
    .Y(_01933_));
 sky130_fd_sc_hd__inv_2 _07995_ (.A(_01856_),
    .Y(_01934_));
 sky130_fd_sc_hd__nand2_1 _07996_ (.A(_01933_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_1 _07997_ (.A(_01935_),
    .B(_01857_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_1 _07998_ (.A(_01936_),
    .B(_01858_),
    .Y(_01937_));
 sky130_fd_sc_hd__nand3_1 _07999_ (.A(_01935_),
    .B(_01857_),
    .C(_01859_),
    .Y(_01938_));
 sky130_fd_sc_hd__nand2_1 _08000_ (.A(_01937_),
    .B(_01938_),
    .Y(_01940_));
 sky130_fd_sc_hd__nand2_1 _08001_ (.A(_00893_),
    .B(_00344_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand2_1 _08002_ (.A(_00384_),
    .B(_00300_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _08003_ (.A(_01941_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_1 _08004_ (.A(_05159_),
    .B(_00410_),
    .Y(_01944_));
 sky130_fd_sc_hd__inv_2 _08005_ (.A(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__nor2_1 _08006_ (.A(_01941_),
    .B(_01942_),
    .Y(_01946_));
 sky130_fd_sc_hd__a21oi_1 _08007_ (.A1(_01943_),
    .A2(_01945_),
    .B1(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _08008_ (.A(_01940_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__inv_2 _08009_ (.A(_01947_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand3_2 _08010_ (.A(_01949_),
    .B(_01938_),
    .C(_01937_),
    .Y(_01951_));
 sky130_fd_sc_hd__a21boi_1 _08011_ (.A1(_01932_),
    .A2(_01948_),
    .B1_N(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__nand2_1 _08012_ (.A(_01919_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__a21o_1 _08013_ (.A1(_01824_),
    .A2(_01825_),
    .B1(_01827_),
    .X(_01954_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(_01954_),
    .B(_01828_),
    .Y(_01955_));
 sky130_fd_sc_hd__a21oi_2 _08015_ (.A1(_01924_),
    .A2(_01929_),
    .B1(_01922_),
    .Y(_01956_));
 sky130_fd_sc_hd__inv_2 _08016_ (.A(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _08017_ (.A(_01955_),
    .B(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__nand3_1 _08018_ (.A(_01954_),
    .B(_01828_),
    .C(_01956_),
    .Y(_01959_));
 sky130_fd_sc_hd__nand2_1 _08019_ (.A(_01958_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__nand2_1 _08020_ (.A(net1),
    .B(_00315_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor3_1 _08021_ (.A(_00187_),
    .B(_00560_),
    .C(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__inv_2 _08022_ (.A(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _08023_ (.A(_01960_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__nand3_1 _08024_ (.A(_01958_),
    .B(_01963_),
    .C(_01959_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _08025_ (.A(_01965_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _08026_ (.A(_01952_),
    .B(_01919_),
    .Y(_01968_));
 sky130_fd_sc_hd__a21oi_1 _08027_ (.A1(_01953_),
    .A2(_01967_),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(_01915_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _08029_ (.A(_00194_),
    .B(_03039_),
    .Y(_01971_));
 sky130_fd_sc_hd__or2_1 _08030_ (.A(_01956_),
    .B(_01955_),
    .X(_01973_));
 sky130_fd_sc_hd__inv_2 _08031_ (.A(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__and2_1 _08032_ (.A(_01960_),
    .B(_01963_),
    .X(_01975_));
 sky130_fd_sc_hd__nor2_1 _08033_ (.A(_01974_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__nand2b_1 _08034_ (.A_N(_01971_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__o21ai_1 _08035_ (.A1(_01974_),
    .A2(_01975_),
    .B1(_01971_),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _08036_ (.A(_01977_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _08037_ (.A(_01969_),
    .B(_01915_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21oi_1 _08038_ (.A1(_01970_),
    .A2(_01979_),
    .B1(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__nand2_1 _08039_ (.A(_01878_),
    .B(_01892_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand2_1 _08040_ (.A(_01982_),
    .B(_01837_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand3_1 _08041_ (.A(_01878_),
    .B(_01892_),
    .C(_01836_),
    .Y(_01985_));
 sky130_fd_sc_hd__nand3_1 _08042_ (.A(_01981_),
    .B(_01984_),
    .C(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_1 _08043_ (.A(_01984_),
    .B(_01985_),
    .Y(_01987_));
 sky130_fd_sc_hd__a21o_1 _08044_ (.A1(_01953_),
    .A2(_01967_),
    .B1(_01968_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_1 _08045_ (.A(_01911_),
    .B(_01870_),
    .Y(_01989_));
 sky130_fd_sc_hd__nand3_1 _08046_ (.A(_01888_),
    .B(_01866_),
    .C(_01913_),
    .Y(_01990_));
 sky130_fd_sc_hd__nand2_1 _08047_ (.A(_01989_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _08048_ (.A(_01988_),
    .B(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand3_1 _08049_ (.A(_01992_),
    .B(_01970_),
    .C(_01979_),
    .Y(_01993_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_01993_),
    .B(_01992_),
    .Y(_01995_));
 sky130_fd_sc_hd__nand2_1 _08051_ (.A(_01987_),
    .B(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__nor2_1 _08052_ (.A(_01971_),
    .B(_01976_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand3_2 _08053_ (.A(_01986_),
    .B(_01996_),
    .C(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_2 _08054_ (.A(_01998_),
    .B(_01996_),
    .Y(_01999_));
 sky130_fd_sc_hd__inv_2 _08055_ (.A(_01800_),
    .Y(_02000_));
 sky130_fd_sc_hd__inv_2 _08056_ (.A(_01893_),
    .Y(_02001_));
 sky130_fd_sc_hd__nand2_1 _08057_ (.A(_02000_),
    .B(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__nand3_1 _08058_ (.A(_02002_),
    .B(_01896_),
    .C(_01894_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _08059_ (.A(_02000_),
    .B(_01893_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand2_1 _08060_ (.A(_02001_),
    .B(_01800_),
    .Y(_02006_));
 sky130_fd_sc_hd__nand3_1 _08061_ (.A(_02004_),
    .B(_01834_),
    .C(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__nand3_2 _08062_ (.A(_01999_),
    .B(_02003_),
    .C(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__inv_2 _08063_ (.A(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_2 _08064_ (.A(_01910_),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__a21o_1 _08065_ (.A1(_01736_),
    .A2(_01731_),
    .B1(_01737_),
    .X(_02011_));
 sky130_fd_sc_hd__nand3_1 _08066_ (.A(_02011_),
    .B(_01743_),
    .C(_01747_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand2_1 _08067_ (.A(_01748_),
    .B(_01738_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_1 _08068_ (.A(_02012_),
    .B(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__nor2_1 _08069_ (.A(_01898_),
    .B(_01908_),
    .Y(_02015_));
 sky130_fd_sc_hd__inv_2 _08070_ (.A(_02015_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand2_1 _08071_ (.A(_02014_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__nand3_1 _08072_ (.A(_02015_),
    .B(_02012_),
    .C(_02013_),
    .Y(_02019_));
 sky130_fd_sc_hd__nand2_1 _08073_ (.A(_02018_),
    .B(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _08074_ (.A(_02010_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_1 _08075_ (.A(_01630_),
    .B(_01753_),
    .Y(_02022_));
 sky130_fd_sc_hd__nand2_1 _08076_ (.A(_02022_),
    .B(_02012_),
    .Y(_02023_));
 sky130_fd_sc_hd__nand2_1 _08077_ (.A(_02023_),
    .B(_01754_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(_02024_),
    .B(_02019_),
    .Y(_02025_));
 sky130_fd_sc_hd__nor2_1 _08079_ (.A(_02017_),
    .B(_02014_),
    .Y(_02026_));
 sky130_fd_sc_hd__nand3_2 _08080_ (.A(_02026_),
    .B(_02023_),
    .C(_01754_),
    .Y(_02028_));
 sky130_fd_sc_hd__nand3_2 _08081_ (.A(_02021_),
    .B(_02025_),
    .C(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand2_1 _08082_ (.A(_01632_),
    .B(_01633_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _08083_ (.A(_02030_),
    .B(_01755_),
    .Y(_02031_));
 sky130_fd_sc_hd__nand3_1 _08084_ (.A(_01632_),
    .B(_01633_),
    .C(_01754_),
    .Y(_02032_));
 sky130_fd_sc_hd__nand3_1 _08085_ (.A(_02031_),
    .B(_02032_),
    .C(_02028_),
    .Y(_02033_));
 sky130_fd_sc_hd__inv_2 _08086_ (.A(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(_02030_),
    .B(_01754_),
    .Y(_02035_));
 sky130_fd_sc_hd__inv_2 _08088_ (.A(_02028_),
    .Y(_02036_));
 sky130_fd_sc_hd__nand3_1 _08089_ (.A(_02035_),
    .B(_01756_),
    .C(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__o21ai_1 _08090_ (.A1(_02029_),
    .A2(_02034_),
    .B1(_02037_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2_1 _08091_ (.A(_01986_),
    .B(_01996_),
    .Y(_02040_));
 sky130_fd_sc_hd__inv_2 _08092_ (.A(_01997_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _08093_ (.A(_02040_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_1 _08094_ (.A(_02042_),
    .B(_01998_),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _08095_ (.A(_04895_),
    .B(_00641_),
    .Y(_02044_));
 sky130_fd_sc_hd__inv_2 _08096_ (.A(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__nand2_1 _08097_ (.A(_00329_),
    .B(_00674_),
    .Y(_02046_));
 sky130_fd_sc_hd__inv_2 _08098_ (.A(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__nand2_1 _08099_ (.A(_02045_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand2_1 _08100_ (.A(_02044_),
    .B(_02046_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _08101_ (.A(_04947_),
    .B(_00751_),
    .Y(_02051_));
 sky130_fd_sc_hd__inv_2 _08102_ (.A(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__a21o_1 _08103_ (.A1(_02048_),
    .A2(_02050_),
    .B1(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__nand3_1 _08104_ (.A(_02048_),
    .B(_02052_),
    .C(_02050_),
    .Y(_02054_));
 sky130_fd_sc_hd__nand2_1 _08105_ (.A(_02053_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__inv_2 _08106_ (.A(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__or2b_1 _08107_ (.A(_01946_),
    .B_N(_01943_),
    .X(_02057_));
 sky130_fd_sc_hd__nand2_1 _08108_ (.A(_02057_),
    .B(_01945_),
    .Y(_02058_));
 sky130_fd_sc_hd__and2b_1 _08109_ (.A_N(_01946_),
    .B(_01943_),
    .X(_02059_));
 sky130_fd_sc_hd__nand2_1 _08110_ (.A(_02059_),
    .B(_01944_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _08111_ (.A(_00384_),
    .B(_00344_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _08112_ (.A(_04895_),
    .B(_00300_),
    .Y(_02063_));
 sky130_fd_sc_hd__nand2_1 _08113_ (.A(_02062_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__nand2_1 _08114_ (.A(_00893_),
    .B(_00410_),
    .Y(_02065_));
 sky130_fd_sc_hd__inv_2 _08115_ (.A(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _08116_ (.A(_02062_),
    .B(_02063_),
    .Y(_02067_));
 sky130_fd_sc_hd__a21oi_1 _08117_ (.A1(_02064_),
    .A2(_02066_),
    .B1(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand3_1 _08118_ (.A(_02058_),
    .B(_02061_),
    .C(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__nand2_1 _08119_ (.A(_02057_),
    .B(_01944_),
    .Y(_02070_));
 sky130_fd_sc_hd__nand2_1 _08120_ (.A(_02059_),
    .B(_01945_),
    .Y(_02072_));
 sky130_fd_sc_hd__nand3b_2 _08121_ (.A_N(_02068_),
    .B(_02070_),
    .C(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__a21boi_1 _08122_ (.A1(_02056_),
    .A2(_02069_),
    .B1_N(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2_1 _08123_ (.A(_01951_),
    .B(_01948_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_1 _08124_ (.A(_02075_),
    .B(_01931_),
    .Y(_02076_));
 sky130_fd_sc_hd__nand3_1 _08125_ (.A(_01951_),
    .B(_01932_),
    .C(_01948_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_1 _08126_ (.A(_02076_),
    .B(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand2_1 _08127_ (.A(_02074_),
    .B(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__o21ai_1 _08128_ (.A1(_00187_),
    .A2(_00560_),
    .B1(_01962_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _08129_ (.A(_01964_),
    .B(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__and2_1 _08130_ (.A(_02054_),
    .B(_02048_),
    .X(_02083_));
 sky130_fd_sc_hd__nor2_1 _08131_ (.A(_02081_),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__inv_2 _08132_ (.A(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_1 _08133_ (.A(_02083_),
    .B(_02081_),
    .Y(_02086_));
 sky130_fd_sc_hd__and2_1 _08134_ (.A(_02085_),
    .B(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__nor2_1 _08135_ (.A(_02078_),
    .B(_02074_),
    .Y(_02088_));
 sky130_fd_sc_hd__a21oi_1 _08136_ (.A1(_02079_),
    .A2(_02087_),
    .B1(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__inv_2 _08137_ (.A(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand2_1 _08138_ (.A(_02077_),
    .B(_01951_),
    .Y(_02091_));
 sky130_fd_sc_hd__nand3_1 _08139_ (.A(_02091_),
    .B(_01882_),
    .C(_01918_),
    .Y(_02092_));
 sky130_fd_sc_hd__nand2_1 _08140_ (.A(_02092_),
    .B(_01953_),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_1 _08141_ (.A(_02094_),
    .B(_01967_),
    .Y(_02095_));
 sky130_fd_sc_hd__nand3b_1 _08142_ (.A_N(_01967_),
    .B(_02092_),
    .C(_01953_),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_1 _08143_ (.A(_02095_),
    .B(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _08144_ (.A(_02090_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__nand3_1 _08145_ (.A(_02089_),
    .B(_02096_),
    .C(_02095_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand3_1 _08146_ (.A(_02098_),
    .B(_02099_),
    .C(_02084_),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_1 _08147_ (.A(_02100_),
    .B(_02098_),
    .Y(_02101_));
 sky130_fd_sc_hd__nand2_1 _08148_ (.A(_01992_),
    .B(_01970_),
    .Y(_02102_));
 sky130_fd_sc_hd__nand3_1 _08149_ (.A(_02102_),
    .B(_01977_),
    .C(_01978_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand3_2 _08150_ (.A(_02101_),
    .B(_01993_),
    .C(_02103_),
    .Y(_02105_));
 sky130_fd_sc_hd__nand2_1 _08151_ (.A(_02043_),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__inv_2 _08152_ (.A(_02105_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand3_4 _08153_ (.A(_02042_),
    .B(_01998_),
    .C(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_1 _08154_ (.A(_02098_),
    .B(_02099_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _08155_ (.A(_02109_),
    .B(_02085_),
    .Y(_02110_));
 sky130_fd_sc_hd__nand2_1 _08156_ (.A(_02110_),
    .B(_02100_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand2_1 _08157_ (.A(_00381_),
    .B(_00232_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _08158_ (.A(_05310_),
    .B(_00234_),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_1 _08159_ (.A(_02112_),
    .B(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__nand2_1 _08160_ (.A(_00384_),
    .B(_00433_),
    .Y(_02116_));
 sky130_fd_sc_hd__inv_2 _08161_ (.A(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _08162_ (.A(_02112_),
    .B(_02113_),
    .Y(_02118_));
 sky130_fd_sc_hd__a21o_1 _08163_ (.A1(_02114_),
    .A2(_02117_),
    .B1(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__inv_2 _08164_ (.A(_02062_),
    .Y(_02120_));
 sky130_fd_sc_hd__inv_2 _08165_ (.A(_02063_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _08166_ (.A(_02120_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(_02122_),
    .B(_02064_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2b_1 _08168_ (.A_N(_02123_),
    .B(_02065_),
    .Y(_02124_));
 sky130_fd_sc_hd__nand2_1 _08169_ (.A(_02123_),
    .B(_02066_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand3b_1 _08170_ (.A_N(_02119_),
    .B(_02124_),
    .C(_02125_),
    .Y(_02127_));
 sky130_fd_sc_hd__nand2_1 _08171_ (.A(_04947_),
    .B(_00641_),
    .Y(_02128_));
 sky130_fd_sc_hd__nand2_1 _08172_ (.A(_05159_),
    .B(_00674_),
    .Y(_02129_));
 sky130_fd_sc_hd__or2_1 _08173_ (.A(_02128_),
    .B(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__nand2_1 _08174_ (.A(_02128_),
    .B(_02129_),
    .Y(_02131_));
 sky130_fd_sc_hd__nand2_1 _08175_ (.A(_02130_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _08176_ (.A(_04958_),
    .B(_00306_),
    .Y(_02133_));
 sky130_fd_sc_hd__or2b_1 _08177_ (.A(_02132_),
    .B_N(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__a21o_1 _08178_ (.A1(_02130_),
    .A2(_02131_),
    .B1(_02133_),
    .X(_02135_));
 sky130_fd_sc_hd__nand2_1 _08179_ (.A(_02134_),
    .B(_02135_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _08180_ (.A(_02124_),
    .B(_02125_),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2_1 _08181_ (.A(_02138_),
    .B(_02119_),
    .Y(_02139_));
 sky130_fd_sc_hd__a21boi_1 _08182_ (.A1(_02127_),
    .A2(_02136_),
    .B1_N(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__nand2_1 _08183_ (.A(_02073_),
    .B(_02069_),
    .Y(_02141_));
 sky130_fd_sc_hd__nand2_1 _08184_ (.A(_02141_),
    .B(_02055_),
    .Y(_02142_));
 sky130_fd_sc_hd__nand3_1 _08185_ (.A(_02073_),
    .B(_02069_),
    .C(_02056_),
    .Y(_02143_));
 sky130_fd_sc_hd__nand2_1 _08186_ (.A(_02142_),
    .B(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__nand2_1 _08187_ (.A(_02140_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand2_1 _08188_ (.A(_04958_),
    .B(_05068_),
    .Y(_02146_));
 sky130_fd_sc_hd__o21a_1 _08189_ (.A1(_02133_),
    .A2(_02132_),
    .B1(_02130_),
    .X(_02147_));
 sky130_fd_sc_hd__nor2_1 _08190_ (.A(_02146_),
    .B(_02147_),
    .Y(_02149_));
 sky130_fd_sc_hd__inv_2 _08191_ (.A(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_1 _08192_ (.A(_02147_),
    .B(_02146_),
    .Y(_02151_));
 sky130_fd_sc_hd__nand2_1 _08193_ (.A(_02150_),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__inv_2 _08194_ (.A(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__nor2_1 _08195_ (.A(_02144_),
    .B(_02140_),
    .Y(_02154_));
 sky130_fd_sc_hd__a21oi_1 _08196_ (.A1(_02145_),
    .A2(_02153_),
    .B1(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _08197_ (.A(_02143_),
    .B(_02073_),
    .Y(_02156_));
 sky130_fd_sc_hd__nand2_1 _08198_ (.A(_02075_),
    .B(_01932_),
    .Y(_02157_));
 sky130_fd_sc_hd__nand3_1 _08199_ (.A(_01951_),
    .B(_01948_),
    .C(_01931_),
    .Y(_02158_));
 sky130_fd_sc_hd__nand2_1 _08200_ (.A(_02157_),
    .B(_02158_),
    .Y(_02160_));
 sky130_fd_sc_hd__nand2_1 _08201_ (.A(_02156_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__nand2_1 _08202_ (.A(_02079_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__nand2_1 _08203_ (.A(_02162_),
    .B(_02087_),
    .Y(_02163_));
 sky130_fd_sc_hd__nand3b_1 _08204_ (.A_N(_02087_),
    .B(_02079_),
    .C(_02161_),
    .Y(_02164_));
 sky130_fd_sc_hd__nand3_1 _08205_ (.A(_02155_),
    .B(_02163_),
    .C(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__inv_2 _08206_ (.A(_02155_),
    .Y(_02166_));
 sky130_fd_sc_hd__nand2_1 _08207_ (.A(_02163_),
    .B(_02164_),
    .Y(_02167_));
 sky130_fd_sc_hd__nand2_1 _08208_ (.A(_02166_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__a21boi_1 _08209_ (.A1(_02165_),
    .A2(_02149_),
    .B1_N(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__nor2_1 _08210_ (.A(_02111_),
    .B(_02169_),
    .Y(_02171_));
 sky130_fd_sc_hd__inv_2 _08211_ (.A(_02101_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _08212_ (.A(_02103_),
    .B(_01993_),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _08213_ (.A(_02172_),
    .B(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand3_2 _08214_ (.A(_02171_),
    .B(_02105_),
    .C(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__inv_2 _08215_ (.A(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__nand3_4 _08216_ (.A(_02106_),
    .B(_02108_),
    .C(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_02003_),
    .B(_02007_),
    .Y(_02178_));
 sky130_fd_sc_hd__inv_2 _08218_ (.A(_01999_),
    .Y(_02179_));
 sky130_fd_sc_hd__nand2_1 _08219_ (.A(_02178_),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_1 _08220_ (.A(_02180_),
    .B(_02008_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_1 _08221_ (.A(_02182_),
    .B(_02108_),
    .Y(_02183_));
 sky130_fd_sc_hd__nand3b_2 _08222_ (.A_N(_02108_),
    .B(_02180_),
    .C(_02008_),
    .Y(_02184_));
 sky130_fd_sc_hd__nand3b_2 _08223_ (.A_N(_02177_),
    .B(_02183_),
    .C(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__nor2_1 _08224_ (.A(_02108_),
    .B(_02182_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand3_1 _08225_ (.A(_02008_),
    .B(_01905_),
    .C(_01909_),
    .Y(_02187_));
 sky130_fd_sc_hd__nand3_2 _08226_ (.A(_02186_),
    .B(_02010_),
    .C(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _08227_ (.A(_02010_),
    .B(_02187_),
    .Y(_02189_));
 sky130_fd_sc_hd__nand2_1 _08228_ (.A(_02189_),
    .B(_02184_),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _08229_ (.A(_02188_),
    .B(_02190_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(_02185_),
    .B(_02191_),
    .Y(_02193_));
 sky130_fd_sc_hd__inv_2 _08231_ (.A(_02010_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand3_1 _08232_ (.A(_02194_),
    .B(_02019_),
    .C(_02018_),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(_02020_),
    .B(_02010_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _08234_ (.A(_02195_),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _08235_ (.A(_02197_),
    .B(_02188_),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _08236_ (.A(_02188_),
    .B(_02197_),
    .Y(_02199_));
 sky130_fd_sc_hd__a21oi_1 _08237_ (.A1(_02193_),
    .A2(_02198_),
    .B1(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__nand2_1 _08238_ (.A(_02025_),
    .B(_02028_),
    .Y(_02201_));
 sky130_fd_sc_hd__nand2_1 _08239_ (.A(_02201_),
    .B(_02195_),
    .Y(_02202_));
 sky130_fd_sc_hd__nand2_1 _08240_ (.A(_02202_),
    .B(_02029_),
    .Y(_02204_));
 sky130_fd_sc_hd__inv_2 _08241_ (.A(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__nand3_1 _08242_ (.A(_02205_),
    .B(_02037_),
    .C(_02033_),
    .Y(_02206_));
 sky130_fd_sc_hd__nor2_1 _08243_ (.A(_02200_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__nor2_1 _08244_ (.A(_02039_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__nand2_1 _08245_ (.A(_02106_),
    .B(_02108_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_1 _08246_ (.A(_02209_),
    .B(_02175_),
    .Y(_02210_));
 sky130_fd_sc_hd__nand2_1 _08247_ (.A(_02210_),
    .B(_02177_),
    .Y(_02211_));
 sky130_fd_sc_hd__a21o_1 _08248_ (.A1(_02165_),
    .A2(_02168_),
    .B1(_02149_),
    .X(_02212_));
 sky130_fd_sc_hd__nand3_1 _08249_ (.A(_02165_),
    .B(_02168_),
    .C(_02149_),
    .Y(_02213_));
 sky130_fd_sc_hd__nand2_1 _08250_ (.A(_02127_),
    .B(_02139_),
    .Y(_02215_));
 sky130_fd_sc_hd__nand3_1 _08251_ (.A(_02215_),
    .B(_02135_),
    .C(_02134_),
    .Y(_02216_));
 sky130_fd_sc_hd__nand3_1 _08252_ (.A(_02127_),
    .B(_02139_),
    .C(_02136_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _08253_ (.A(_02216_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2b_1 _08254_ (.A_N(_02118_),
    .B(_02114_),
    .Y(_02219_));
 sky130_fd_sc_hd__xor2_1 _08255_ (.A(_02117_),
    .B(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__a22o_1 _08256_ (.A1(_05310_),
    .A2(_00232_),
    .B1(_00194_),
    .B2(_00234_),
    .X(_02221_));
 sky130_fd_sc_hd__nand2_1 _08257_ (.A(_00381_),
    .B(_00433_),
    .Y(_02222_));
 sky130_fd_sc_hd__inv_2 _08258_ (.A(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__and4_1 _08259_ (.A(_05310_),
    .B(_00194_),
    .C(_00234_),
    .D(_00232_),
    .X(_02224_));
 sky130_fd_sc_hd__a21oi_1 _08260_ (.A1(_02221_),
    .A2(_02223_),
    .B1(_02224_),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _08261_ (.A(_02220_),
    .B(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__and4_1 _08262_ (.A(_00893_),
    .B(_00194_),
    .C(_00303_),
    .D(_00301_),
    .X(_02228_));
 sky130_fd_sc_hd__inv_2 _08263_ (.A(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__a22o_1 _08264_ (.A1(_00893_),
    .A2(_00303_),
    .B1(_00194_),
    .B2(_00301_),
    .X(_02230_));
 sky130_fd_sc_hd__and2_1 _08265_ (.A(_02229_),
    .B(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__nor2_1 _08266_ (.A(_02226_),
    .B(_02220_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21oi_1 _08267_ (.A1(_02227_),
    .A2(_02231_),
    .B1(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__nand2_1 _08268_ (.A(_02218_),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _08269_ (.A(_02233_),
    .B(_02218_),
    .Y(_02235_));
 sky130_fd_sc_hd__a21oi_1 _08270_ (.A1(_02234_),
    .A2(_02228_),
    .B1(_02235_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2b_1 _08271_ (.A_N(_02154_),
    .B(_02145_),
    .Y(_02238_));
 sky130_fd_sc_hd__xor2_1 _08272_ (.A(_02153_),
    .B(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__nor2_1 _08273_ (.A(_02237_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand3_2 _08274_ (.A(_02212_),
    .B(_02213_),
    .C(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _08275_ (.A(_02213_),
    .B(_02168_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand3_1 _08276_ (.A(_02242_),
    .B(_02100_),
    .C(_02110_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand2_1 _08277_ (.A(_02169_),
    .B(_02111_),
    .Y(_02244_));
 sky130_fd_sc_hd__nand2_1 _08278_ (.A(_02243_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _08279_ (.A(_02241_),
    .B(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_1 _08280_ (.A(_02105_),
    .B(_02174_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand2_1 _08281_ (.A(_02248_),
    .B(_02243_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand3_2 _08282_ (.A(_02246_),
    .B(_02249_),
    .C(_02175_),
    .Y(_02250_));
 sky130_fd_sc_hd__nand2_1 _08283_ (.A(_02211_),
    .B(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__inv_2 _08284_ (.A(_02250_),
    .Y(_02252_));
 sky130_fd_sc_hd__nand3_4 _08285_ (.A(_02210_),
    .B(_02252_),
    .C(_02177_),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_1 _08286_ (.A(_02251_),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__nand2_1 _08287_ (.A(_02249_),
    .B(_02175_),
    .Y(_02255_));
 sky130_fd_sc_hd__inv_2 _08288_ (.A(_02241_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand3_1 _08289_ (.A(_02256_),
    .B(_02243_),
    .C(_02244_),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_1 _08290_ (.A(_02255_),
    .B(_02257_),
    .Y(_02259_));
 sky130_fd_sc_hd__nand2_1 _08291_ (.A(_02250_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__nand2_1 _08292_ (.A(_02212_),
    .B(_02213_),
    .Y(_02261_));
 sky130_fd_sc_hd__inv_2 _08293_ (.A(_02240_),
    .Y(_02262_));
 sky130_fd_sc_hd__nand2_1 _08294_ (.A(_02261_),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__nand2_1 _08295_ (.A(_02263_),
    .B(_02241_),
    .Y(_02264_));
 sky130_fd_sc_hd__inv_2 _08296_ (.A(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2b_1 _08297_ (.A_N(_02235_),
    .B(_02234_),
    .Y(_02266_));
 sky130_fd_sc_hd__or2_1 _08298_ (.A(_02229_),
    .B(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__nand2_1 _08299_ (.A(_02266_),
    .B(_02229_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand2b_1 _08300_ (.A_N(_02232_),
    .B(_02227_),
    .Y(_02270_));
 sky130_fd_sc_hd__xor2_1 _08301_ (.A(_02231_),
    .B(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__inv_2 _08302_ (.A(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__inv_2 _08303_ (.A(_02221_),
    .Y(_02273_));
 sky130_fd_sc_hd__or3_1 _08304_ (.A(_02222_),
    .B(_02224_),
    .C(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__o21ai_1 _08305_ (.A1(_02224_),
    .A2(_02273_),
    .B1(_02222_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_1 _08306_ (.A(_02274_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__nand2_1 _08307_ (.A(_05310_),
    .B(_00433_),
    .Y(_02277_));
 sky130_fd_sc_hd__inv_2 _08308_ (.A(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__and3_1 _08309_ (.A(_02278_),
    .B(_00194_),
    .C(_00232_),
    .X(_02279_));
 sky130_fd_sc_hd__inv_2 _08310_ (.A(_02279_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_1 _08311_ (.A(_02276_),
    .B(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__nand3_1 _08312_ (.A(_02274_),
    .B(_02275_),
    .C(_02279_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _08313_ (.A(_00384_),
    .B(_00303_),
    .Y(_02284_));
 sky130_fd_sc_hd__inv_2 _08314_ (.A(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__nand3_1 _08315_ (.A(_02282_),
    .B(_02283_),
    .C(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__nand2_1 _08316_ (.A(_02286_),
    .B(_02283_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand2_1 _08317_ (.A(_02272_),
    .B(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__inv_2 _08318_ (.A(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand3_2 _08319_ (.A(_02267_),
    .B(_02268_),
    .C(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _08320_ (.A(_02239_),
    .B(_02237_),
    .Y(_02292_));
 sky130_fd_sc_hd__nand2_1 _08321_ (.A(_02262_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__nor2_1 _08322_ (.A(_02290_),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_1 _08323_ (.A(_02265_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__nand2_1 _08324_ (.A(_02245_),
    .B(_02241_),
    .Y(_02296_));
 sky130_fd_sc_hd__nand2_1 _08325_ (.A(_02257_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _08326_ (.A(_02295_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2b_1 _08327_ (.A(_02260_),
    .B_N(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__inv_2 _08328_ (.A(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__nand2_1 _08329_ (.A(_02254_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__nand3_1 _08330_ (.A(_02299_),
    .B(_02251_),
    .C(_02253_),
    .Y(_02303_));
 sky130_fd_sc_hd__xor2_1 _08331_ (.A(_02228_),
    .B(_02266_),
    .X(_02304_));
 sky130_fd_sc_hd__nand2_1 _08332_ (.A(_02304_),
    .B(_02288_),
    .Y(_02305_));
 sky130_fd_sc_hd__a21o_1 _08333_ (.A1(_02282_),
    .A2(_02283_),
    .B1(_02285_),
    .X(_02306_));
 sky130_fd_sc_hd__nand2_1 _08334_ (.A(_02306_),
    .B(_02286_),
    .Y(_02307_));
 sky130_fd_sc_hd__inv_2 _08335_ (.A(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__inv_2 _08336_ (.A(_00381_),
    .Y(_02309_));
 sky130_fd_sc_hd__inv_2 _08337_ (.A(_00674_),
    .Y(_02310_));
 sky130_fd_sc_hd__inv_2 _08338_ (.A(_04958_),
    .Y(_02311_));
 sky130_fd_sc_hd__inv_2 _08339_ (.A(_00232_),
    .Y(_02312_));
 sky130_fd_sc_hd__o21ai_1 _08340_ (.A1(_02311_),
    .A2(_02312_),
    .B1(_02277_),
    .Y(_02314_));
 sky130_fd_sc_hd__nand2_1 _08341_ (.A(_02281_),
    .B(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__or3_1 _08342_ (.A(_02309_),
    .B(_02310_),
    .C(_02315_),
    .X(_02316_));
 sky130_fd_sc_hd__inv_2 _08343_ (.A(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__nand2_1 _08344_ (.A(_02308_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__or2_1 _08345_ (.A(_02287_),
    .B(_02272_),
    .X(_02319_));
 sky130_fd_sc_hd__nand2_1 _08346_ (.A(_02319_),
    .B(_02288_),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _08347_ (.A(_02318_),
    .B(_02320_),
    .Y(_02321_));
 sky130_fd_sc_hd__a21o_1 _08348_ (.A1(_02305_),
    .A2(_02290_),
    .B1(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__nand3_1 _08349_ (.A(_02321_),
    .B(_02305_),
    .C(_02290_),
    .Y(_02323_));
 sky130_fd_sc_hd__o21ai_1 _08350_ (.A1(_02309_),
    .A2(_02310_),
    .B1(_02315_),
    .Y(_02325_));
 sky130_fd_sc_hd__and3_1 _08351_ (.A(_02278_),
    .B(_00194_),
    .C(_00303_),
    .X(_02326_));
 sky130_fd_sc_hd__and3_1 _08352_ (.A(_02316_),
    .B(_02325_),
    .C(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__nand3b_1 _08353_ (.A_N(_02320_),
    .B(_02308_),
    .C(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_02323_),
    .B(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _08355_ (.A(_02293_),
    .B(_02290_),
    .Y(_02330_));
 sky130_fd_sc_hd__and4_1 _08356_ (.A(_02265_),
    .B(_02322_),
    .C(_02329_),
    .D(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__nand2_1 _08357_ (.A(_02297_),
    .B(_02295_),
    .Y(_02332_));
 sky130_fd_sc_hd__nand2_1 _08358_ (.A(_02331_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__nor2_1 _08359_ (.A(_02260_),
    .B(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__nand3_1 _08360_ (.A(_02301_),
    .B(_02303_),
    .C(_02334_),
    .Y(_02336_));
 sky130_fd_sc_hd__nand2_1 _08361_ (.A(_02336_),
    .B(_02303_),
    .Y(_02337_));
 sky130_fd_sc_hd__nand2_1 _08362_ (.A(_02183_),
    .B(_02184_),
    .Y(_02338_));
 sky130_fd_sc_hd__nand2_1 _08363_ (.A(_02338_),
    .B(_02177_),
    .Y(_02339_));
 sky130_fd_sc_hd__a21o_1 _08364_ (.A1(_02339_),
    .A2(_02185_),
    .B1(_02253_),
    .X(_02340_));
 sky130_fd_sc_hd__and2_1 _08365_ (.A(_02339_),
    .B(_02185_),
    .X(_02341_));
 sky130_fd_sc_hd__nand2_1 _08366_ (.A(_02341_),
    .B(_02253_),
    .Y(_02342_));
 sky130_fd_sc_hd__nand2_1 _08367_ (.A(_02340_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__nand2_1 _08368_ (.A(_02337_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__nand2b_1 _08369_ (.A_N(_02253_),
    .B(_02341_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand2_1 _08370_ (.A(_02344_),
    .B(_02345_),
    .Y(_02347_));
 sky130_fd_sc_hd__inv_2 _08371_ (.A(_02188_),
    .Y(_02348_));
 sky130_fd_sc_hd__nand2_1 _08372_ (.A(_02197_),
    .B(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hd__nand3_1 _08373_ (.A(_02188_),
    .B(_02195_),
    .C(_02196_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2_1 _08374_ (.A(_02349_),
    .B(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__inv_2 _08375_ (.A(_02193_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _08376_ (.A(_02191_),
    .B(_02185_),
    .Y(_02353_));
 sky130_fd_sc_hd__nand3_1 _08377_ (.A(_02351_),
    .B(_02352_),
    .C(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _08378_ (.A(_02354_),
    .B(_02206_),
    .Y(_02355_));
 sky130_fd_sc_hd__nand2_1 _08379_ (.A(_02347_),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__nand2_1 _08380_ (.A(_02208_),
    .B(_02356_),
    .Y(_02358_));
 sky130_fd_sc_hd__inv_4 _08381_ (.A(_01769_),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _08382_ (.A(_01768_),
    .B(_01756_),
    .Y(_02360_));
 sky130_fd_sc_hd__nand2_1 _08383_ (.A(_02359_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__nor2_1 _08384_ (.A(_01633_),
    .B(_01764_),
    .Y(_02362_));
 sky130_fd_sc_hd__xor2_2 _08385_ (.A(_02362_),
    .B(_01776_),
    .X(_02363_));
 sky130_fd_sc_hd__nor3_1 _08386_ (.A(_02361_),
    .B(_02363_),
    .C(_01501_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand3_1 _08387_ (.A(_01790_),
    .B(_02358_),
    .C(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _08388_ (.A(_01789_),
    .B(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _08389_ (.A(_01521_),
    .B(_04645_),
    .Y(_02367_));
 sky130_fd_sc_hd__inv_2 _08390_ (.A(net5),
    .Y(_02369_));
 sky130_fd_sc_hd__nand2_1 _08391_ (.A(_01334_),
    .B(_05114_),
    .Y(_02370_));
 sky130_fd_sc_hd__nor3_1 _08392_ (.A(_01267_),
    .B(_02369_),
    .C(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__o21ai_2 _08393_ (.A1(_01267_),
    .A2(_02369_),
    .B1(_02370_),
    .Y(_02372_));
 sky130_fd_sc_hd__inv_2 _08394_ (.A(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__nor2_1 _08395_ (.A(_02371_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__xor2_1 _08396_ (.A(_02367_),
    .B(_02374_),
    .X(_02375_));
 sky130_fd_sc_hd__inv_2 _08397_ (.A(net64),
    .Y(_02376_));
 sky130_fd_sc_hd__inv_2 _08398_ (.A(_00960_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_1 _08399_ (.A(_05096_),
    .B(_04128_),
    .Y(_02378_));
 sky130_fd_sc_hd__o21ai_1 _08400_ (.A1(_02376_),
    .A2(_02377_),
    .B1(_02378_),
    .Y(_02380_));
 sky130_fd_sc_hd__nand2_1 _08401_ (.A(_02687_),
    .B(_02214_),
    .Y(_02381_));
 sky130_fd_sc_hd__inv_2 _08402_ (.A(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor3_1 _08403_ (.A(_02376_),
    .B(_02377_),
    .C(_02378_),
    .Y(_02383_));
 sky130_fd_sc_hd__a21oi_1 _08404_ (.A1(_02380_),
    .A2(_02382_),
    .B1(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__inv_2 _08405_ (.A(_00520_),
    .Y(_02385_));
 sky130_fd_sc_hd__nand2_1 _08406_ (.A(_05096_),
    .B(_00960_),
    .Y(_02386_));
 sky130_fd_sc_hd__nor3_1 _08407_ (.A(_02376_),
    .B(_02385_),
    .C(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__o21ai_2 _08408_ (.A1(_02376_),
    .A2(_02385_),
    .B1(_02386_),
    .Y(_02388_));
 sky130_fd_sc_hd__inv_2 _08409_ (.A(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__nand2_1 _08410_ (.A(_02687_),
    .B(_04128_),
    .Y(_02391_));
 sky130_fd_sc_hd__o21ai_1 _08411_ (.A1(_02387_),
    .A2(_02389_),
    .B1(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__inv_2 _08412_ (.A(_02391_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand3b_1 _08413_ (.A_N(_02387_),
    .B(_02393_),
    .C(_02388_),
    .Y(_02394_));
 sky130_fd_sc_hd__nand2_1 _08414_ (.A(_02392_),
    .B(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__or2_1 _08415_ (.A(_02384_),
    .B(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(_02395_),
    .B(_02384_),
    .Y(_02397_));
 sky130_fd_sc_hd__nand3b_1 _08417_ (.A_N(_02375_),
    .B(_02396_),
    .C(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__inv_2 _08418_ (.A(_02384_),
    .Y(_02399_));
 sky130_fd_sc_hd__or2_1 _08419_ (.A(_02399_),
    .B(_02395_),
    .X(_02400_));
 sky130_fd_sc_hd__nand2_1 _08420_ (.A(_02395_),
    .B(_02399_),
    .Y(_02402_));
 sky130_fd_sc_hd__nand3_1 _08421_ (.A(_02400_),
    .B(_02375_),
    .C(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__nand2_1 _08422_ (.A(_02398_),
    .B(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__nand2_1 _08423_ (.A(_02203_),
    .B(_00520_),
    .Y(_02405_));
 sky130_fd_sc_hd__nand2_1 _08424_ (.A(_00315_),
    .B(_00311_),
    .Y(_02406_));
 sky130_fd_sc_hd__nand2_1 _08425_ (.A(_05068_),
    .B(_00355_),
    .Y(_02407_));
 sky130_fd_sc_hd__or2_1 _08426_ (.A(_02406_),
    .B(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__nand2_1 _08427_ (.A(_02406_),
    .B(_02407_),
    .Y(_02409_));
 sky130_fd_sc_hd__nand2_1 _08428_ (.A(_02408_),
    .B(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__or2_1 _08429_ (.A(_02405_),
    .B(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__nand2_1 _08430_ (.A(_02410_),
    .B(_02405_),
    .Y(_02413_));
 sky130_fd_sc_hd__nand2_1 _08431_ (.A(_02411_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__nand2_1 _08432_ (.A(_00535_),
    .B(_00528_),
    .Y(_02415_));
 sky130_fd_sc_hd__inv_2 _08433_ (.A(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__nand2_1 _08434_ (.A(_02414_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__nand2_1 _08435_ (.A(_00568_),
    .B(_00559_),
    .Y(_02418_));
 sky130_fd_sc_hd__nor2_1 _08436_ (.A(_02416_),
    .B(_02414_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21oi_2 _08437_ (.A1(_02417_),
    .A2(_02418_),
    .B1(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__inv_2 _08438_ (.A(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__nand2_1 _08439_ (.A(_02404_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__nand3_1 _08440_ (.A(_02398_),
    .B(_02403_),
    .C(_02420_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_1 _08441_ (.A(_02422_),
    .B(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__nand2_1 _08442_ (.A(_00611_),
    .B(_00605_),
    .Y(_02426_));
 sky130_fd_sc_hd__inv_2 _08443_ (.A(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__inv_2 _08444_ (.A(_02383_),
    .Y(_02428_));
 sky130_fd_sc_hd__nand2_1 _08445_ (.A(_02428_),
    .B(_02380_),
    .Y(_02429_));
 sky130_fd_sc_hd__or2b_1 _08446_ (.A(_02429_),
    .B_N(_02382_),
    .X(_02430_));
 sky130_fd_sc_hd__nand2_1 _08447_ (.A(_02429_),
    .B(_02381_),
    .Y(_02431_));
 sky130_fd_sc_hd__nand2_1 _08448_ (.A(_02430_),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_1 _08449_ (.A(_02432_),
    .B(_02426_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand3_1 _08450_ (.A(_02430_),
    .B(_02427_),
    .C(_02431_),
    .Y(_02435_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(_02433_),
    .B(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__inv_2 _08452_ (.A(net4),
    .Y(_02437_));
 sky130_fd_sc_hd__nand2_1 _08453_ (.A(_01521_),
    .B(_05114_),
    .Y(_02438_));
 sky130_fd_sc_hd__or3_1 _08454_ (.A(_02437_),
    .B(_01267_),
    .C(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__o21ai_1 _08455_ (.A1(_02437_),
    .A2(_01267_),
    .B1(_02438_),
    .Y(_02440_));
 sky130_fd_sc_hd__nand2_1 _08456_ (.A(_03105_),
    .B(_04645_),
    .Y(_02441_));
 sky130_fd_sc_hd__inv_2 _08457_ (.A(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__a21o_1 _08458_ (.A1(_02439_),
    .A2(_02440_),
    .B1(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__nor3_1 _08459_ (.A(_02437_),
    .B(_01267_),
    .C(_02438_),
    .Y(_02444_));
 sky130_fd_sc_hd__nand3b_1 _08460_ (.A_N(_02444_),
    .B(_02442_),
    .C(_02440_),
    .Y(_02446_));
 sky130_fd_sc_hd__nand2_1 _08461_ (.A(_02443_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__inv_2 _08462_ (.A(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__nand2_1 _08463_ (.A(_02436_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__o21ai_2 _08464_ (.A1(_02427_),
    .A2(_02432_),
    .B1(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__nand2_1 _08465_ (.A(_02425_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__nand3b_1 _08466_ (.A_N(_02450_),
    .B(_02422_),
    .C(_02424_),
    .Y(_02452_));
 sky130_fd_sc_hd__nand2_1 _08467_ (.A(_02451_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__inv_2 _08468_ (.A(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__nand2_1 _08469_ (.A(_00433_),
    .B(_00526_),
    .Y(_02455_));
 sky130_fd_sc_hd__nand2_1 _08470_ (.A(_00344_),
    .B(_05049_),
    .Y(_02457_));
 sky130_fd_sc_hd__nand2_1 _08471_ (.A(_00234_),
    .B(_01895_),
    .Y(_02458_));
 sky130_fd_sc_hd__or2_1 _08472_ (.A(_02457_),
    .B(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__nand2_1 _08473_ (.A(_02457_),
    .B(_02458_),
    .Y(_02460_));
 sky130_fd_sc_hd__nand2_1 _08474_ (.A(_02459_),
    .B(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__or2_1 _08475_ (.A(_02455_),
    .B(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__nand2_1 _08476_ (.A(_02461_),
    .B(_02455_),
    .Y(_02463_));
 sky130_fd_sc_hd__nand2_1 _08477_ (.A(_02462_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _08478_ (.A(_00545_),
    .B(_00539_),
    .Y(_02465_));
 sky130_fd_sc_hd__inv_2 _08479_ (.A(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__nand2_1 _08480_ (.A(_02464_),
    .B(_02466_),
    .Y(_02468_));
 sky130_fd_sc_hd__nand2_1 _08481_ (.A(_00306_),
    .B(_00421_),
    .Y(_02469_));
 sky130_fd_sc_hd__nand2_1 _08482_ (.A(_00301_),
    .B(_00685_),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_1 _08483_ (.A(_00303_),
    .B(net17),
    .Y(_02471_));
 sky130_fd_sc_hd__or2_1 _08484_ (.A(_02470_),
    .B(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__nand2_1 _08485_ (.A(_02470_),
    .B(_02471_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand2_1 _08486_ (.A(_02472_),
    .B(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__or2_1 _08487_ (.A(_02469_),
    .B(_02474_),
    .X(_02475_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(_02474_),
    .B(_02469_),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_1 _08489_ (.A(_02475_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__inv_2 _08490_ (.A(_02477_),
    .Y(_02479_));
 sky130_fd_sc_hd__nand3_1 _08491_ (.A(_02462_),
    .B(_02465_),
    .C(_02463_),
    .Y(_02480_));
 sky130_fd_sc_hd__nand3_1 _08492_ (.A(_02468_),
    .B(_02479_),
    .C(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__nand2_1 _08493_ (.A(_02481_),
    .B(_02480_),
    .Y(_02482_));
 sky130_fd_sc_hd__nand2_1 _08494_ (.A(_00433_),
    .B(net17),
    .Y(_02483_));
 sky130_fd_sc_hd__nand2_1 _08495_ (.A(_00344_),
    .B(_00526_),
    .Y(_02484_));
 sky130_fd_sc_hd__nand2_1 _08496_ (.A(_00300_),
    .B(_05049_),
    .Y(_02485_));
 sky130_fd_sc_hd__or2_1 _08497_ (.A(_02484_),
    .B(_02485_),
    .X(_02486_));
 sky130_fd_sc_hd__nand2_1 _08498_ (.A(_02484_),
    .B(_02485_),
    .Y(_02487_));
 sky130_fd_sc_hd__nand2_1 _08499_ (.A(_02486_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__or2_1 _08500_ (.A(_02483_),
    .B(_02488_),
    .X(_02490_));
 sky130_fd_sc_hd__nand2_1 _08501_ (.A(_02488_),
    .B(_02483_),
    .Y(_02491_));
 sky130_fd_sc_hd__nand2_1 _08502_ (.A(_02490_),
    .B(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__o21ai_1 _08503_ (.A1(_02455_),
    .A2(_02461_),
    .B1(_02459_),
    .Y(_02493_));
 sky130_fd_sc_hd__inv_2 _08504_ (.A(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__nand2_1 _08505_ (.A(_02492_),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand3_1 _08506_ (.A(_02493_),
    .B(_02490_),
    .C(_02491_),
    .Y(_02496_));
 sky130_fd_sc_hd__nand2_1 _08507_ (.A(_02495_),
    .B(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__inv_2 _08508_ (.A(net18),
    .Y(_02498_));
 sky130_fd_sc_hd__nand2_1 _08509_ (.A(_00301_),
    .B(_01895_),
    .Y(_02499_));
 sky130_fd_sc_hd__nor3_1 _08510_ (.A(_02310_),
    .B(_02498_),
    .C(_02499_),
    .Y(_02501_));
 sky130_fd_sc_hd__inv_2 _08511_ (.A(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__o21ai_1 _08512_ (.A1(_02310_),
    .A2(_02498_),
    .B1(_02499_),
    .Y(_02503_));
 sky130_fd_sc_hd__nand2_1 _08513_ (.A(_02502_),
    .B(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__nand2_1 _08514_ (.A(_00306_),
    .B(_00685_),
    .Y(_02505_));
 sky130_fd_sc_hd__inv_2 _08515_ (.A(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__nand2b_1 _08516_ (.A_N(_02504_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _08517_ (.A(_02504_),
    .B(_02505_),
    .Y(_02508_));
 sky130_fd_sc_hd__nand2_1 _08518_ (.A(_02507_),
    .B(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__nand2_1 _08519_ (.A(_02497_),
    .B(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__inv_2 _08520_ (.A(_02509_),
    .Y(_02512_));
 sky130_fd_sc_hd__nand3_1 _08521_ (.A(_02512_),
    .B(_02495_),
    .C(_02496_),
    .Y(_02513_));
 sky130_fd_sc_hd__nand3_2 _08522_ (.A(_02482_),
    .B(_02510_),
    .C(_02513_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand2_1 _08523_ (.A(_02510_),
    .B(_02513_),
    .Y(_02515_));
 sky130_fd_sc_hd__a21boi_1 _08524_ (.A1(_02468_),
    .A2(_02479_),
    .B1_N(_02480_),
    .Y(_02516_));
 sky130_fd_sc_hd__nand2_1 _08525_ (.A(_02515_),
    .B(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(_02514_),
    .B(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__inv_2 _08527_ (.A(_00421_),
    .Y(_02519_));
 sky130_fd_sc_hd__nand2_1 _08528_ (.A(_00315_),
    .B(_00355_),
    .Y(_02520_));
 sky130_fd_sc_hd__or3_1 _08529_ (.A(_00560_),
    .B(_02519_),
    .C(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__o21ai_1 _08530_ (.A1(_00560_),
    .A2(_02519_),
    .B1(_02520_),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _08531_ (.A(_02521_),
    .B(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand2_1 _08532_ (.A(_02203_),
    .B(_00311_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand2_1 _08533_ (.A(_02524_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__nand3b_1 _08534_ (.A_N(_02525_),
    .B(_02521_),
    .C(_02523_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2_1 _08535_ (.A(_02526_),
    .B(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__o21a_1 _08536_ (.A1(_02469_),
    .A2(_02474_),
    .B1(_02472_),
    .X(_02529_));
 sky130_fd_sc_hd__inv_2 _08537_ (.A(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__nand2_1 _08538_ (.A(_02528_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand3_1 _08539_ (.A(_02526_),
    .B(_02527_),
    .C(_02529_),
    .Y(_02532_));
 sky130_fd_sc_hd__nand2_1 _08540_ (.A(_02531_),
    .B(_02532_),
    .Y(_02534_));
 sky130_fd_sc_hd__nand2_1 _08541_ (.A(_02411_),
    .B(_02408_),
    .Y(_02535_));
 sky130_fd_sc_hd__nand2_1 _08542_ (.A(_02534_),
    .B(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__nand3b_1 _08543_ (.A_N(_02535_),
    .B(_02531_),
    .C(_02532_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2_1 _08544_ (.A(_02536_),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2_1 _08545_ (.A(_02518_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__inv_2 _08546_ (.A(_02538_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand3_2 _08547_ (.A(_02540_),
    .B(_02514_),
    .C(_02517_),
    .Y(_02541_));
 sky130_fd_sc_hd__nand2_1 _08548_ (.A(_02539_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_1 _08549_ (.A(_02468_),
    .B(_02480_),
    .Y(_02543_));
 sky130_fd_sc_hd__nand2_1 _08550_ (.A(_02543_),
    .B(_02477_),
    .Y(_02545_));
 sky130_fd_sc_hd__nand2_1 _08551_ (.A(_02545_),
    .B(_02481_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand2_1 _08552_ (.A(_00551_),
    .B(_00550_),
    .Y(_02547_));
 sky130_fd_sc_hd__inv_2 _08553_ (.A(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__nand2_1 _08554_ (.A(_02546_),
    .B(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2_1 _08555_ (.A(_02414_),
    .B(_02415_),
    .Y(_02550_));
 sky130_fd_sc_hd__nand3_1 _08556_ (.A(_02416_),
    .B(_02411_),
    .C(_02413_),
    .Y(_02551_));
 sky130_fd_sc_hd__nand2_1 _08557_ (.A(_02550_),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(_02552_),
    .B(_02418_),
    .Y(_02553_));
 sky130_fd_sc_hd__nand3b_1 _08559_ (.A_N(_02418_),
    .B(_02550_),
    .C(_02551_),
    .Y(_02554_));
 sky130_fd_sc_hd__nand2_1 _08560_ (.A(_02553_),
    .B(_02554_),
    .Y(_02556_));
 sky130_fd_sc_hd__inv_2 _08561_ (.A(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__nand3_1 _08562_ (.A(_02545_),
    .B(_02547_),
    .C(_02481_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand3_1 _08563_ (.A(_02549_),
    .B(_02557_),
    .C(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_1 _08564_ (.A(_02559_),
    .B(_02558_),
    .Y(_02560_));
 sky130_fd_sc_hd__inv_2 _08565_ (.A(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__nand2_1 _08566_ (.A(_02542_),
    .B(_02561_),
    .Y(_02562_));
 sky130_fd_sc_hd__nand3_2 _08567_ (.A(_02560_),
    .B(_02539_),
    .C(_02541_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand3_2 _08568_ (.A(_02454_),
    .B(_02562_),
    .C(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__nand2_1 _08569_ (.A(_02564_),
    .B(_02563_),
    .Y(_02565_));
 sky130_fd_sc_hd__nand2_1 _08570_ (.A(_02541_),
    .B(_02514_),
    .Y(_02567_));
 sky130_fd_sc_hd__nand2_1 _08571_ (.A(_02490_),
    .B(_02486_),
    .Y(_02568_));
 sky130_fd_sc_hd__nand2_1 _08572_ (.A(_00433_),
    .B(net18),
    .Y(_02569_));
 sky130_fd_sc_hd__nand2_1 _08573_ (.A(_00344_),
    .B(net17),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _08574_ (.A(_00300_),
    .B(_00526_),
    .Y(_02571_));
 sky130_fd_sc_hd__or2_1 _08575_ (.A(_02570_),
    .B(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__nand2_1 _08576_ (.A(_02570_),
    .B(_02571_),
    .Y(_02573_));
 sky130_fd_sc_hd__nand2_1 _08577_ (.A(_02572_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__or2_1 _08578_ (.A(_02569_),
    .B(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_1 _08579_ (.A(_02574_),
    .B(_02569_),
    .Y(_02576_));
 sky130_fd_sc_hd__nand3_1 _08580_ (.A(_02568_),
    .B(_02575_),
    .C(_02576_),
    .Y(_02578_));
 sky130_fd_sc_hd__nand2_1 _08581_ (.A(_02575_),
    .B(_02576_),
    .Y(_02579_));
 sky130_fd_sc_hd__o21a_1 _08582_ (.A1(_02483_),
    .A2(_02488_),
    .B1(_02486_),
    .X(_02580_));
 sky130_fd_sc_hd__nand2_1 _08583_ (.A(_02579_),
    .B(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__nand2_1 _08584_ (.A(_02578_),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__inv_2 _08585_ (.A(net19),
    .Y(_02583_));
 sky130_fd_sc_hd__nand2_1 _08586_ (.A(_00301_),
    .B(_05049_),
    .Y(_02584_));
 sky130_fd_sc_hd__nor3_1 _08587_ (.A(_02310_),
    .B(_02583_),
    .C(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__o21ai_2 _08588_ (.A1(_02310_),
    .A2(_02583_),
    .B1(_02584_),
    .Y(_02586_));
 sky130_fd_sc_hd__inv_2 _08589_ (.A(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand2_1 _08590_ (.A(_00306_),
    .B(_01895_),
    .Y(_02589_));
 sky130_fd_sc_hd__o21ai_1 _08591_ (.A1(_02585_),
    .A2(_02587_),
    .B1(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__inv_2 _08592_ (.A(_02589_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand3b_1 _08593_ (.A_N(_02585_),
    .B(_02591_),
    .C(_02586_),
    .Y(_02592_));
 sky130_fd_sc_hd__nand2_1 _08594_ (.A(_02590_),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__nand2_1 _08595_ (.A(_02582_),
    .B(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__inv_2 _08596_ (.A(_02593_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand3_1 _08597_ (.A(_02578_),
    .B(_02595_),
    .C(_02581_),
    .Y(_02596_));
 sky130_fd_sc_hd__nand2_1 _08598_ (.A(_02594_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__a21boi_1 _08599_ (.A1(_02512_),
    .A2(_02495_),
    .B1_N(_02496_),
    .Y(_02598_));
 sky130_fd_sc_hd__nand2_1 _08600_ (.A(_02597_),
    .B(_02598_),
    .Y(_02600_));
 sky130_fd_sc_hd__nand2_1 _08601_ (.A(_02513_),
    .B(_02496_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand3_2 _08602_ (.A(_02601_),
    .B(_02594_),
    .C(_02596_),
    .Y(_02602_));
 sky130_fd_sc_hd__nand2_1 _08603_ (.A(_02600_),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__nand2_1 _08604_ (.A(_02527_),
    .B(_02521_),
    .Y(_02604_));
 sky130_fd_sc_hd__nand2_1 _08605_ (.A(_02203_),
    .B(_00355_),
    .Y(_02605_));
 sky130_fd_sc_hd__inv_2 _08606_ (.A(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__nand2_1 _08607_ (.A(_00315_),
    .B(_00421_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand2_1 _08608_ (.A(_05068_),
    .B(_00685_),
    .Y(_02608_));
 sky130_fd_sc_hd__xor2_1 _08609_ (.A(_02607_),
    .B(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__or2_1 _08610_ (.A(_02606_),
    .B(_02609_),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_1 _08611_ (.A(_02609_),
    .B(_02606_),
    .Y(_02612_));
 sky130_fd_sc_hd__nand2_1 _08612_ (.A(_02611_),
    .B(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21oi_2 _08613_ (.A1(_02503_),
    .A2(_02506_),
    .B1(_02501_),
    .Y(_02614_));
 sky130_fd_sc_hd__inv_2 _08614_ (.A(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _08615_ (.A(_02613_),
    .B(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand3_1 _08616_ (.A(_02611_),
    .B(_02612_),
    .C(_02614_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand3b_1 _08617_ (.A_N(_02604_),
    .B(_02616_),
    .C(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__nand2_1 _08618_ (.A(_02616_),
    .B(_02617_),
    .Y(_02619_));
 sky130_fd_sc_hd__nand2_1 _08619_ (.A(_02619_),
    .B(_02604_),
    .Y(_02620_));
 sky130_fd_sc_hd__nand2_1 _08620_ (.A(_02618_),
    .B(_02620_),
    .Y(_02622_));
 sky130_fd_sc_hd__nand2_1 _08621_ (.A(_02603_),
    .B(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__inv_2 _08622_ (.A(_02622_),
    .Y(_02624_));
 sky130_fd_sc_hd__nand3_2 _08623_ (.A(_02600_),
    .B(_02602_),
    .C(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__nand3_2 _08624_ (.A(_02567_),
    .B(_02623_),
    .C(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand2_1 _08625_ (.A(_02623_),
    .B(_02625_),
    .Y(_02627_));
 sky130_fd_sc_hd__a21boi_1 _08626_ (.A1(_02540_),
    .A2(_02517_),
    .B1_N(_02514_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2_1 _08627_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__nand2_1 _08628_ (.A(_02626_),
    .B(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2_1 _08629_ (.A(_02528_),
    .B(_02529_),
    .Y(_02631_));
 sky130_fd_sc_hd__nor2_1 _08630_ (.A(_02529_),
    .B(_02528_),
    .Y(_02633_));
 sky130_fd_sc_hd__a21oi_2 _08631_ (.A1(_02631_),
    .A2(_02535_),
    .B1(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(_05096_),
    .B(_00520_),
    .Y(_02635_));
 sky130_fd_sc_hd__nor3_1 _08633_ (.A(_02376_),
    .B(_00561_),
    .C(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__o21ai_2 _08634_ (.A1(_02376_),
    .A2(_00561_),
    .B1(_02635_),
    .Y(_02637_));
 sky130_fd_sc_hd__inv_2 _08635_ (.A(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__nand2_1 _08636_ (.A(_02687_),
    .B(_00960_),
    .Y(_02639_));
 sky130_fd_sc_hd__o21ai_1 _08637_ (.A1(_02636_),
    .A2(_02638_),
    .B1(_02639_),
    .Y(_02640_));
 sky130_fd_sc_hd__inv_2 _08638_ (.A(_02639_),
    .Y(_02641_));
 sky130_fd_sc_hd__nand3b_1 _08639_ (.A_N(_02636_),
    .B(_02641_),
    .C(_02637_),
    .Y(_02642_));
 sky130_fd_sc_hd__nand2_1 _08640_ (.A(_02640_),
    .B(_02642_),
    .Y(_02644_));
 sky130_fd_sc_hd__a21oi_1 _08641_ (.A1(_02388_),
    .A2(_02393_),
    .B1(_02387_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand2_1 _08642_ (.A(_02644_),
    .B(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand3b_1 _08643_ (.A_N(_02645_),
    .B(_02640_),
    .C(_02642_),
    .Y(_02647_));
 sky130_fd_sc_hd__nand2_1 _08644_ (.A(_02646_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__nand2_1 _08645_ (.A(_01334_),
    .B(_04645_),
    .Y(_02649_));
 sky130_fd_sc_hd__inv_2 _08646_ (.A(_04128_),
    .Y(_02650_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(_02214_),
    .B(_05114_),
    .Y(_02651_));
 sky130_fd_sc_hd__nor3_1 _08648_ (.A(_01267_),
    .B(_02650_),
    .C(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hd__o21ai_1 _08649_ (.A1(_01267_),
    .A2(_02650_),
    .B1(_02651_),
    .Y(_02653_));
 sky130_fd_sc_hd__inv_2 _08650_ (.A(_02653_),
    .Y(_02655_));
 sky130_fd_sc_hd__nor2_1 _08651_ (.A(_02652_),
    .B(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__xor2_1 _08652_ (.A(_02649_),
    .B(_02656_),
    .X(_02657_));
 sky130_fd_sc_hd__nand2_1 _08653_ (.A(_02648_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__nand3b_1 _08654_ (.A_N(_02657_),
    .B(_02646_),
    .C(_02647_),
    .Y(_02659_));
 sky130_fd_sc_hd__nand3_1 _08655_ (.A(_02634_),
    .B(_02658_),
    .C(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__inv_2 _08656_ (.A(_02634_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand2_1 _08657_ (.A(_02659_),
    .B(_02658_),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_1 _08658_ (.A(_02661_),
    .B(_02662_),
    .Y(_02663_));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_02660_),
    .B(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand2_1 _08660_ (.A(_02398_),
    .B(_02396_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(_02664_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand3b_1 _08662_ (.A_N(_02666_),
    .B(_02660_),
    .C(_02663_),
    .Y(_02668_));
 sky130_fd_sc_hd__nand2_1 _08663_ (.A(_02667_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(_02630_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__inv_2 _08665_ (.A(_02669_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand3_2 _08666_ (.A(_02626_),
    .B(_02671_),
    .C(_02629_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand3_2 _08667_ (.A(_02565_),
    .B(_02670_),
    .C(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand2_1 _08668_ (.A(_02670_),
    .B(_02672_),
    .Y(_02674_));
 sky130_fd_sc_hd__a21boi_1 _08669_ (.A1(_02454_),
    .A2(_02562_),
    .B1_N(_02563_),
    .Y(_02675_));
 sky130_fd_sc_hd__nand2_2 _08670_ (.A(_02674_),
    .B(_02675_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_1 _08671_ (.A(_02673_),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__inv_2 _08672_ (.A(_02489_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_1 _08673_ (.A(_05113_),
    .B(_04899_),
    .Y(_02680_));
 sky130_fd_sc_hd__or3_1 _08674_ (.A(_02679_),
    .B(_00188_),
    .C(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__o21ai_1 _08675_ (.A1(_02679_),
    .A2(_00188_),
    .B1(_02680_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand2_1 _08676_ (.A(_02681_),
    .B(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _08677_ (.A(_05278_),
    .B(_04888_),
    .Y(_02684_));
 sky130_fd_sc_hd__nand2_1 _08678_ (.A(_02683_),
    .B(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__nand3b_2 _08679_ (.A_N(_02684_),
    .B(_02681_),
    .C(_02682_),
    .Y(_02686_));
 sky130_fd_sc_hd__nand2_1 _08680_ (.A(_02685_),
    .B(_02686_),
    .Y(_02688_));
 sky130_fd_sc_hd__nand2_1 _08681_ (.A(_02446_),
    .B(_02439_),
    .Y(_02689_));
 sky130_fd_sc_hd__inv_2 _08682_ (.A(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__nand2_1 _08683_ (.A(_02688_),
    .B(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_00138_),
    .B(_04888_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _08685_ (.A(_05278_),
    .B(_04899_),
    .Y(_02693_));
 sky130_fd_sc_hd__nand2_1 _08686_ (.A(_05113_),
    .B(_04897_),
    .Y(_02694_));
 sky130_fd_sc_hd__or2_1 _08687_ (.A(_02693_),
    .B(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(_02693_),
    .B(_02694_),
    .Y(_02696_));
 sky130_fd_sc_hd__nand2_1 _08689_ (.A(_02695_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__or2_1 _08690_ (.A(_02692_),
    .B(_02697_),
    .X(_02699_));
 sky130_fd_sc_hd__nand2_1 _08691_ (.A(_02699_),
    .B(_02695_),
    .Y(_02700_));
 sky130_fd_sc_hd__nand3_2 _08692_ (.A(_02685_),
    .B(_02686_),
    .C(_02689_),
    .Y(_02701_));
 sky130_fd_sc_hd__a21boi_1 _08693_ (.A1(_02691_),
    .A2(_02700_),
    .B1_N(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__nand2_1 _08694_ (.A(_02686_),
    .B(_02681_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(_05113_),
    .B(_04888_),
    .Y(_02704_));
 sky130_fd_sc_hd__inv_2 _08696_ (.A(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(_03105_),
    .B(_04899_),
    .Y(_02706_));
 sky130_fd_sc_hd__nand2_1 _08698_ (.A(_01532_),
    .B(_04897_),
    .Y(_02707_));
 sky130_fd_sc_hd__xor2_1 _08699_ (.A(_02706_),
    .B(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__or2_1 _08700_ (.A(_02705_),
    .B(_02708_),
    .X(_02710_));
 sky130_fd_sc_hd__nand2_1 _08701_ (.A(_02708_),
    .B(_02705_),
    .Y(_02711_));
 sky130_fd_sc_hd__nand2_1 _08702_ (.A(_02710_),
    .B(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__inv_2 _08703_ (.A(_02367_),
    .Y(_02713_));
 sky130_fd_sc_hd__a21oi_2 _08704_ (.A1(_02372_),
    .A2(_02713_),
    .B1(_02371_),
    .Y(_02714_));
 sky130_fd_sc_hd__inv_2 _08705_ (.A(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand2_1 _08706_ (.A(_02712_),
    .B(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__nand3_1 _08707_ (.A(_02710_),
    .B(_02711_),
    .C(_02714_),
    .Y(_02717_));
 sky130_fd_sc_hd__nand3b_1 _08708_ (.A_N(_02703_),
    .B(_02716_),
    .C(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__nand2_1 _08709_ (.A(_02716_),
    .B(_02717_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_02719_),
    .B(_02703_),
    .Y(_02721_));
 sky130_fd_sc_hd__nand3_1 _08711_ (.A(_02702_),
    .B(_02718_),
    .C(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__nand3_1 _08712_ (.A(_02691_),
    .B(_02701_),
    .C(_02700_),
    .Y(_02723_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(_02723_),
    .B(_02701_),
    .Y(_02724_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(_02718_),
    .B(_02721_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_1 _08715_ (.A(_02724_),
    .B(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__nand2_1 _08716_ (.A(_02722_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__inv_2 _08717_ (.A(_02797_),
    .Y(_02728_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(_00329_),
    .B(_04933_),
    .Y(_02729_));
 sky130_fd_sc_hd__o21ai_2 _08719_ (.A1(_02728_),
    .A2(_05179_),
    .B1(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__nand2_1 _08720_ (.A(_04634_),
    .B(_04941_),
    .Y(_02732_));
 sky130_fd_sc_hd__inv_2 _08721_ (.A(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__nor3_1 _08722_ (.A(_02728_),
    .B(_05179_),
    .C(_02729_),
    .Y(_02734_));
 sky130_fd_sc_hd__a21oi_1 _08723_ (.A1(_02730_),
    .A2(_02733_),
    .B1(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__inv_2 _08724_ (.A(_02555_),
    .Y(_02736_));
 sky130_fd_sc_hd__nand2_1 _08725_ (.A(_02797_),
    .B(_04933_),
    .Y(_02737_));
 sky130_fd_sc_hd__nor3_1 _08726_ (.A(_02736_),
    .B(_05179_),
    .C(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__inv_2 _08727_ (.A(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__o21ai_1 _08728_ (.A1(_02736_),
    .A2(_05179_),
    .B1(_02737_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand2_1 _08729_ (.A(_00329_),
    .B(_04941_),
    .Y(_02741_));
 sky130_fd_sc_hd__a21bo_1 _08730_ (.A1(_02739_),
    .A2(_02740_),
    .B1_N(_02741_),
    .X(_02743_));
 sky130_fd_sc_hd__nand3b_1 _08731_ (.A_N(_02741_),
    .B(_02739_),
    .C(_02740_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand2_1 _08732_ (.A(_02743_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__nor2_1 _08733_ (.A(_02735_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__nand2_1 _08734_ (.A(_02745_),
    .B(_02735_),
    .Y(_02747_));
 sky130_fd_sc_hd__inv_2 _08735_ (.A(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__nand2_1 _08736_ (.A(_00682_),
    .B(_04880_),
    .Y(_02749_));
 sky130_fd_sc_hd__inv_2 _08737_ (.A(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__inv_2 _08738_ (.A(net46),
    .Y(_02751_));
 sky130_fd_sc_hd__inv_2 _08739_ (.A(_04634_),
    .Y(_02752_));
 sky130_fd_sc_hd__nand2_1 _08740_ (.A(_05191_),
    .B(_04814_),
    .Y(_02754_));
 sky130_fd_sc_hd__nor3_1 _08741_ (.A(_02751_),
    .B(_02752_),
    .C(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__o21ai_1 _08742_ (.A1(_02751_),
    .A2(_02752_),
    .B1(_02754_),
    .Y(_02756_));
 sky130_fd_sc_hd__nor2b_1 _08743_ (.A(_02755_),
    .B_N(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__or2_1 _08744_ (.A(_02750_),
    .B(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(_02757_),
    .B(_02750_),
    .Y(_02759_));
 sky130_fd_sc_hd__nand2_1 _08746_ (.A(_02758_),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__o21ai_1 _08747_ (.A1(_02746_),
    .A2(_02748_),
    .B1(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__inv_2 _08748_ (.A(_02746_),
    .Y(_02762_));
 sky130_fd_sc_hd__inv_2 _08749_ (.A(_02760_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand3_1 _08750_ (.A(_02762_),
    .B(_02763_),
    .C(_02747_),
    .Y(_02765_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(_02761_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__inv_2 _08752_ (.A(_02766_),
    .Y(_02767_));
 sky130_fd_sc_hd__nand2_1 _08753_ (.A(_02727_),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand3_1 _08754_ (.A(_02722_),
    .B(_02766_),
    .C(_02726_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2_1 _08755_ (.A(_02768_),
    .B(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _08756_ (.A(_02404_),
    .B(_02420_),
    .Y(_02771_));
 sky130_fd_sc_hd__nor2_1 _08757_ (.A(_02420_),
    .B(_02404_),
    .Y(_02772_));
 sky130_fd_sc_hd__a21oi_2 _08758_ (.A1(_02771_),
    .A2(_02450_),
    .B1(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__inv_2 _08759_ (.A(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_02770_),
    .B(_02774_),
    .Y(_02776_));
 sky130_fd_sc_hd__nand3_1 _08761_ (.A(_02773_),
    .B(_02768_),
    .C(_02769_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _08762_ (.A(_02776_),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand2_1 _08763_ (.A(_02691_),
    .B(_02701_),
    .Y(_02779_));
 sky130_fd_sc_hd__inv_2 _08764_ (.A(_02700_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2_1 _08765_ (.A(_02779_),
    .B(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(_02781_),
    .B(_02723_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2_1 _08767_ (.A(_02697_),
    .B(_02692_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand2_1 _08768_ (.A(_02699_),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__nand2_1 _08769_ (.A(_00599_),
    .B(_00593_),
    .Y(_02785_));
 sky130_fd_sc_hd__inv_2 _08770_ (.A(_02785_),
    .Y(_02787_));
 sky130_fd_sc_hd__nand2_1 _08771_ (.A(_02784_),
    .B(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _08772_ (.A(_00657_),
    .B(_00651_),
    .Y(_02789_));
 sky130_fd_sc_hd__nor2_1 _08773_ (.A(_02787_),
    .B(_02784_),
    .Y(_02790_));
 sky130_fd_sc_hd__a21oi_2 _08774_ (.A1(_02788_),
    .A2(_02789_),
    .B1(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__inv_2 _08775_ (.A(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__nand2_1 _08776_ (.A(_02782_),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand3_1 _08777_ (.A(_02781_),
    .B(_02791_),
    .C(_02723_),
    .Y(_02794_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(_02793_),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__inv_2 _08779_ (.A(_02730_),
    .Y(_02796_));
 sky130_fd_sc_hd__o21ai_1 _08780_ (.A1(_02734_),
    .A2(_02796_),
    .B1(_02732_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand3b_1 _08781_ (.A_N(_02734_),
    .B(_02733_),
    .C(_02730_),
    .Y(_02799_));
 sky130_fd_sc_hd__nand2_1 _08782_ (.A(_02798_),
    .B(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__nand2_1 _08783_ (.A(_00893_),
    .B(_04941_),
    .Y(_02801_));
 sky130_fd_sc_hd__inv_2 _08784_ (.A(_00329_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _08785_ (.A(_05159_),
    .B(_04933_),
    .Y(_02803_));
 sky130_fd_sc_hd__nor3_1 _08786_ (.A(_02802_),
    .B(_05179_),
    .C(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__inv_2 _08787_ (.A(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__o21ai_1 _08788_ (.A1(_02802_),
    .A2(_05179_),
    .B1(_02803_),
    .Y(_02806_));
 sky130_fd_sc_hd__nand3b_1 _08789_ (.A_N(_02801_),
    .B(_02805_),
    .C(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _08790_ (.A(_02807_),
    .B(_02805_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2b_1 _08791_ (.A_N(_02800_),
    .B(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__nand2b_1 _08792_ (.A_N(_02809_),
    .B(_02800_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand2_1 _08793_ (.A(_00682_),
    .B(_00381_),
    .Y(_02812_));
 sky130_fd_sc_hd__nand2_1 _08794_ (.A(_05191_),
    .B(_00384_),
    .Y(_02813_));
 sky130_fd_sc_hd__nor3_1 _08795_ (.A(_02751_),
    .B(_05178_),
    .C(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__o21ai_1 _08796_ (.A1(_02751_),
    .A2(_05178_),
    .B1(_02813_),
    .Y(_02815_));
 sky130_fd_sc_hd__inv_2 _08797_ (.A(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__nor2_1 _08798_ (.A(_02814_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__xor2_1 _08799_ (.A(_02812_),
    .B(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__inv_2 _08800_ (.A(_02818_),
    .Y(_02820_));
 sky130_fd_sc_hd__a21o_1 _08801_ (.A1(_02810_),
    .A2(_02811_),
    .B1(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__nand3_1 _08802_ (.A(_02810_),
    .B(_02811_),
    .C(_02820_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _08803_ (.A(_02821_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__inv_2 _08804_ (.A(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_02795_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__or2_1 _08806_ (.A(_02791_),
    .B(_02782_),
    .X(_02826_));
 sky130_fd_sc_hd__nand2_1 _08807_ (.A(_02825_),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__nand2_1 _08808_ (.A(_02778_),
    .B(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__nand3b_1 _08809_ (.A_N(_02827_),
    .B(_02776_),
    .C(_02777_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _08810_ (.A(_02828_),
    .B(_02829_),
    .Y(_02831_));
 sky130_fd_sc_hd__nand2_1 _08811_ (.A(_02678_),
    .B(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__inv_2 _08812_ (.A(_02831_),
    .Y(_02833_));
 sky130_fd_sc_hd__nand3_2 _08813_ (.A(_02673_),
    .B(_02833_),
    .C(_02677_),
    .Y(_02834_));
 sky130_fd_sc_hd__nand2_1 _08814_ (.A(_02832_),
    .B(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__nand3_1 _08815_ (.A(_02823_),
    .B(_02793_),
    .C(_02794_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand2_1 _08816_ (.A(_02825_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__nand3_1 _08817_ (.A(_02447_),
    .B(_02433_),
    .C(_02435_),
    .Y(_02838_));
 sky130_fd_sc_hd__nand2_1 _08818_ (.A(_02449_),
    .B(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__nand2_1 _08819_ (.A(_00579_),
    .B(_00573_),
    .Y(_02840_));
 sky130_fd_sc_hd__inv_2 _08820_ (.A(_02840_),
    .Y(_02842_));
 sky130_fd_sc_hd__nand2_1 _08821_ (.A(_02839_),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__nand2_1 _08822_ (.A(_00617_),
    .B(_00616_),
    .Y(_02844_));
 sky130_fd_sc_hd__nor2_1 _08823_ (.A(_02842_),
    .B(_02839_),
    .Y(_02845_));
 sky130_fd_sc_hd__a21oi_2 _08824_ (.A1(_02843_),
    .A2(_02844_),
    .B1(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__inv_2 _08825_ (.A(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__nand2_1 _08826_ (.A(_02837_),
    .B(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hd__nand3_1 _08827_ (.A(_02846_),
    .B(_02825_),
    .C(_02836_),
    .Y(_02849_));
 sky130_fd_sc_hd__nand2_1 _08828_ (.A(_02848_),
    .B(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__nand2_1 _08829_ (.A(_00658_),
    .B(_00659_),
    .Y(_02851_));
 sky130_fd_sc_hd__nor2_1 _08830_ (.A(_00659_),
    .B(_00658_),
    .Y(_02853_));
 sky130_fd_sc_hd__a21oi_1 _08831_ (.A1(_02851_),
    .A2(_00665_),
    .B1(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__nand2_1 _08832_ (.A(_02784_),
    .B(_02785_),
    .Y(_02855_));
 sky130_fd_sc_hd__nand3_1 _08833_ (.A(_02787_),
    .B(_02699_),
    .C(_02783_),
    .Y(_02856_));
 sky130_fd_sc_hd__nand2_1 _08834_ (.A(_02855_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(_02857_),
    .B(_02789_),
    .Y(_02858_));
 sky130_fd_sc_hd__nand3b_1 _08836_ (.A_N(_02789_),
    .B(_02855_),
    .C(_02856_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_1 _08837_ (.A(_02858_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__inv_2 _08838_ (.A(_02854_),
    .Y(_02861_));
 sky130_fd_sc_hd__nand2_1 _08839_ (.A(_02860_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__nand3_1 _08840_ (.A(_02858_),
    .B(_02859_),
    .C(_02854_),
    .Y(_02864_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(_02862_),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(_00694_),
    .B(_00691_),
    .Y(_02866_));
 sky130_fd_sc_hd__inv_2 _08843_ (.A(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__a21bo_1 _08844_ (.A1(_02805_),
    .A2(_02806_),
    .B1_N(_02801_),
    .X(_02868_));
 sky130_fd_sc_hd__nand3_1 _08845_ (.A(_02867_),
    .B(_02868_),
    .C(_02807_),
    .Y(_02869_));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(_02868_),
    .B(_02807_),
    .Y(_02870_));
 sky130_fd_sc_hd__nand2_1 _08847_ (.A(_02870_),
    .B(_02866_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_1 _08848_ (.A(_02869_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(_00682_),
    .B(_05310_),
    .Y(_02873_));
 sky130_fd_sc_hd__inv_2 _08850_ (.A(_04880_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _08851_ (.A(_05191_),
    .B(_00381_),
    .Y(_02876_));
 sky130_fd_sc_hd__nor3_1 _08852_ (.A(_02751_),
    .B(_02875_),
    .C(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__o21ai_1 _08853_ (.A1(_02751_),
    .A2(_02875_),
    .B1(_02876_),
    .Y(_02878_));
 sky130_fd_sc_hd__inv_2 _08854_ (.A(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__nor2_1 _08855_ (.A(_02877_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__xor2_1 _08856_ (.A(_02873_),
    .B(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__inv_2 _08857_ (.A(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__nand2_1 _08858_ (.A(_02872_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand3_1 _08859_ (.A(_02869_),
    .B(_02881_),
    .C(_02871_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _08860_ (.A(_02883_),
    .B(_02884_),
    .Y(_02886_));
 sky130_fd_sc_hd__inv_2 _08861_ (.A(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__nand2_1 _08862_ (.A(_02865_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__o21ai_1 _08863_ (.A1(_02854_),
    .A2(_02860_),
    .B1(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__nand2_1 _08864_ (.A(_02850_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__nand3b_1 _08865_ (.A_N(_02889_),
    .B(_02848_),
    .C(_02849_),
    .Y(_02891_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_02890_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__inv_2 _08867_ (.A(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(_02562_),
    .B(_02563_),
    .Y(_02894_));
 sky130_fd_sc_hd__nand2_1 _08869_ (.A(_02894_),
    .B(_02453_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_02895_),
    .B(_02564_),
    .Y(_02897_));
 sky130_fd_sc_hd__nand2_1 _08871_ (.A(_02839_),
    .B(_02840_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand3_1 _08872_ (.A(_02449_),
    .B(_02838_),
    .C(_02842_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _08873_ (.A(_02898_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(_02900_),
    .B(_02844_),
    .Y(_02901_));
 sky130_fd_sc_hd__nand3b_1 _08875_ (.A_N(_02844_),
    .B(_02898_),
    .C(_02899_),
    .Y(_02902_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__inv_2 _08877_ (.A(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2_1 _08878_ (.A(_02549_),
    .B(_02558_),
    .Y(_02905_));
 sky130_fd_sc_hd__nand2_1 _08879_ (.A(_02905_),
    .B(_02556_),
    .Y(_02906_));
 sky130_fd_sc_hd__nand2_1 _08880_ (.A(_02906_),
    .B(_02559_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand2_1 _08881_ (.A(_00582_),
    .B(_00555_),
    .Y(_02909_));
 sky130_fd_sc_hd__inv_2 _08882_ (.A(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__nand2_2 _08883_ (.A(_02908_),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__nand3_2 _08884_ (.A(_02906_),
    .B(_02909_),
    .C(_02559_),
    .Y(_02912_));
 sky130_fd_sc_hd__a21boi_2 _08885_ (.A1(_02904_),
    .A2(_02911_),
    .B1_N(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(_02897_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__nor2_1 _08887_ (.A(_02913_),
    .B(_02897_),
    .Y(_02915_));
 sky130_fd_sc_hd__a21oi_2 _08888_ (.A1(_02893_),
    .A2(_02914_),
    .B1(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__inv_2 _08889_ (.A(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__nand2_1 _08890_ (.A(_02835_),
    .B(_02917_),
    .Y(_02919_));
 sky130_fd_sc_hd__nand3_1 _08891_ (.A(_02916_),
    .B(_02832_),
    .C(_02834_),
    .Y(_02920_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__nand2_1 _08893_ (.A(_02837_),
    .B(_02846_),
    .Y(_02922_));
 sky130_fd_sc_hd__nor2_1 _08894_ (.A(_02846_),
    .B(_02837_),
    .Y(_02923_));
 sky130_fd_sc_hd__a21oi_1 _08895_ (.A1(_02922_),
    .A2(_02889_),
    .B1(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__inv_2 _08896_ (.A(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_1 _08897_ (.A(net51),
    .B(_04958_),
    .Y(_02926_));
 sky130_fd_sc_hd__inv_2 _08898_ (.A(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__nand2_1 _08899_ (.A(net50),
    .B(_05310_),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_1 _08900_ (.A(net49),
    .B(_00381_),
    .Y(_02930_));
 sky130_fd_sc_hd__xor2_1 _08901_ (.A(_02928_),
    .B(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__or2_1 _08902_ (.A(_02927_),
    .B(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_1 _08903_ (.A(_02931_),
    .B(_02927_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _08904_ (.A(_02932_),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__inv_2 _08905_ (.A(_02812_),
    .Y(_02935_));
 sky130_fd_sc_hd__a21oi_1 _08906_ (.A1(_02815_),
    .A2(_02935_),
    .B1(_02814_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand2_1 _08907_ (.A(_02934_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand3b_1 _08908_ (.A_N(_02936_),
    .B(_02932_),
    .C(_02933_),
    .Y(_02938_));
 sky130_fd_sc_hd__nand2_1 _08909_ (.A(_02937_),
    .B(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__and4_1 _08910_ (.A(net49),
    .B(net50),
    .C(_04947_),
    .D(net1),
    .X(_02941_));
 sky130_fd_sc_hd__inv_2 _08911_ (.A(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2_1 _08912_ (.A(_02939_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand3_1 _08913_ (.A(_02937_),
    .B(_02938_),
    .C(_02941_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_1 _08914_ (.A(_02943_),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__a21boi_1 _08915_ (.A1(_02811_),
    .A2(_02820_),
    .B1_N(_02810_),
    .Y(_02946_));
 sky130_fd_sc_hd__nor2_1 _08916_ (.A(_02945_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__nand2_1 _08917_ (.A(_02946_),
    .B(_02945_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2b_1 _08918_ (.A_N(_02947_),
    .B(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__a22o_1 _08919_ (.A1(net49),
    .A2(_05310_),
    .B1(net50),
    .B2(_04958_),
    .X(_02950_));
 sky130_fd_sc_hd__nand2_1 _08920_ (.A(_02942_),
    .B(_02950_),
    .Y(_02952_));
 sky130_fd_sc_hd__o21ba_1 _08921_ (.A1(_02873_),
    .A2(_02879_),
    .B1_N(_02877_),
    .X(_02953_));
 sky130_fd_sc_hd__nor2_1 _08922_ (.A(_02952_),
    .B(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__inv_2 _08923_ (.A(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__nand2_1 _08924_ (.A(_02949_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__nand3b_1 _08925_ (.A_N(_02947_),
    .B(_02954_),
    .C(_02948_),
    .Y(_02957_));
 sky130_fd_sc_hd__nand2_1 _08926_ (.A(_02956_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand2_1 _08927_ (.A(_02953_),
    .B(_02952_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand2_1 _08928_ (.A(_02955_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__nand2_1 _08929_ (.A(_02870_),
    .B(_02867_),
    .Y(_02961_));
 sky130_fd_sc_hd__nor2_1 _08930_ (.A(_02867_),
    .B(_02870_),
    .Y(_02963_));
 sky130_fd_sc_hd__a21oi_1 _08931_ (.A1(_02961_),
    .A2(_02882_),
    .B1(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__nor2_1 _08932_ (.A(_02960_),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__inv_2 _08933_ (.A(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__nand2_1 _08934_ (.A(net49),
    .B(_00194_),
    .Y(_02967_));
 sky130_fd_sc_hd__and2_1 _08935_ (.A(_00683_),
    .B(_00679_),
    .X(_02968_));
 sky130_fd_sc_hd__nor2_1 _08936_ (.A(_02967_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2_1 _08937_ (.A(_02964_),
    .B(_02960_),
    .Y(_02970_));
 sky130_fd_sc_hd__nand3_1 _08938_ (.A(_02966_),
    .B(_02969_),
    .C(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__nand2_1 _08939_ (.A(_02971_),
    .B(_02966_),
    .Y(_02972_));
 sky130_fd_sc_hd__inv_2 _08940_ (.A(_02972_),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_1 _08941_ (.A(_02958_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__nand3_1 _08942_ (.A(_02956_),
    .B(_02972_),
    .C(_02957_),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(_02975_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__inv_2 _08944_ (.A(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__nand2_1 _08945_ (.A(_02925_),
    .B(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__nand2_1 _08946_ (.A(_02924_),
    .B(_02977_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand2_1 _08947_ (.A(_02979_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__a21o_1 _08948_ (.A1(_02966_),
    .A2(_02970_),
    .B1(_02969_),
    .X(_02982_));
 sky130_fd_sc_hd__nand2_1 _08949_ (.A(_02968_),
    .B(_02967_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2b_1 _08950_ (.A_N(_02969_),
    .B(_02983_),
    .Y(_02985_));
 sky130_fd_sc_hd__and2_1 _08951_ (.A(_00702_),
    .B(_00698_),
    .X(_02986_));
 sky130_fd_sc_hd__nor2_1 _08952_ (.A(_02985_),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__nand3_1 _08953_ (.A(_02982_),
    .B(_02971_),
    .C(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__nand2_1 _08954_ (.A(_02981_),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand3b_1 _08955_ (.A_N(_02988_),
    .B(_02979_),
    .C(_02980_),
    .Y(_02990_));
 sky130_fd_sc_hd__nand2_1 _08956_ (.A(_02989_),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__inv_2 _08957_ (.A(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__nand2_1 _08958_ (.A(_02921_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__nand3_1 _08959_ (.A(_02919_),
    .B(_02920_),
    .C(_02991_),
    .Y(_02994_));
 sky130_fd_sc_hd__nand2_1 _08960_ (.A(_02993_),
    .B(_02994_),
    .Y(_02996_));
 sky130_fd_sc_hd__nand3_1 _08961_ (.A(_02904_),
    .B(_02912_),
    .C(_02911_),
    .Y(_02997_));
 sky130_fd_sc_hd__nand2_1 _08962_ (.A(_02997_),
    .B(_02912_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand2_1 _08963_ (.A(_02897_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__nand3_1 _08964_ (.A(_02913_),
    .B(_02895_),
    .C(_02564_),
    .Y(_03000_));
 sky130_fd_sc_hd__nand2_1 _08965_ (.A(_02999_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__nand2_1 _08966_ (.A(_03001_),
    .B(_02893_),
    .Y(_03002_));
 sky130_fd_sc_hd__nand3_1 _08967_ (.A(_02999_),
    .B(_03000_),
    .C(_02892_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(_03002_),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_02911_),
    .B(_02912_),
    .Y(_03005_));
 sky130_fd_sc_hd__nand2_1 _08970_ (.A(_03005_),
    .B(_02903_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _08971_ (.A(_02997_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__nand2_2 _08972_ (.A(_00636_),
    .B(_00587_),
    .Y(_03009_));
 sky130_fd_sc_hd__inv_2 _08973_ (.A(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(_03008_),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__or2_1 _08975_ (.A(_00625_),
    .B(_00622_),
    .X(_03012_));
 sky130_fd_sc_hd__nand2_1 _08976_ (.A(_00632_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__inv_2 _08977_ (.A(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand3_1 _08978_ (.A(_02886_),
    .B(_02862_),
    .C(_02864_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand3_1 _08979_ (.A(_03014_),
    .B(_02888_),
    .C(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__nand2_1 _08980_ (.A(_02888_),
    .B(_03015_),
    .Y(_03018_));
 sky130_fd_sc_hd__nand2_1 _08981_ (.A(_03018_),
    .B(_03013_),
    .Y(_03019_));
 sky130_fd_sc_hd__nand2_1 _08982_ (.A(_03016_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__nor2_1 _08983_ (.A(_00671_),
    .B(_00668_),
    .Y(_03021_));
 sky130_fd_sc_hd__inv_2 _08984_ (.A(_00708_),
    .Y(_03022_));
 sky130_fd_sc_hd__nor2_1 _08985_ (.A(_03021_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__inv_2 _08986_ (.A(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__nand2_1 _08987_ (.A(_03020_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nand3_1 _08988_ (.A(_03016_),
    .B(_03019_),
    .C(_03023_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand2_1 _08989_ (.A(_03025_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__inv_2 _08990_ (.A(_03027_),
    .Y(_03029_));
 sky130_fd_sc_hd__nor2_1 _08991_ (.A(_03010_),
    .B(_03008_),
    .Y(_03030_));
 sky130_fd_sc_hd__a21oi_2 _08992_ (.A1(_03011_),
    .A2(_03029_),
    .B1(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__nand2_1 _08993_ (.A(_03004_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__nand2_1 _08994_ (.A(_03018_),
    .B(_03014_),
    .Y(_03033_));
 sky130_fd_sc_hd__nor2_1 _08995_ (.A(_03014_),
    .B(_03018_),
    .Y(_03034_));
 sky130_fd_sc_hd__a21oi_1 _08996_ (.A1(_03033_),
    .A2(_03024_),
    .B1(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__inv_2 _08997_ (.A(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__nand2_1 _08998_ (.A(_02982_),
    .B(_02971_),
    .Y(_03037_));
 sky130_fd_sc_hd__inv_2 _08999_ (.A(_02987_),
    .Y(_03038_));
 sky130_fd_sc_hd__nand2_1 _09000_ (.A(_03037_),
    .B(_03038_),
    .Y(_03040_));
 sky130_fd_sc_hd__nand3_1 _09001_ (.A(_03036_),
    .B(_02988_),
    .C(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__nand2_1 _09002_ (.A(_03040_),
    .B(_02988_),
    .Y(_03042_));
 sky130_fd_sc_hd__nand2_1 _09003_ (.A(_03042_),
    .B(_03035_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand2_1 _09004_ (.A(_03041_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__nand2_1 _09005_ (.A(_02986_),
    .B(_02985_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(_03038_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__or2_1 _09007_ (.A(_00739_),
    .B(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__nand2_1 _09008_ (.A(_03044_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__nand3b_1 _09009_ (.A_N(_03047_),
    .B(_03041_),
    .C(_03043_),
    .Y(_03049_));
 sky130_fd_sc_hd__nand2_1 _09010_ (.A(_03048_),
    .B(_03049_),
    .Y(_03051_));
 sky130_fd_sc_hd__inv_2 _09011_ (.A(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__nor2_1 _09012_ (.A(_03031_),
    .B(_03004_),
    .Y(_03053_));
 sky130_fd_sc_hd__a21oi_2 _09013_ (.A1(_03032_),
    .A2(_03052_),
    .B1(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__inv_2 _09014_ (.A(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_02996_),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__nand3_1 _09016_ (.A(_03054_),
    .B(_02993_),
    .C(_02994_),
    .Y(_03057_));
 sky130_fd_sc_hd__nand2_1 _09017_ (.A(_03056_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand2_1 _09018_ (.A(_03049_),
    .B(_03041_),
    .Y(_03059_));
 sky130_fd_sc_hd__inv_2 _09019_ (.A(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__nand2_1 _09020_ (.A(_03058_),
    .B(_03060_),
    .Y(_03062_));
 sky130_fd_sc_hd__nand3_1 _09021_ (.A(_03056_),
    .B(_03057_),
    .C(_03059_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand2_1 _09022_ (.A(_03062_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__inv_2 _09023_ (.A(_03031_),
    .Y(_03065_));
 sky130_fd_sc_hd__nand2_1 _09024_ (.A(_03004_),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__nand3_1 _09025_ (.A(_03031_),
    .B(_03002_),
    .C(_03003_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _09026_ (.A(_03066_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__nand2_1 _09027_ (.A(_03068_),
    .B(_03052_),
    .Y(_03069_));
 sky130_fd_sc_hd__nand3_1 _09028_ (.A(_03066_),
    .B(_03067_),
    .C(_03051_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand2_1 _09029_ (.A(_03069_),
    .B(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__nand2_1 _09030_ (.A(_03008_),
    .B(_03009_),
    .Y(_03073_));
 sky130_fd_sc_hd__nand3_1 _09031_ (.A(_03010_),
    .B(_02997_),
    .C(_03007_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _09032_ (.A(_03073_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2_1 _09033_ (.A(_03075_),
    .B(_03029_),
    .Y(_03076_));
 sky130_fd_sc_hd__nand3_1 _09034_ (.A(_03073_),
    .B(_03074_),
    .C(_03027_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand2_1 _09035_ (.A(_03076_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__nand3_1 _09036_ (.A(_00644_),
    .B(_00636_),
    .C(_00639_),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_1 _09037_ (.A(_00727_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__inv_2 _09038_ (.A(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__nand2_1 _09039_ (.A(_03078_),
    .B(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__nand2_1 _09040_ (.A(_03046_),
    .B(_00739_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2_1 _09041_ (.A(_03047_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__o21a_1 _09042_ (.A1(_00710_),
    .A2(_00713_),
    .B1(_00723_),
    .X(_03086_));
 sky130_fd_sc_hd__nor2_1 _09043_ (.A(_03085_),
    .B(_03086_),
    .Y(_03087_));
 sky130_fd_sc_hd__nand2_1 _09044_ (.A(_03086_),
    .B(_03085_),
    .Y(_03088_));
 sky130_fd_sc_hd__nor2b_1 _09045_ (.A(_03087_),
    .B_N(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__nor2_1 _09046_ (.A(_03081_),
    .B(_03078_),
    .Y(_03090_));
 sky130_fd_sc_hd__a21oi_2 _09047_ (.A1(_03082_),
    .A2(_03089_),
    .B1(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__nand2_1 _09048_ (.A(_03071_),
    .B(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__nor2_1 _09049_ (.A(_03091_),
    .B(_03071_),
    .Y(_03093_));
 sky130_fd_sc_hd__a21oi_1 _09050_ (.A1(_03092_),
    .A2(_03087_),
    .B1(_03093_),
    .Y(_03095_));
 sky130_fd_sc_hd__inv_2 _09051_ (.A(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_2 _09052_ (.A(_03064_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__nand3_1 _09053_ (.A(_03095_),
    .B(_03062_),
    .C(_03063_),
    .Y(_03098_));
 sky130_fd_sc_hd__nand2_1 _09054_ (.A(_03097_),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__nand2_1 _09055_ (.A(_03078_),
    .B(_03080_),
    .Y(_03100_));
 sky130_fd_sc_hd__nand3_1 _09056_ (.A(_03081_),
    .B(_03076_),
    .C(_03077_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _09057_ (.A(_03100_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__nand2_1 _09058_ (.A(_03102_),
    .B(_03089_),
    .Y(_03103_));
 sky130_fd_sc_hd__nand3b_1 _09059_ (.A_N(_03089_),
    .B(_03100_),
    .C(_03101_),
    .Y(_03104_));
 sky130_fd_sc_hd__nand2_1 _09060_ (.A(_03103_),
    .B(_03104_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2_1 _09061_ (.A(_00730_),
    .B(_00733_),
    .Y(_03107_));
 sky130_fd_sc_hd__nor2_1 _09062_ (.A(_00733_),
    .B(_00730_),
    .Y(_03108_));
 sky130_fd_sc_hd__a21oi_2 _09063_ (.A1(_03107_),
    .A2(_00748_),
    .B1(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__nand2_1 _09064_ (.A(_03106_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__nor2_1 _09065_ (.A(_03109_),
    .B(_03106_),
    .Y(_03111_));
 sky130_fd_sc_hd__a21oi_2 _09066_ (.A1(_03110_),
    .A2(_00744_),
    .B1(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__inv_2 _09067_ (.A(_03091_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _09068_ (.A(_03071_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__nand3_1 _09069_ (.A(_03069_),
    .B(_03091_),
    .C(_03070_),
    .Y(_03115_));
 sky130_fd_sc_hd__nand2_1 _09070_ (.A(_03114_),
    .B(_03115_),
    .Y(_03117_));
 sky130_fd_sc_hd__nand2_1 _09071_ (.A(_03117_),
    .B(_03087_),
    .Y(_03118_));
 sky130_fd_sc_hd__nand3b_1 _09072_ (.A_N(_03087_),
    .B(_03114_),
    .C(_03115_),
    .Y(_03119_));
 sky130_fd_sc_hd__nand2_1 _09073_ (.A(_03118_),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__nor2_1 _09074_ (.A(_03112_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__inv_2 _09075_ (.A(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_1 _09076_ (.A(_03099_),
    .B(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__nand3_2 _09077_ (.A(_03097_),
    .B(_03121_),
    .C(_03098_),
    .Y(_03124_));
 sky130_fd_sc_hd__nand2_1 _09078_ (.A(_03123_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__inv_2 _09079_ (.A(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(_02990_),
    .B(_02979_),
    .Y(_03128_));
 sky130_fd_sc_hd__nand2_1 _09081_ (.A(_02835_),
    .B(_02916_),
    .Y(_03129_));
 sky130_fd_sc_hd__nor2_1 _09082_ (.A(_02916_),
    .B(_02835_),
    .Y(_03130_));
 sky130_fd_sc_hd__a21o_1 _09083_ (.A1(_03129_),
    .A2(_02992_),
    .B1(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__nand2_1 _09084_ (.A(_02770_),
    .B(_02773_),
    .Y(_03132_));
 sky130_fd_sc_hd__nor2_1 _09085_ (.A(_02773_),
    .B(_02770_),
    .Y(_03133_));
 sky130_fd_sc_hd__a21o_1 _09086_ (.A1(_03132_),
    .A2(_02827_),
    .B1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__inv_2 _09087_ (.A(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__a21oi_1 _09088_ (.A1(_02763_),
    .A2(_02747_),
    .B1(_02746_),
    .Y(_03136_));
 sky130_fd_sc_hd__inv_2 _09089_ (.A(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__nand2_1 _09090_ (.A(net51),
    .B(_05310_),
    .Y(_03139_));
 sky130_fd_sc_hd__inv_2 _09091_ (.A(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__nand2_1 _09092_ (.A(net50),
    .B(_00381_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand2_1 _09093_ (.A(net49),
    .B(_00384_),
    .Y(_03142_));
 sky130_fd_sc_hd__xor2_1 _09094_ (.A(_03141_),
    .B(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__or2_1 _09095_ (.A(_03140_),
    .B(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_03143_),
    .B(_03140_),
    .Y(_03145_));
 sky130_fd_sc_hd__a21oi_2 _09097_ (.A1(_02756_),
    .A2(_02750_),
    .B1(_02755_),
    .Y(_03146_));
 sky130_fd_sc_hd__a21o_1 _09098_ (.A1(_03144_),
    .A2(_03145_),
    .B1(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__inv_2 _09099_ (.A(net49),
    .Y(_03148_));
 sky130_fd_sc_hd__nor3_1 _09100_ (.A(_03148_),
    .B(_02309_),
    .C(_02928_),
    .Y(_03150_));
 sky130_fd_sc_hd__inv_2 _09101_ (.A(_02933_),
    .Y(_03151_));
 sky130_fd_sc_hd__nor2_1 _09102_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__nand3_1 _09103_ (.A(_03144_),
    .B(_03145_),
    .C(_03146_),
    .Y(_03153_));
 sky130_fd_sc_hd__nand3_1 _09104_ (.A(_03147_),
    .B(_03152_),
    .C(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__nand2_1 _09105_ (.A(_03147_),
    .B(_03153_),
    .Y(_03155_));
 sky130_fd_sc_hd__o21ai_2 _09106_ (.A1(_03150_),
    .A2(_03151_),
    .B1(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__nand3_2 _09107_ (.A(_03137_),
    .B(_03154_),
    .C(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__nand2_1 _09108_ (.A(_03156_),
    .B(_03154_),
    .Y(_03158_));
 sky130_fd_sc_hd__nand2_1 _09109_ (.A(_03158_),
    .B(_03136_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_1 _09110_ (.A(_03157_),
    .B(_03159_),
    .Y(_03161_));
 sky130_fd_sc_hd__nand2_1 _09111_ (.A(_02944_),
    .B(_02938_),
    .Y(_03162_));
 sky130_fd_sc_hd__inv_2 _09112_ (.A(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__nand2_1 _09113_ (.A(_03161_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__nand3_2 _09114_ (.A(_03157_),
    .B(_03159_),
    .C(_03162_),
    .Y(_03165_));
 sky130_fd_sc_hd__nand2_1 _09115_ (.A(_03164_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__a21oi_1 _09116_ (.A1(_02948_),
    .A2(_02954_),
    .B1(_02947_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand2_1 _09117_ (.A(_03166_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__inv_2 _09118_ (.A(_03167_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand3_2 _09119_ (.A(_03169_),
    .B(_03164_),
    .C(_03165_),
    .Y(_03170_));
 sky130_fd_sc_hd__nand2_1 _09120_ (.A(_03168_),
    .B(_03170_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand2_1 _09121_ (.A(net52),
    .B(_00194_),
    .Y(_03173_));
 sky130_fd_sc_hd__nand2_1 _09122_ (.A(_03172_),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand3b_2 _09123_ (.A_N(_03173_),
    .B(_03168_),
    .C(_03170_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand2_1 _09124_ (.A(_03174_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand2_1 _09125_ (.A(_03135_),
    .B(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__nand3_2 _09126_ (.A(_03134_),
    .B(_03174_),
    .C(_03175_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_1 _09127_ (.A(_03177_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(_03179_),
    .B(_02976_),
    .Y(_03180_));
 sky130_fd_sc_hd__inv_2 _09129_ (.A(_02976_),
    .Y(_03181_));
 sky130_fd_sc_hd__nand3_1 _09130_ (.A(_03177_),
    .B(_03178_),
    .C(_03181_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2_1 _09131_ (.A(_03180_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__inv_2 _09132_ (.A(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_1 _09133_ (.A(_02834_),
    .B(_02673_),
    .Y(_03186_));
 sky130_fd_sc_hd__nand2_1 _09134_ (.A(_02672_),
    .B(_02626_),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_1 _09135_ (.A(_02575_),
    .B(_02572_),
    .Y(_03188_));
 sky130_fd_sc_hd__nand2_1 _09136_ (.A(_00433_),
    .B(net19),
    .Y(_03189_));
 sky130_fd_sc_hd__inv_2 _09137_ (.A(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(_00232_),
    .B(net18),
    .Y(_03191_));
 sky130_fd_sc_hd__nand2_1 _09139_ (.A(_00234_),
    .B(net17),
    .Y(_03192_));
 sky130_fd_sc_hd__xor2_1 _09140_ (.A(_03191_),
    .B(_03192_),
    .X(_03194_));
 sky130_fd_sc_hd__or2_1 _09141_ (.A(_03190_),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__nand2_1 _09142_ (.A(_03194_),
    .B(_03190_),
    .Y(_03196_));
 sky130_fd_sc_hd__nand2_1 _09143_ (.A(_03195_),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__nand2b_1 _09144_ (.A_N(_03188_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__nand3_1 _09145_ (.A(_03188_),
    .B(_03195_),
    .C(_03196_),
    .Y(_03199_));
 sky130_fd_sc_hd__nand2_1 _09146_ (.A(_03198_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _09147_ (.A(_00301_),
    .B(_00526_),
    .Y(_03201_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(_00303_),
    .B(net20),
    .Y(_03202_));
 sky130_fd_sc_hd__xor2_1 _09149_ (.A(_03201_),
    .B(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__a21o_1 _09150_ (.A1(_00306_),
    .A2(_05049_),
    .B1(_03203_),
    .X(_03205_));
 sky130_fd_sc_hd__nand3_1 _09151_ (.A(_03203_),
    .B(_00306_),
    .C(_05049_),
    .Y(_03206_));
 sky130_fd_sc_hd__nand2_1 _09152_ (.A(_03205_),
    .B(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__nand2_1 _09153_ (.A(_03200_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__nand3b_1 _09154_ (.A_N(_03207_),
    .B(_03198_),
    .C(_03199_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_1 _09155_ (.A(_03208_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_1 _09156_ (.A(_02596_),
    .B(_02578_),
    .Y(_03211_));
 sky130_fd_sc_hd__inv_2 _09157_ (.A(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(_03210_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__nand3_1 _09159_ (.A(_03211_),
    .B(_03208_),
    .C(_03209_),
    .Y(_03214_));
 sky130_fd_sc_hd__nand2_1 _09160_ (.A(_03213_),
    .B(_03214_),
    .Y(_03216_));
 sky130_fd_sc_hd__nand2_1 _09161_ (.A(_02203_),
    .B(_00421_),
    .Y(_03217_));
 sky130_fd_sc_hd__inv_2 _09162_ (.A(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__inv_2 _09163_ (.A(_01895_),
    .Y(_03219_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(_00315_),
    .B(_00685_),
    .Y(_03220_));
 sky130_fd_sc_hd__nor3_1 _09165_ (.A(_00560_),
    .B(_03219_),
    .C(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__o21ai_1 _09166_ (.A1(_00560_),
    .A2(_03219_),
    .B1(_03220_),
    .Y(_03222_));
 sky130_fd_sc_hd__nor2b_1 _09167_ (.A(_03221_),
    .B_N(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__or2_1 _09168_ (.A(_03218_),
    .B(_03223_),
    .X(_03224_));
 sky130_fd_sc_hd__nand2_1 _09169_ (.A(_03223_),
    .B(_03218_),
    .Y(_03225_));
 sky130_fd_sc_hd__nand2_1 _09170_ (.A(_03224_),
    .B(_03225_),
    .Y(_03227_));
 sky130_fd_sc_hd__a21oi_1 _09171_ (.A1(_02586_),
    .A2(_02591_),
    .B1(_02585_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_1 _09172_ (.A(_03227_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand3b_1 _09173_ (.A_N(_03228_),
    .B(_03224_),
    .C(_03225_),
    .Y(_03230_));
 sky130_fd_sc_hd__nand2_1 _09174_ (.A(_03229_),
    .B(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__o21a_1 _09175_ (.A1(_02607_),
    .A2(_02608_),
    .B1(_02612_),
    .X(_03232_));
 sky130_fd_sc_hd__nand2_1 _09176_ (.A(_03231_),
    .B(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__nand3b_1 _09177_ (.A_N(_03232_),
    .B(_03229_),
    .C(_03230_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_1 _09178_ (.A(_03233_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__nand2_1 _09179_ (.A(_03216_),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__inv_2 _09180_ (.A(_03235_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand3_1 _09181_ (.A(_03213_),
    .B(_03238_),
    .C(_03214_),
    .Y(_03239_));
 sky130_fd_sc_hd__nand2_1 _09182_ (.A(_03236_),
    .B(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__a21boi_1 _09183_ (.A1(_02624_),
    .A2(_02600_),
    .B1_N(_02602_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _09184_ (.A(_03240_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__nand2_1 _09185_ (.A(_02625_),
    .B(_02602_),
    .Y(_03243_));
 sky130_fd_sc_hd__nand3_1 _09186_ (.A(_03243_),
    .B(_03236_),
    .C(_03239_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand2_1 _09187_ (.A(_03242_),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__nand2_1 _09188_ (.A(_02687_),
    .B(_00520_),
    .Y(_03246_));
 sky130_fd_sc_hd__inv_2 _09189_ (.A(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _09190_ (.A(_05096_),
    .B(_00311_),
    .Y(_03249_));
 sky130_fd_sc_hd__nand2_1 _09191_ (.A(_03039_),
    .B(_00355_),
    .Y(_03250_));
 sky130_fd_sc_hd__xor2_1 _09192_ (.A(_03249_),
    .B(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__or2_1 _09193_ (.A(_03247_),
    .B(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_03251_),
    .B(_03247_),
    .Y(_03253_));
 sky130_fd_sc_hd__a21oi_1 _09195_ (.A1(_02637_),
    .A2(_02641_),
    .B1(_02636_),
    .Y(_03254_));
 sky130_fd_sc_hd__a21bo_1 _09196_ (.A1(_03252_),
    .A2(_03253_),
    .B1_N(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__nand3b_1 _09197_ (.A_N(_03254_),
    .B(_03252_),
    .C(_03253_),
    .Y(_03256_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(_03255_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__nand2_1 _09199_ (.A(_02214_),
    .B(_04645_),
    .Y(_03258_));
 sky130_fd_sc_hd__nand2_1 _09200_ (.A(_05114_),
    .B(_04128_),
    .Y(_03260_));
 sky130_fd_sc_hd__nor3_1 _09201_ (.A(_01267_),
    .B(_02377_),
    .C(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__o21ai_1 _09202_ (.A1(_01267_),
    .A2(_02377_),
    .B1(_03260_),
    .Y(_03262_));
 sky130_fd_sc_hd__inv_2 _09203_ (.A(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_1 _09204_ (.A(_03261_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__xor2_1 _09205_ (.A(_03258_),
    .B(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__nand2_1 _09206_ (.A(_03257_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand3b_1 _09207_ (.A_N(_03265_),
    .B(_03255_),
    .C(_03256_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand2_1 _09208_ (.A(_03266_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_1 _09209_ (.A(_02613_),
    .B(_02614_),
    .Y(_03269_));
 sky130_fd_sc_hd__nor2_1 _09210_ (.A(_02614_),
    .B(_02613_),
    .Y(_03271_));
 sky130_fd_sc_hd__a21oi_2 _09211_ (.A1(_03269_),
    .A2(_02604_),
    .B1(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__inv_2 _09212_ (.A(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__nand2_1 _09213_ (.A(_03268_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand3_1 _09214_ (.A(_03266_),
    .B(_03267_),
    .C(_03272_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand2_1 _09215_ (.A(_03274_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_1 _09216_ (.A(_02659_),
    .B(_02647_),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_1 _09217_ (.A(_03276_),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand3b_1 _09218_ (.A_N(_03277_),
    .B(_03274_),
    .C(_03275_),
    .Y(_03279_));
 sky130_fd_sc_hd__nand2_1 _09219_ (.A(_03278_),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__nand2_1 _09220_ (.A(_03245_),
    .B(_03280_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand3b_1 _09221_ (.A_N(_03280_),
    .B(_03242_),
    .C(_03244_),
    .Y(_03283_));
 sky130_fd_sc_hd__nand3_2 _09222_ (.A(_03187_),
    .B(_03282_),
    .C(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _09223_ (.A(_03282_),
    .B(_03283_),
    .Y(_03285_));
 sky130_fd_sc_hd__a21boi_1 _09224_ (.A1(_02671_),
    .A2(_02629_),
    .B1_N(_02626_),
    .Y(_03286_));
 sky130_fd_sc_hd__nand2_1 _09225_ (.A(_03285_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2_1 _09226_ (.A(_03284_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__inv_2 _09227_ (.A(_01532_),
    .Y(_03289_));
 sky130_fd_sc_hd__nor3_1 _09228_ (.A(_03289_),
    .B(_00188_),
    .C(_02706_),
    .Y(_03290_));
 sky130_fd_sc_hd__inv_2 _09229_ (.A(_02711_),
    .Y(_03291_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(_03105_),
    .B(_04888_),
    .Y(_03293_));
 sky130_fd_sc_hd__inv_2 _09231_ (.A(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__nand2_1 _09232_ (.A(_01532_),
    .B(_04899_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand2_1 _09233_ (.A(_01334_),
    .B(_04897_),
    .Y(_03296_));
 sky130_fd_sc_hd__xor2_1 _09234_ (.A(_03295_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__or2_1 _09235_ (.A(_03294_),
    .B(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(_03297_),
    .B(_03294_),
    .Y(_03299_));
 sky130_fd_sc_hd__inv_2 _09237_ (.A(_02649_),
    .Y(_03300_));
 sky130_fd_sc_hd__a21oi_1 _09238_ (.A1(_02653_),
    .A2(_03300_),
    .B1(_02652_),
    .Y(_03301_));
 sky130_fd_sc_hd__a21o_1 _09239_ (.A1(_03298_),
    .A2(_03299_),
    .B1(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__nand3_1 _09240_ (.A(_03298_),
    .B(_03299_),
    .C(_03301_),
    .Y(_03304_));
 sky130_fd_sc_hd__nand2_1 _09241_ (.A(_03302_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__o21ai_1 _09242_ (.A1(_03290_),
    .A2(_03291_),
    .B1(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__nor2_1 _09243_ (.A(_03290_),
    .B(_03291_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand3_1 _09244_ (.A(_03302_),
    .B(_03307_),
    .C(_03304_),
    .Y(_03308_));
 sky130_fd_sc_hd__nand2_1 _09245_ (.A(_03306_),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__nand2_1 _09246_ (.A(_02712_),
    .B(_02714_),
    .Y(_03310_));
 sky130_fd_sc_hd__nor2_1 _09247_ (.A(_02714_),
    .B(_02712_),
    .Y(_03311_));
 sky130_fd_sc_hd__a21oi_2 _09248_ (.A1(_03310_),
    .A2(_02703_),
    .B1(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__inv_2 _09249_ (.A(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _09250_ (.A(_03309_),
    .B(_03313_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand3_1 _09251_ (.A(_03306_),
    .B(_03312_),
    .C(_03308_),
    .Y(_03316_));
 sky130_fd_sc_hd__nand2_1 _09252_ (.A(_03315_),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__nand2_1 _09253_ (.A(_00138_),
    .B(_04941_),
    .Y(_03318_));
 sky130_fd_sc_hd__inv_2 _09254_ (.A(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(_05278_),
    .B(_04933_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand2_1 _09256_ (.A(_05113_),
    .B(_04936_),
    .Y(_03321_));
 sky130_fd_sc_hd__xor2_1 _09257_ (.A(_03320_),
    .B(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__or2_1 _09258_ (.A(_03319_),
    .B(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_03322_),
    .B(_03319_),
    .Y(_03324_));
 sky130_fd_sc_hd__nand2_1 _09260_ (.A(_03323_),
    .B(_03324_),
    .Y(_03326_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(_02744_),
    .B(_02739_),
    .Y(_03327_));
 sky130_fd_sc_hd__inv_2 _09262_ (.A(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__or2_1 _09263_ (.A(_03326_),
    .B(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__nand2_1 _09264_ (.A(_03328_),
    .B(_03326_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand2_1 _09265_ (.A(_00682_),
    .B(_00893_),
    .Y(_03331_));
 sky130_fd_sc_hd__inv_2 _09266_ (.A(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand2_1 _09267_ (.A(_05191_),
    .B(_05159_),
    .Y(_03333_));
 sky130_fd_sc_hd__nor3_1 _09268_ (.A(_02751_),
    .B(_02802_),
    .C(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__o21ai_1 _09269_ (.A1(_02751_),
    .A2(_02802_),
    .B1(_03333_),
    .Y(_03335_));
 sky130_fd_sc_hd__or2b_1 _09270_ (.A(_03334_),
    .B_N(_03335_),
    .X(_03337_));
 sky130_fd_sc_hd__xor2_1 _09271_ (.A(_03332_),
    .B(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__inv_2 _09272_ (.A(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__a21o_1 _09273_ (.A1(_03329_),
    .A2(_03330_),
    .B1(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__nand3_1 _09274_ (.A(_03329_),
    .B(_03339_),
    .C(_03330_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand2_1 _09275_ (.A(_03340_),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__inv_2 _09276_ (.A(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2_1 _09277_ (.A(_03317_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__nand3_1 _09278_ (.A(_03315_),
    .B(_03342_),
    .C(_03316_),
    .Y(_03345_));
 sky130_fd_sc_hd__nand2_1 _09279_ (.A(_03344_),
    .B(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__nand2_1 _09280_ (.A(_02634_),
    .B(_02662_),
    .Y(_03348_));
 sky130_fd_sc_hd__nor2_1 _09281_ (.A(_02662_),
    .B(_02634_),
    .Y(_03349_));
 sky130_fd_sc_hd__a21oi_2 _09282_ (.A1(_03348_),
    .A2(_02666_),
    .B1(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__inv_2 _09283_ (.A(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _09284_ (.A(_03346_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand3_1 _09285_ (.A(_03344_),
    .B(_03345_),
    .C(_03350_),
    .Y(_03353_));
 sky130_fd_sc_hd__nand2_1 _09286_ (.A(_03352_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__nor2_1 _09287_ (.A(_02725_),
    .B(_02702_),
    .Y(_03355_));
 sky130_fd_sc_hd__inv_2 _09288_ (.A(_02768_),
    .Y(_03356_));
 sky130_fd_sc_hd__nor2_1 _09289_ (.A(_03355_),
    .B(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__inv_2 _09290_ (.A(_03357_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand2_1 _09291_ (.A(_03354_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__nand3_1 _09292_ (.A(_03352_),
    .B(_03353_),
    .C(_03357_),
    .Y(_03361_));
 sky130_fd_sc_hd__nand2_1 _09293_ (.A(_03360_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand2_1 _09294_ (.A(_03288_),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand3b_2 _09295_ (.A_N(_03362_),
    .B(_03284_),
    .C(_03287_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand3_2 _09296_ (.A(_03186_),
    .B(_03363_),
    .C(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__nand2_1 _09297_ (.A(_03363_),
    .B(_03364_),
    .Y(_03366_));
 sky130_fd_sc_hd__a21boi_1 _09298_ (.A1(_02833_),
    .A2(_02677_),
    .B1_N(_02673_),
    .Y(_03367_));
 sky130_fd_sc_hd__nand2_1 _09299_ (.A(_03366_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand3_2 _09300_ (.A(_03185_),
    .B(_03365_),
    .C(_03368_),
    .Y(_03370_));
 sky130_fd_sc_hd__nand2_1 _09301_ (.A(_03365_),
    .B(_03368_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_1 _09302_ (.A(_03371_),
    .B(_03184_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand3_2 _09303_ (.A(_03131_),
    .B(_03370_),
    .C(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__nand2_1 _09304_ (.A(_03372_),
    .B(_03370_),
    .Y(_03374_));
 sky130_fd_sc_hd__a21oi_1 _09305_ (.A1(_03129_),
    .A2(_02992_),
    .B1(_03130_),
    .Y(_03375_));
 sky130_fd_sc_hd__nand2_1 _09306_ (.A(_03374_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand3b_1 _09307_ (.A_N(_03128_),
    .B(_03373_),
    .C(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _09308_ (.A(_03374_),
    .B(_03131_),
    .Y(_03378_));
 sky130_fd_sc_hd__nand3_1 _09309_ (.A(_03372_),
    .B(_03375_),
    .C(_03370_),
    .Y(_03379_));
 sky130_fd_sc_hd__nand3_1 _09310_ (.A(_03378_),
    .B(_03379_),
    .C(_03128_),
    .Y(_03381_));
 sky130_fd_sc_hd__nand2_1 _09311_ (.A(_03377_),
    .B(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__nand2_1 _09312_ (.A(_02996_),
    .B(_03054_),
    .Y(_03383_));
 sky130_fd_sc_hd__nor2_1 _09313_ (.A(_03054_),
    .B(_02996_),
    .Y(_03384_));
 sky130_fd_sc_hd__a21oi_1 _09314_ (.A1(_03383_),
    .A2(_03059_),
    .B1(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__inv_2 _09315_ (.A(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__nand2_2 _09316_ (.A(_03382_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand3_1 _09317_ (.A(_03377_),
    .B(_03385_),
    .C(_03381_),
    .Y(_03388_));
 sky130_fd_sc_hd__nand2_1 _09318_ (.A(_03387_),
    .B(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__inv_2 _09319_ (.A(_03097_),
    .Y(_03390_));
 sky130_fd_sc_hd__nand2_1 _09320_ (.A(_03389_),
    .B(_03390_),
    .Y(_03392_));
 sky130_fd_sc_hd__nand3_1 _09321_ (.A(_03387_),
    .B(_03388_),
    .C(_03097_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_1 _09322_ (.A(_03392_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_1 _09323_ (.A(_03126_),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__nor2_1 _09324_ (.A(_00754_),
    .B(_00752_),
    .Y(_03396_));
 sky130_fd_sc_hd__inv_2 _09325_ (.A(_00759_),
    .Y(_03397_));
 sky130_fd_sc_hd__inv_2 _09326_ (.A(_03109_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_1 _09327_ (.A(_03106_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__nand3_1 _09328_ (.A(_03103_),
    .B(_03104_),
    .C(_03109_),
    .Y(_03400_));
 sky130_fd_sc_hd__nand2_1 _09329_ (.A(_03399_),
    .B(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__nand2_1 _09330_ (.A(_03401_),
    .B(_00745_),
    .Y(_03403_));
 sky130_fd_sc_hd__nand3_1 _09331_ (.A(_03399_),
    .B(_03400_),
    .C(_00744_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand2_1 _09332_ (.A(_03403_),
    .B(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__o21ai_2 _09333_ (.A1(_03396_),
    .A2(_03397_),
    .B1(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__inv_2 _09334_ (.A(_03112_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _09335_ (.A(_03120_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__nand3_1 _09336_ (.A(_03112_),
    .B(_03118_),
    .C(_03119_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand2_1 _09337_ (.A(_03408_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__xnor2_1 _09338_ (.A(_03406_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__nor2_1 _09339_ (.A(_03396_),
    .B(_03397_),
    .Y(_03412_));
 sky130_fd_sc_hd__nand3_1 _09340_ (.A(_03412_),
    .B(_03404_),
    .C(_03403_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_03406_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_1 _09342_ (.A(_03415_),
    .B(_00761_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand3b_1 _09343_ (.A_N(_00761_),
    .B(_03406_),
    .C(_03414_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _09344_ (.A(_03416_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__inv_2 _09345_ (.A(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_1 _09346_ (.A(_03411_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__nor2_1 _09347_ (.A(_03395_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__nand2_1 _09348_ (.A(_02366_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__inv_2 _09349_ (.A(_03124_),
    .Y(_03423_));
 sky130_fd_sc_hd__nand2_1 _09350_ (.A(_03394_),
    .B(_03423_),
    .Y(_03425_));
 sky130_fd_sc_hd__or2_1 _09351_ (.A(_03097_),
    .B(_03389_),
    .X(_03426_));
 sky130_fd_sc_hd__nand2_1 _09352_ (.A(_03425_),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__nor2_1 _09353_ (.A(_00761_),
    .B(_03415_),
    .Y(_03428_));
 sky130_fd_sc_hd__nand3_1 _09354_ (.A(_03406_),
    .B(_03408_),
    .C(_03409_),
    .Y(_03429_));
 sky130_fd_sc_hd__a21oi_1 _09355_ (.A1(_03408_),
    .A2(_03409_),
    .B1(_03406_),
    .Y(_03430_));
 sky130_fd_sc_hd__a21oi_1 _09356_ (.A1(_03428_),
    .A2(_03429_),
    .B1(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__nor2_1 _09357_ (.A(_03431_),
    .B(_03395_),
    .Y(_03432_));
 sky130_fd_sc_hd__nor2_1 _09358_ (.A(_03427_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_1 _09359_ (.A(_03422_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand2_1 _09360_ (.A(_00433_),
    .B(net20),
    .Y(_03436_));
 sky130_fd_sc_hd__and4_1 _09361_ (.A(_00234_),
    .B(_00232_),
    .C(net18),
    .D(net19),
    .X(_03437_));
 sky130_fd_sc_hd__a22o_1 _09362_ (.A1(_00234_),
    .A2(net18),
    .B1(_00232_),
    .B2(net19),
    .X(_03438_));
 sky130_fd_sc_hd__nand2b_1 _09363_ (.A_N(_03437_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__or2_1 _09364_ (.A(_03436_),
    .B(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__nand2_1 _09365_ (.A(_03439_),
    .B(_03436_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(_03440_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__o21a_1 _09367_ (.A1(_03191_),
    .A2(_03192_),
    .B1(_03196_),
    .X(_03443_));
 sky130_fd_sc_hd__nand2_1 _09368_ (.A(_03442_),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand3b_2 _09369_ (.A_N(_03443_),
    .B(_03440_),
    .C(_03441_),
    .Y(_03445_));
 sky130_fd_sc_hd__nand2_1 _09370_ (.A(_00306_),
    .B(_00526_),
    .Y(_03447_));
 sky130_fd_sc_hd__inv_2 _09371_ (.A(net21),
    .Y(_03448_));
 sky130_fd_sc_hd__nand2_1 _09372_ (.A(_00301_),
    .B(net17),
    .Y(_03449_));
 sky130_fd_sc_hd__nor3_1 _09373_ (.A(_02310_),
    .B(_03448_),
    .C(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__o21ai_1 _09374_ (.A1(_02310_),
    .A2(_03448_),
    .B1(_03449_),
    .Y(_03451_));
 sky130_fd_sc_hd__and2b_1 _09375_ (.A_N(_03450_),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__xor2_1 _09376_ (.A(_03447_),
    .B(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__inv_2 _09377_ (.A(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__a21o_1 _09378_ (.A1(_03444_),
    .A2(_03445_),
    .B1(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__nand3_2 _09379_ (.A(_03444_),
    .B(_03445_),
    .C(_03454_),
    .Y(_03456_));
 sky130_fd_sc_hd__nand2_1 _09380_ (.A(_03455_),
    .B(_03456_),
    .Y(_03458_));
 sky130_fd_sc_hd__and2_1 _09381_ (.A(_03209_),
    .B(_03199_),
    .X(_03459_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(_03458_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__nand3b_1 _09383_ (.A_N(_03459_),
    .B(_03455_),
    .C(_03456_),
    .Y(_03461_));
 sky130_fd_sc_hd__nand2_1 _09384_ (.A(_03460_),
    .B(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(_02203_),
    .B(_00685_),
    .Y(_03463_));
 sky130_fd_sc_hd__and4_1 _09386_ (.A(_05068_),
    .B(_00315_),
    .C(_01895_),
    .D(_05049_),
    .X(_03464_));
 sky130_fd_sc_hd__a22o_1 _09387_ (.A1(_05068_),
    .A2(_05049_),
    .B1(_00315_),
    .B2(_01895_),
    .X(_03465_));
 sky130_fd_sc_hd__nand2b_1 _09388_ (.A_N(_03464_),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__or2_1 _09389_ (.A(_03463_),
    .B(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__nand2_1 _09390_ (.A(_03466_),
    .B(_03463_),
    .Y(_03469_));
 sky130_fd_sc_hd__nand2_1 _09391_ (.A(_03467_),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__inv_2 _09392_ (.A(net20),
    .Y(_03471_));
 sky130_fd_sc_hd__nor3_1 _09393_ (.A(_02310_),
    .B(_03471_),
    .C(_03201_),
    .Y(_03472_));
 sky130_fd_sc_hd__inv_2 _09394_ (.A(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__nand2_1 _09395_ (.A(_03206_),
    .B(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__or2b_1 _09396_ (.A(_03470_),
    .B_N(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__nand3_1 _09397_ (.A(_03470_),
    .B(_03473_),
    .C(_03206_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _09398_ (.A(_03475_),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__inv_2 _09399_ (.A(_03225_),
    .Y(_03478_));
 sky130_fd_sc_hd__nor2_1 _09400_ (.A(_03221_),
    .B(_03478_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2_1 _09401_ (.A(_03477_),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__inv_2 _09402_ (.A(_03480_),
    .Y(_03482_));
 sky130_fd_sc_hd__nand3_1 _09403_ (.A(_03475_),
    .B(_03482_),
    .C(_03476_),
    .Y(_03483_));
 sky130_fd_sc_hd__nand2_1 _09404_ (.A(_03481_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__nand2_1 _09405_ (.A(_03462_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__inv_2 _09406_ (.A(_03484_),
    .Y(_03486_));
 sky130_fd_sc_hd__nand3_1 _09407_ (.A(_03460_),
    .B(_03461_),
    .C(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__nand2_1 _09408_ (.A(_03485_),
    .B(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__and2_1 _09409_ (.A(_03239_),
    .B(_03214_),
    .X(_03489_));
 sky130_fd_sc_hd__nand2_1 _09410_ (.A(_03488_),
    .B(_03489_),
    .Y(_03491_));
 sky130_fd_sc_hd__nand3b_2 _09411_ (.A_N(_03489_),
    .B(_03485_),
    .C(_03487_),
    .Y(_03492_));
 sky130_fd_sc_hd__nand2_1 _09412_ (.A(_03491_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__o21a_1 _09413_ (.A1(_03249_),
    .A2(_03250_),
    .B1(_03253_),
    .X(_03494_));
 sky130_fd_sc_hd__nand2_1 _09414_ (.A(_02687_),
    .B(_00311_),
    .Y(_03495_));
 sky130_fd_sc_hd__inv_2 _09415_ (.A(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__and4_1 _09416_ (.A(_03039_),
    .B(_05096_),
    .C(_00355_),
    .D(_00421_),
    .X(_03497_));
 sky130_fd_sc_hd__inv_2 _09417_ (.A(_03497_),
    .Y(_03498_));
 sky130_fd_sc_hd__a22o_1 _09418_ (.A1(_03039_),
    .A2(_00421_),
    .B1(_05096_),
    .B2(_00355_),
    .X(_03499_));
 sky130_fd_sc_hd__and2_1 _09419_ (.A(_03498_),
    .B(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__or2_1 _09420_ (.A(_03496_),
    .B(_03500_),
    .X(_03502_));
 sky130_fd_sc_hd__nand2_1 _09421_ (.A(_03500_),
    .B(_03496_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand2_1 _09422_ (.A(_03502_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__or2_1 _09423_ (.A(_03494_),
    .B(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(_03504_),
    .B(_03494_),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2_1 _09425_ (.A(_03505_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__and4_1 _09426_ (.A(_03248_),
    .B(_05114_),
    .C(_00960_),
    .D(_00520_),
    .X(_03508_));
 sky130_fd_sc_hd__a22o_1 _09427_ (.A1(_03248_),
    .A2(_00520_),
    .B1(_05114_),
    .B2(_00960_),
    .X(_03509_));
 sky130_fd_sc_hd__and2b_1 _09428_ (.A_N(_03508_),
    .B(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__nand2_1 _09429_ (.A(_04128_),
    .B(_04645_),
    .Y(_03511_));
 sky130_fd_sc_hd__or2b_1 _09430_ (.A(_03510_),
    .B_N(_03511_),
    .X(_03513_));
 sky130_fd_sc_hd__or2b_1 _09431_ (.A(_03511_),
    .B_N(_03510_),
    .X(_03514_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(_03513_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _09433_ (.A(_03507_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand3b_1 _09434_ (.A_N(_03515_),
    .B(_03505_),
    .C(_03506_),
    .Y(_03517_));
 sky130_fd_sc_hd__nand2_1 _09435_ (.A(_03516_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2_1 _09436_ (.A(_03234_),
    .B(_03230_),
    .Y(_03519_));
 sky130_fd_sc_hd__nand2_1 _09437_ (.A(_03518_),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__inv_2 _09438_ (.A(_03519_),
    .Y(_03521_));
 sky130_fd_sc_hd__nand3_1 _09439_ (.A(_03516_),
    .B(_03517_),
    .C(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__nand2_1 _09440_ (.A(_03520_),
    .B(_03522_),
    .Y(_03524_));
 sky130_fd_sc_hd__nand2_1 _09441_ (.A(_03267_),
    .B(_03256_),
    .Y(_03525_));
 sky130_fd_sc_hd__nand2_1 _09442_ (.A(_03524_),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand3b_1 _09443_ (.A_N(_03525_),
    .B(_03520_),
    .C(_03522_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_03526_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__nand2_1 _09445_ (.A(_03493_),
    .B(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__inv_2 _09446_ (.A(_03528_),
    .Y(_03530_));
 sky130_fd_sc_hd__nand3_1 _09447_ (.A(_03530_),
    .B(_03491_),
    .C(_03492_),
    .Y(_03531_));
 sky130_fd_sc_hd__nand2_1 _09448_ (.A(_03529_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__and2_1 _09449_ (.A(_03283_),
    .B(_03244_),
    .X(_03533_));
 sky130_fd_sc_hd__nand2_1 _09450_ (.A(_03532_),
    .B(_03533_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand3b_2 _09451_ (.A_N(_03533_),
    .B(_03529_),
    .C(_03531_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_03535_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__nand2_1 _09453_ (.A(_01532_),
    .B(_04888_),
    .Y(_03538_));
 sky130_fd_sc_hd__and4_1 _09454_ (.A(_01334_),
    .B(_02214_),
    .C(_04897_),
    .D(_04899_),
    .X(_03539_));
 sky130_fd_sc_hd__a22o_1 _09455_ (.A1(_01334_),
    .A2(_04899_),
    .B1(_02214_),
    .B2(_04897_),
    .X(_03540_));
 sky130_fd_sc_hd__nand2b_1 _09456_ (.A_N(_03539_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__or2_1 _09457_ (.A(_03538_),
    .B(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__nand2_1 _09458_ (.A(_03541_),
    .B(_03538_),
    .Y(_03543_));
 sky130_fd_sc_hd__inv_2 _09459_ (.A(_03261_),
    .Y(_03544_));
 sky130_fd_sc_hd__o21a_1 _09460_ (.A1(_03258_),
    .A2(_03263_),
    .B1(_03544_),
    .X(_03546_));
 sky130_fd_sc_hd__inv_2 _09461_ (.A(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__a21o_1 _09462_ (.A1(_03542_),
    .A2(_03543_),
    .B1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__nand3_1 _09463_ (.A(_03542_),
    .B(_03543_),
    .C(_03547_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _09464_ (.A(_03548_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__o21a_1 _09465_ (.A1(_03295_),
    .A2(_03296_),
    .B1(_03299_),
    .X(_03551_));
 sky130_fd_sc_hd__nand2_1 _09466_ (.A(_03550_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__nand3b_1 _09467_ (.A_N(_03551_),
    .B(_03548_),
    .C(_03549_),
    .Y(_03553_));
 sky130_fd_sc_hd__nand2_1 _09468_ (.A(_03552_),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__nand2_1 _09469_ (.A(_03298_),
    .B(_03299_),
    .Y(_03555_));
 sky130_fd_sc_hd__or2_1 _09470_ (.A(_03301_),
    .B(_03555_),
    .X(_03557_));
 sky130_fd_sc_hd__nand2_1 _09471_ (.A(_03306_),
    .B(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__nand2_1 _09472_ (.A(_03554_),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__inv_2 _09473_ (.A(_03558_),
    .Y(_03560_));
 sky130_fd_sc_hd__nand3_1 _09474_ (.A(_03552_),
    .B(_03553_),
    .C(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__o21a_1 _09475_ (.A1(_03320_),
    .A2(_03321_),
    .B1(_03324_),
    .X(_03562_));
 sky130_fd_sc_hd__nand2_1 _09476_ (.A(_05278_),
    .B(_04941_),
    .Y(_03563_));
 sky130_fd_sc_hd__and4_1 _09477_ (.A(_03105_),
    .B(_05113_),
    .C(_04936_),
    .D(_04933_),
    .X(_03564_));
 sky130_fd_sc_hd__inv_2 _09478_ (.A(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a22o_1 _09479_ (.A1(_03105_),
    .A2(_04936_),
    .B1(_05113_),
    .B2(_04933_),
    .X(_03566_));
 sky130_fd_sc_hd__nand2_1 _09480_ (.A(_03565_),
    .B(_03566_),
    .Y(_03568_));
 sky130_fd_sc_hd__or2_1 _09481_ (.A(_03563_),
    .B(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__nand2_1 _09482_ (.A(_03568_),
    .B(_03563_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_03569_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__nor2_1 _09484_ (.A(_03562_),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__inv_2 _09485_ (.A(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__nand2_1 _09486_ (.A(_03571_),
    .B(_03562_),
    .Y(_03574_));
 sky130_fd_sc_hd__nand2_1 _09487_ (.A(_00682_),
    .B(_05159_),
    .Y(_03575_));
 sky130_fd_sc_hd__and4_1 _09488_ (.A(net46),
    .B(_05191_),
    .C(_00138_),
    .D(_00329_),
    .X(_03576_));
 sky130_fd_sc_hd__a22o_1 _09489_ (.A1(net46),
    .A2(_00138_),
    .B1(_05191_),
    .B2(_00329_),
    .X(_03577_));
 sky130_fd_sc_hd__and2b_1 _09490_ (.A_N(_03576_),
    .B(_03577_),
    .X(_03579_));
 sky130_fd_sc_hd__xor2_1 _09491_ (.A(_03575_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__inv_2 _09492_ (.A(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__a21o_1 _09493_ (.A1(_03573_),
    .A2(_03574_),
    .B1(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__nand3_1 _09494_ (.A(_03573_),
    .B(_03581_),
    .C(_03574_),
    .Y(_03583_));
 sky130_fd_sc_hd__nand2_1 _09495_ (.A(_03582_),
    .B(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__a21o_1 _09496_ (.A1(_03559_),
    .A2(_03561_),
    .B1(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__nand3_1 _09497_ (.A(_03559_),
    .B(_03561_),
    .C(_03584_),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_1 _09498_ (.A(_03585_),
    .B(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__o21a_1 _09499_ (.A1(_03268_),
    .A2(_03272_),
    .B1(_03278_),
    .X(_03588_));
 sky130_fd_sc_hd__inv_2 _09500_ (.A(_03588_),
    .Y(_03590_));
 sky130_fd_sc_hd__nand2_1 _09501_ (.A(_03587_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__nand3_1 _09502_ (.A(_03585_),
    .B(_03586_),
    .C(_03588_),
    .Y(_03592_));
 sky130_fd_sc_hd__nand2_1 _09503_ (.A(_03591_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__o21ai_2 _09504_ (.A1(_03312_),
    .A2(_03309_),
    .B1(_03344_),
    .Y(_03594_));
 sky130_fd_sc_hd__nand2_1 _09505_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__nand3b_1 _09506_ (.A_N(_03594_),
    .B(_03591_),
    .C(_03592_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_1 _09507_ (.A(_03595_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__nand2_1 _09508_ (.A(_03537_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__inv_2 _09509_ (.A(_03597_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand3_2 _09510_ (.A(_03599_),
    .B(_03535_),
    .C(_03536_),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_1 _09511_ (.A(_03598_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__and2_1 _09512_ (.A(_03364_),
    .B(_03284_),
    .X(_03603_));
 sky130_fd_sc_hd__nand2_1 _09513_ (.A(_03602_),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__nand3b_2 _09514_ (.A_N(_03603_),
    .B(_03598_),
    .C(_03601_),
    .Y(_03605_));
 sky130_fd_sc_hd__nand2_1 _09515_ (.A(_03604_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__a21oi_1 _09516_ (.A1(_03335_),
    .A2(_03332_),
    .B1(_03334_),
    .Y(_03607_));
 sky130_fd_sc_hd__and4_1 _09517_ (.A(net49),
    .B(net50),
    .C(_04814_),
    .D(_04880_),
    .X(_03608_));
 sky130_fd_sc_hd__inv_2 _09518_ (.A(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__a22o_1 _09519_ (.A1(net49),
    .A2(_00893_),
    .B1(net50),
    .B2(_00384_),
    .X(_03610_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(_03609_),
    .B(_03610_),
    .Y(_03612_));
 sky130_fd_sc_hd__inv_2 _09521_ (.A(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__nand2_1 _09522_ (.A(net51),
    .B(_00381_),
    .Y(_03614_));
 sky130_fd_sc_hd__inv_2 _09523_ (.A(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _09524_ (.A(_03613_),
    .B(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_1 _09525_ (.A(_03612_),
    .B(_03614_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _09526_ (.A(_03616_),
    .B(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__or2_1 _09527_ (.A(_03607_),
    .B(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__nand2_1 _09528_ (.A(_03618_),
    .B(_03607_),
    .Y(_03620_));
 sky130_fd_sc_hd__o21a_1 _09529_ (.A1(_03141_),
    .A2(_03142_),
    .B1(_03145_),
    .X(_03621_));
 sky130_fd_sc_hd__inv_2 _09530_ (.A(_03621_),
    .Y(_03623_));
 sky130_fd_sc_hd__a21o_1 _09531_ (.A1(_03619_),
    .A2(_03620_),
    .B1(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__nand3_1 _09532_ (.A(_03619_),
    .B(_03623_),
    .C(_03620_),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_1 _09533_ (.A(_03624_),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand2_1 _09534_ (.A(_03341_),
    .B(_03329_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_03626_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__inv_2 _09536_ (.A(_03627_),
    .Y(_03629_));
 sky130_fd_sc_hd__nand3_1 _09537_ (.A(_03624_),
    .B(_03629_),
    .C(_03625_),
    .Y(_03630_));
 sky130_fd_sc_hd__nand2_1 _09538_ (.A(_03628_),
    .B(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_1 _09539_ (.A(_03144_),
    .B(_03145_),
    .Y(_03632_));
 sky130_fd_sc_hd__o21ai_2 _09540_ (.A1(_03632_),
    .A2(_03146_),
    .B1(_03156_),
    .Y(_03634_));
 sky130_fd_sc_hd__nand2_1 _09541_ (.A(_03631_),
    .B(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__nand3b_1 _09542_ (.A_N(_03634_),
    .B(_03628_),
    .C(_03630_),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(_03635_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__nand2_1 _09544_ (.A(_03165_),
    .B(_03157_),
    .Y(_03638_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_03637_),
    .B(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__inv_2 _09546_ (.A(_03638_),
    .Y(_03640_));
 sky130_fd_sc_hd__nand3_1 _09547_ (.A(_03635_),
    .B(_03636_),
    .C(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__nand2_1 _09548_ (.A(_03639_),
    .B(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__inv_2 _09549_ (.A(net52),
    .Y(_03643_));
 sky130_fd_sc_hd__inv_2 _09550_ (.A(net53),
    .Y(_03645_));
 sky130_fd_sc_hd__or4_2 _09551_ (.A(_03643_),
    .B(_03645_),
    .C(_00187_),
    .D(_02311_),
    .X(_03646_));
 sky130_fd_sc_hd__a22o_1 _09552_ (.A1(net52),
    .A2(_05310_),
    .B1(net53),
    .B2(_00194_),
    .X(_03647_));
 sky130_fd_sc_hd__nand3_1 _09553_ (.A(_03642_),
    .B(_03646_),
    .C(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(_03646_),
    .B(_03647_),
    .Y(_03649_));
 sky130_fd_sc_hd__nand3_1 _09555_ (.A(_03639_),
    .B(_03641_),
    .C(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(_03648_),
    .B(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__nor2_1 _09557_ (.A(_03350_),
    .B(_03346_),
    .Y(_03652_));
 sky130_fd_sc_hd__inv_2 _09558_ (.A(_03360_),
    .Y(_03653_));
 sky130_fd_sc_hd__nor2_1 _09559_ (.A(_03652_),
    .B(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__inv_2 _09560_ (.A(_03654_),
    .Y(_03656_));
 sky130_fd_sc_hd__nand2_1 _09561_ (.A(_03651_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand3_1 _09562_ (.A(_03648_),
    .B(_03650_),
    .C(_03654_),
    .Y(_03658_));
 sky130_fd_sc_hd__nand2_1 _09563_ (.A(_03657_),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_1 _09564_ (.A(_03175_),
    .B(_03170_),
    .Y(_03660_));
 sky130_fd_sc_hd__nand2_1 _09565_ (.A(_03659_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__nand3b_1 _09566_ (.A_N(_03660_),
    .B(_03657_),
    .C(_03658_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand2_1 _09567_ (.A(_03661_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__nand2_1 _09568_ (.A(_03606_),
    .B(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__inv_2 _09569_ (.A(_03663_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand3_2 _09570_ (.A(_03665_),
    .B(_03604_),
    .C(_03605_),
    .Y(_03667_));
 sky130_fd_sc_hd__nand2_1 _09571_ (.A(_03664_),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__and2_1 _09572_ (.A(_03370_),
    .B(_03365_),
    .X(_03669_));
 sky130_fd_sc_hd__nand2_1 _09573_ (.A(_03668_),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand3b_1 _09574_ (.A_N(_03669_),
    .B(_03664_),
    .C(_03667_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _09575_ (.A(_03670_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_1 _09576_ (.A(_03183_),
    .B(_03178_),
    .Y(_03673_));
 sky130_fd_sc_hd__inv_2 _09577_ (.A(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__nand2_1 _09578_ (.A(_03672_),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand3_1 _09579_ (.A(_03670_),
    .B(_03671_),
    .C(_03673_),
    .Y(_03676_));
 sky130_fd_sc_hd__nand2_1 _09580_ (.A(_03675_),
    .B(_03676_),
    .Y(_03678_));
 sky130_fd_sc_hd__nand3_1 _09581_ (.A(_03373_),
    .B(_03376_),
    .C(_03128_),
    .Y(_03679_));
 sky130_fd_sc_hd__nand3_1 _09582_ (.A(_03678_),
    .B(_03373_),
    .C(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__nand2_1 _09583_ (.A(_03679_),
    .B(_03373_),
    .Y(_03681_));
 sky130_fd_sc_hd__nand3_2 _09584_ (.A(_03675_),
    .B(_03676_),
    .C(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _09585_ (.A(_03680_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_03683_),
    .B(_03387_),
    .Y(_03684_));
 sky130_fd_sc_hd__inv_2 _09587_ (.A(_03387_),
    .Y(_03685_));
 sky130_fd_sc_hd__nand3_2 _09588_ (.A(_03680_),
    .B(_03685_),
    .C(_03682_),
    .Y(_03686_));
 sky130_fd_sc_hd__nand2_1 _09589_ (.A(_03684_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__nand2_1 _09590_ (.A(_02687_),
    .B(_00355_),
    .Y(_03689_));
 sky130_fd_sc_hd__and4_1 _09591_ (.A(_03039_),
    .B(_05096_),
    .C(_00421_),
    .D(_00685_),
    .X(_03690_));
 sky130_fd_sc_hd__inv_2 _09592_ (.A(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__a22o_1 _09593_ (.A1(_03039_),
    .A2(_00685_),
    .B1(_05096_),
    .B2(_00421_),
    .X(_03692_));
 sky130_fd_sc_hd__nand2_1 _09594_ (.A(_03691_),
    .B(_03692_),
    .Y(_03693_));
 sky130_fd_sc_hd__or2_1 _09595_ (.A(_03689_),
    .B(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__nand2_1 _09596_ (.A(_03693_),
    .B(_03689_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_1 _09597_ (.A(_03694_),
    .B(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__and2_1 _09598_ (.A(_03503_),
    .B(_03498_),
    .X(_03697_));
 sky130_fd_sc_hd__or2_1 _09599_ (.A(_03696_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_03697_),
    .B(_03696_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand2_1 _09601_ (.A(_03698_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__nand2_1 _09602_ (.A(_04645_),
    .B(_00960_),
    .Y(_03702_));
 sky130_fd_sc_hd__and4_1 _09603_ (.A(_03248_),
    .B(_05114_),
    .C(_00520_),
    .D(_00311_),
    .X(_03703_));
 sky130_fd_sc_hd__inv_2 _09604_ (.A(_03703_),
    .Y(_03704_));
 sky130_fd_sc_hd__a22o_1 _09605_ (.A1(_03248_),
    .A2(_00311_),
    .B1(_05114_),
    .B2(_00520_),
    .X(_03705_));
 sky130_fd_sc_hd__nand2_1 _09606_ (.A(_03704_),
    .B(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__xnor2_1 _09607_ (.A(_03702_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__nand2_1 _09608_ (.A(_03701_),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__nand3b_1 _09609_ (.A_N(_03707_),
    .B(_03698_),
    .C(_03700_),
    .Y(_03709_));
 sky130_fd_sc_hd__nand2_1 _09610_ (.A(_03708_),
    .B(_03709_),
    .Y(_03711_));
 sky130_fd_sc_hd__and2_1 _09611_ (.A(_03483_),
    .B(_03475_),
    .X(_03712_));
 sky130_fd_sc_hd__nor2_1 _09612_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__nand2_1 _09613_ (.A(_03712_),
    .B(_03711_),
    .Y(_03714_));
 sky130_fd_sc_hd__inv_2 _09614_ (.A(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__nand2_1 _09615_ (.A(_03517_),
    .B(_03505_),
    .Y(_03716_));
 sky130_fd_sc_hd__o21bai_1 _09616_ (.A1(_03713_),
    .A2(_03715_),
    .B1_N(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__nand3b_1 _09617_ (.A_N(_03713_),
    .B(_03716_),
    .C(_03714_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_1 _09618_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__inv_2 _09619_ (.A(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand2_1 _09620_ (.A(_03487_),
    .B(_03461_),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _09621_ (.A(_00433_),
    .B(net21),
    .Y(_03723_));
 sky130_fd_sc_hd__and4_1 _09622_ (.A(_00234_),
    .B(_00232_),
    .C(net19),
    .D(net20),
    .X(_03724_));
 sky130_fd_sc_hd__a22o_1 _09623_ (.A1(_00234_),
    .A2(net19),
    .B1(_00232_),
    .B2(net20),
    .X(_03725_));
 sky130_fd_sc_hd__nand2b_1 _09624_ (.A_N(_03724_),
    .B(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__or2_1 _09625_ (.A(_03723_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__nand2_1 _09626_ (.A(_03726_),
    .B(_03723_),
    .Y(_03728_));
 sky130_fd_sc_hd__a31o_1 _09627_ (.A1(_03438_),
    .A2(_00433_),
    .A3(net20),
    .B1(_03437_),
    .X(_03729_));
 sky130_fd_sc_hd__a21o_1 _09628_ (.A1(_03727_),
    .A2(_03728_),
    .B1(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__nand3_1 _09629_ (.A(_03727_),
    .B(_03729_),
    .C(_03728_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand2_1 _09630_ (.A(_03730_),
    .B(_03731_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand2_1 _09631_ (.A(_00306_),
    .B(net17),
    .Y(_03734_));
 sky130_fd_sc_hd__and4_1 _09632_ (.A(_00303_),
    .B(_00301_),
    .C(net18),
    .D(net22),
    .X(_03735_));
 sky130_fd_sc_hd__inv_2 _09633_ (.A(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__a22o_1 _09634_ (.A1(_00303_),
    .A2(net22),
    .B1(_00301_),
    .B2(net18),
    .X(_03737_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_03736_),
    .B(_03737_),
    .Y(_03738_));
 sky130_fd_sc_hd__xnor2_1 _09636_ (.A(_03734_),
    .B(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_03733_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__nand3b_1 _09638_ (.A_N(_03739_),
    .B(_03730_),
    .C(_03731_),
    .Y(_03741_));
 sky130_fd_sc_hd__nand2_1 _09639_ (.A(_03740_),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand3_1 _09640_ (.A(_03742_),
    .B(_03445_),
    .C(_03456_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(_03456_),
    .B(_03445_),
    .Y(_03745_));
 sky130_fd_sc_hd__nand3_1 _09642_ (.A(_03740_),
    .B(_03741_),
    .C(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__nand2_1 _09643_ (.A(_03744_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__a31oi_1 _09644_ (.A1(_03451_),
    .A2(_00306_),
    .A3(_00526_),
    .B1(_03450_),
    .Y(_03748_));
 sky130_fd_sc_hd__nand2_1 _09645_ (.A(_02203_),
    .B(_01895_),
    .Y(_03749_));
 sky130_fd_sc_hd__and4_1 _09646_ (.A(_05068_),
    .B(_00315_),
    .C(_05049_),
    .D(_00526_),
    .X(_03750_));
 sky130_fd_sc_hd__inv_2 _09647_ (.A(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__a22o_1 _09648_ (.A1(_05068_),
    .A2(_00526_),
    .B1(_00315_),
    .B2(_05049_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_1 _09649_ (.A(_03751_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__or2_1 _09650_ (.A(_03749_),
    .B(_03753_),
    .X(_03755_));
 sky130_fd_sc_hd__nand2_1 _09651_ (.A(_03753_),
    .B(_03749_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_1 _09652_ (.A(_03755_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__nor2_1 _09653_ (.A(_03748_),
    .B(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__inv_2 _09654_ (.A(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__nand2_1 _09655_ (.A(_03757_),
    .B(_03748_),
    .Y(_03760_));
 sky130_fd_sc_hd__a31o_1 _09656_ (.A1(_03465_),
    .A2(_02203_),
    .A3(_00685_),
    .B1(_03464_),
    .X(_03761_));
 sky130_fd_sc_hd__a21o_1 _09657_ (.A1(_03759_),
    .A2(_03760_),
    .B1(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__nand3_1 _09658_ (.A(_03759_),
    .B(_03761_),
    .C(_03760_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand2_1 _09659_ (.A(_03762_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__nand2_1 _09660_ (.A(_03747_),
    .B(_03764_),
    .Y(_03766_));
 sky130_fd_sc_hd__nand3b_2 _09661_ (.A_N(_03764_),
    .B(_03744_),
    .C(_03746_),
    .Y(_03767_));
 sky130_fd_sc_hd__nand3_2 _09662_ (.A(_03722_),
    .B(_03766_),
    .C(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand2_1 _09663_ (.A(_03766_),
    .B(_03767_),
    .Y(_03769_));
 sky130_fd_sc_hd__inv_2 _09664_ (.A(_03722_),
    .Y(_03770_));
 sky130_fd_sc_hd__nand2_1 _09665_ (.A(_03769_),
    .B(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__nand3_2 _09666_ (.A(_03720_),
    .B(_03768_),
    .C(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand2_1 _09667_ (.A(_03771_),
    .B(_03768_),
    .Y(_03773_));
 sky130_fd_sc_hd__nand2_1 _09668_ (.A(_03773_),
    .B(_03719_),
    .Y(_03774_));
 sky130_fd_sc_hd__nand2_1 _09669_ (.A(_03772_),
    .B(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(_03531_),
    .B(_03492_),
    .Y(_03777_));
 sky130_fd_sc_hd__inv_2 _09671_ (.A(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__nand2_1 _09672_ (.A(_03775_),
    .B(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__nand3_2 _09673_ (.A(_03777_),
    .B(_03772_),
    .C(_03774_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2_1 _09674_ (.A(_03779_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__a31o_1 _09675_ (.A1(_03509_),
    .A2(_04128_),
    .A3(_04645_),
    .B1(_03508_),
    .X(_03782_));
 sky130_fd_sc_hd__inv_2 _09676_ (.A(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _09677_ (.A(_01334_),
    .B(_04888_),
    .Y(_03784_));
 sky130_fd_sc_hd__and4_1 _09678_ (.A(_02214_),
    .B(_04128_),
    .C(_04897_),
    .D(_04899_),
    .X(_03785_));
 sky130_fd_sc_hd__inv_2 _09679_ (.A(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__a22o_1 _09680_ (.A1(_02214_),
    .A2(_04899_),
    .B1(_04128_),
    .B2(_04897_),
    .X(_03788_));
 sky130_fd_sc_hd__nand2_1 _09681_ (.A(_03786_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__or2_1 _09682_ (.A(_03784_),
    .B(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__nand2_1 _09683_ (.A(_03789_),
    .B(_03784_),
    .Y(_03791_));
 sky130_fd_sc_hd__nand2_1 _09684_ (.A(_03790_),
    .B(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__nor2_1 _09685_ (.A(_03783_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__inv_2 _09686_ (.A(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__nand2_1 _09687_ (.A(_03792_),
    .B(_03783_),
    .Y(_03795_));
 sky130_fd_sc_hd__a31o_1 _09688_ (.A1(_03540_),
    .A2(_01532_),
    .A3(_04888_),
    .B1(_03539_),
    .X(_03796_));
 sky130_fd_sc_hd__a21o_1 _09689_ (.A1(_03794_),
    .A2(_03795_),
    .B1(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__nand3_1 _09690_ (.A(_03794_),
    .B(_03796_),
    .C(_03795_),
    .Y(_03799_));
 sky130_fd_sc_hd__nand2_1 _09691_ (.A(_03797_),
    .B(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__nand2_1 _09692_ (.A(_03553_),
    .B(_03549_),
    .Y(_03801_));
 sky130_fd_sc_hd__inv_2 _09693_ (.A(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2b_1 _09694_ (.A_N(_03800_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _09695_ (.A(_03800_),
    .B(_03801_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand2_1 _09696_ (.A(_03803_),
    .B(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__nand2_1 _09697_ (.A(_05113_),
    .B(_04941_),
    .Y(_03806_));
 sky130_fd_sc_hd__inv_2 _09698_ (.A(_04933_),
    .Y(_03807_));
 sky130_fd_sc_hd__or4_1 _09699_ (.A(_02679_),
    .B(_03289_),
    .C(_05179_),
    .D(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__a22o_1 _09700_ (.A1(_03105_),
    .A2(_04933_),
    .B1(_01532_),
    .B2(_04936_),
    .X(_03810_));
 sky130_fd_sc_hd__nand2_1 _09701_ (.A(_03808_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__or2_1 _09702_ (.A(_03806_),
    .B(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__nand2_1 _09703_ (.A(_03811_),
    .B(_03806_),
    .Y(_03813_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_03812_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__nand2_1 _09705_ (.A(_03569_),
    .B(_03565_),
    .Y(_03815_));
 sky130_fd_sc_hd__inv_2 _09706_ (.A(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _09707_ (.A(_03814_),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand3_1 _09708_ (.A(_03812_),
    .B(_03815_),
    .C(_03813_),
    .Y(_03818_));
 sky130_fd_sc_hd__nand2_1 _09709_ (.A(_03817_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__nand2_1 _09710_ (.A(_00682_),
    .B(_00329_),
    .Y(_03821_));
 sky130_fd_sc_hd__inv_2 _09711_ (.A(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__and4_1 _09712_ (.A(net46),
    .B(_05191_),
    .C(_05278_),
    .D(_00138_),
    .X(_03823_));
 sky130_fd_sc_hd__a22o_1 _09713_ (.A1(net46),
    .A2(_05278_),
    .B1(_05191_),
    .B2(_00138_),
    .X(_03824_));
 sky130_fd_sc_hd__or2b_1 _09714_ (.A(_03823_),
    .B_N(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__xor2_1 _09715_ (.A(_03822_),
    .B(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__nand2_1 _09716_ (.A(_03819_),
    .B(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__inv_2 _09717_ (.A(_03826_),
    .Y(_03828_));
 sky130_fd_sc_hd__nand3_1 _09718_ (.A(_03817_),
    .B(_03828_),
    .C(_03818_),
    .Y(_03829_));
 sky130_fd_sc_hd__nand2_1 _09719_ (.A(_03827_),
    .B(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__inv_2 _09720_ (.A(_03830_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _09721_ (.A(_03805_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand3_1 _09722_ (.A(_03803_),
    .B(_03830_),
    .C(_03804_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_1 _09723_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__nand2_1 _09724_ (.A(_03518_),
    .B(_03521_),
    .Y(_03836_));
 sky130_fd_sc_hd__nor2_1 _09725_ (.A(_03521_),
    .B(_03518_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21oi_2 _09726_ (.A1(_03836_),
    .A2(_03525_),
    .B1(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__inv_2 _09727_ (.A(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__nand2_1 _09728_ (.A(_03835_),
    .B(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__nand3_1 _09729_ (.A(_03833_),
    .B(_03834_),
    .C(_03838_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2_1 _09730_ (.A(_03840_),
    .B(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__o21ai_2 _09731_ (.A1(_03560_),
    .A2(_03554_),
    .B1(_03585_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _09732_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__nand3b_1 _09733_ (.A_N(_03844_),
    .B(_03840_),
    .C(_03841_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_1 _09734_ (.A(_03845_),
    .B(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__nand2_1 _09735_ (.A(_03781_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__inv_2 _09736_ (.A(_03847_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand3_2 _09737_ (.A(_03849_),
    .B(_03779_),
    .C(_03780_),
    .Y(_03850_));
 sky130_fd_sc_hd__nand2_1 _09738_ (.A(_03848_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__nand2_1 _09739_ (.A(_03601_),
    .B(_03536_),
    .Y(_03852_));
 sky130_fd_sc_hd__inv_2 _09740_ (.A(_03852_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_03851_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand3_2 _09742_ (.A(_03852_),
    .B(_03848_),
    .C(_03850_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand2_1 _09743_ (.A(_03855_),
    .B(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__and2_1 _09744_ (.A(_03583_),
    .B(_03573_),
    .X(_03858_));
 sky130_fd_sc_hd__and4_1 _09745_ (.A(net49),
    .B(net50),
    .C(_05159_),
    .D(_00893_),
    .X(_03859_));
 sky130_fd_sc_hd__inv_2 _09746_ (.A(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__a22o_1 _09747_ (.A1(net49),
    .A2(_05159_),
    .B1(net50),
    .B2(_00893_),
    .X(_03861_));
 sky130_fd_sc_hd__nand2_1 _09748_ (.A(_03860_),
    .B(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _09749_ (.A(net51),
    .B(_00384_),
    .Y(_03863_));
 sky130_fd_sc_hd__inv_2 _09750_ (.A(_03863_),
    .Y(_03865_));
 sky130_fd_sc_hd__nand2b_1 _09751_ (.A_N(_03862_),
    .B(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _09752_ (.A(_03862_),
    .B(_03863_),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _09753_ (.A(_03866_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__a31o_1 _09754_ (.A1(_03577_),
    .A2(_00682_),
    .A3(_05159_),
    .B1(_03576_),
    .X(_03869_));
 sky130_fd_sc_hd__inv_2 _09755_ (.A(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__nor2_1 _09756_ (.A(_03868_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__inv_2 _09757_ (.A(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__nand2_1 _09758_ (.A(_03870_),
    .B(_03868_),
    .Y(_03873_));
 sky130_fd_sc_hd__nand2_1 _09759_ (.A(_03616_),
    .B(_03609_),
    .Y(_03874_));
 sky130_fd_sc_hd__a21o_1 _09760_ (.A1(_03872_),
    .A2(_03873_),
    .B1(_03874_),
    .X(_03876_));
 sky130_fd_sc_hd__nand3_1 _09761_ (.A(_03872_),
    .B(_03874_),
    .C(_03873_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _09762_ (.A(_03876_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__nor2_1 _09763_ (.A(_03858_),
    .B(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__nand2_1 _09764_ (.A(_03878_),
    .B(_03858_),
    .Y(_03880_));
 sky130_fd_sc_hd__inv_2 _09765_ (.A(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__nand2_1 _09766_ (.A(_03625_),
    .B(_03619_),
    .Y(_03882_));
 sky130_fd_sc_hd__o21bai_1 _09767_ (.A1(_03879_),
    .A2(_03881_),
    .B1_N(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__nand3b_1 _09768_ (.A_N(_03879_),
    .B(_03882_),
    .C(_03880_),
    .Y(_03884_));
 sky130_fd_sc_hd__nand2_1 _09769_ (.A(_03883_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _09770_ (.A(_03626_),
    .B(_03629_),
    .Y(_03887_));
 sky130_fd_sc_hd__nor2_1 _09771_ (.A(_03629_),
    .B(_03626_),
    .Y(_03888_));
 sky130_fd_sc_hd__a21oi_2 _09772_ (.A1(_03887_),
    .A2(_03634_),
    .B1(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__inv_2 _09773_ (.A(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _09774_ (.A(_03885_),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__nand3_1 _09775_ (.A(_03883_),
    .B(_03884_),
    .C(_03889_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _09776_ (.A(_03891_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__inv_2 _09777_ (.A(net54),
    .Y(_03894_));
 sky130_fd_sc_hd__and4_1 _09778_ (.A(net52),
    .B(net53),
    .C(_00381_),
    .D(_04947_),
    .X(_03895_));
 sky130_fd_sc_hd__inv_2 _09779_ (.A(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__a22o_1 _09780_ (.A1(net52),
    .A2(_00381_),
    .B1(net53),
    .B2(_05310_),
    .X(_03898_));
 sky130_fd_sc_hd__nand2_1 _09781_ (.A(_03896_),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__or3_1 _09782_ (.A(_03894_),
    .B(_02311_),
    .C(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__o21ai_1 _09783_ (.A1(_03894_),
    .A2(_02311_),
    .B1(_03899_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _09784_ (.A(_03900_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__or2_1 _09785_ (.A(_03646_),
    .B(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__nand2_1 _09786_ (.A(_03902_),
    .B(_03646_),
    .Y(_03904_));
 sky130_fd_sc_hd__nand2_1 _09787_ (.A(_03903_),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__inv_2 _09788_ (.A(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__nand2_1 _09789_ (.A(_03893_),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__nand3_1 _09790_ (.A(_03891_),
    .B(_03892_),
    .C(_03905_),
    .Y(_03909_));
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(_03907_),
    .B(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _09792_ (.A(_03587_),
    .B(_03588_),
    .Y(_03911_));
 sky130_fd_sc_hd__nor2_1 _09793_ (.A(_03588_),
    .B(_03587_),
    .Y(_03912_));
 sky130_fd_sc_hd__a21oi_2 _09794_ (.A1(_03911_),
    .A2(_03594_),
    .B1(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__inv_2 _09795_ (.A(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__nand2_1 _09796_ (.A(_03910_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand3_1 _09797_ (.A(_03907_),
    .B(_03913_),
    .C(_03909_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2_1 _09798_ (.A(_03915_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__nor2_1 _09799_ (.A(_03640_),
    .B(_03637_),
    .Y(_03918_));
 sky130_fd_sc_hd__inv_2 _09800_ (.A(_03648_),
    .Y(_03920_));
 sky130_fd_sc_hd__nor2_1 _09801_ (.A(_03918_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__inv_2 _09802_ (.A(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__nand2_1 _09803_ (.A(_03917_),
    .B(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand3_1 _09804_ (.A(_03915_),
    .B(_03921_),
    .C(_03916_),
    .Y(_03924_));
 sky130_fd_sc_hd__nand2_1 _09805_ (.A(_03923_),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _09806_ (.A(_03857_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__inv_2 _09807_ (.A(_03925_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand3_1 _09808_ (.A(_03927_),
    .B(_03855_),
    .C(_03856_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand2_1 _09809_ (.A(_03926_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _09810_ (.A(_03667_),
    .B(_03605_),
    .Y(_03931_));
 sky130_fd_sc_hd__inv_2 _09811_ (.A(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _09812_ (.A(_03929_),
    .B(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__nand3_1 _09813_ (.A(_03931_),
    .B(_03926_),
    .C(_03928_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand2_1 _09814_ (.A(_03933_),
    .B(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__nor2_1 _09815_ (.A(_03654_),
    .B(_03651_),
    .Y(_03936_));
 sky130_fd_sc_hd__inv_2 _09816_ (.A(_03661_),
    .Y(_03937_));
 sky130_fd_sc_hd__nor2_1 _09817_ (.A(_03936_),
    .B(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__nand2_2 _09818_ (.A(_03935_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__nand3b_2 _09819_ (.A_N(_03938_),
    .B(_03933_),
    .C(_03934_),
    .Y(_03940_));
 sky130_fd_sc_hd__nand2_1 _09820_ (.A(_03939_),
    .B(_03940_),
    .Y(_03942_));
 sky130_fd_sc_hd__nand2_1 _09821_ (.A(_03676_),
    .B(_03671_),
    .Y(_03943_));
 sky130_fd_sc_hd__inv_2 _09822_ (.A(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__nand2_1 _09823_ (.A(_03942_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__nand3_1 _09824_ (.A(_03943_),
    .B(_03939_),
    .C(_03940_),
    .Y(_03946_));
 sky130_fd_sc_hd__nand2_1 _09825_ (.A(_03945_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _09826_ (.A(_03947_),
    .B(_03682_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand3b_1 _09827_ (.A_N(_03682_),
    .B(_03945_),
    .C(_03946_),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_2 _09828_ (.A(_03948_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__nor2_1 _09829_ (.A(_03687_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__nand2_1 _09830_ (.A(_03434_),
    .B(_03951_),
    .Y(_03953_));
 sky130_fd_sc_hd__nor2_1 _09831_ (.A(_03682_),
    .B(_03947_),
    .Y(_03954_));
 sky130_fd_sc_hd__nor2_1 _09832_ (.A(_03686_),
    .B(_03950_),
    .Y(_03955_));
 sky130_fd_sc_hd__nor2_1 _09833_ (.A(_03954_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand2_1 _09834_ (.A(_03953_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__and2_1 _09835_ (.A(_03940_),
    .B(_03934_),
    .X(_03958_));
 sky130_fd_sc_hd__nand2_1 _09836_ (.A(_03928_),
    .B(_03856_),
    .Y(_03959_));
 sky130_fd_sc_hd__inv_2 _09837_ (.A(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__a21boi_2 _09838_ (.A1(_03817_),
    .A2(_03828_),
    .B1_N(_03818_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand2_1 _09839_ (.A(_03866_),
    .B(_03860_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(net51),
    .B(_00893_),
    .Y(_03964_));
 sky130_fd_sc_hd__inv_2 _09841_ (.A(net50),
    .Y(_03965_));
 sky130_fd_sc_hd__or4_2 _09842_ (.A(_03148_),
    .B(_03965_),
    .C(_02802_),
    .D(_02752_),
    .X(_03966_));
 sky130_fd_sc_hd__a22o_1 _09843_ (.A1(net49),
    .A2(_00329_),
    .B1(net50),
    .B2(_05159_),
    .X(_03967_));
 sky130_fd_sc_hd__nand2_1 _09844_ (.A(_03966_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__or2_1 _09845_ (.A(_03964_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__nand2_1 _09846_ (.A(_03968_),
    .B(_03964_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _09847_ (.A(_03969_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__a21oi_2 _09848_ (.A1(_03824_),
    .A2(_03822_),
    .B1(_03823_),
    .Y(_03972_));
 sky130_fd_sc_hd__inv_2 _09849_ (.A(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _09850_ (.A(_03971_),
    .B(_03973_),
    .Y(_03975_));
 sky130_fd_sc_hd__nand3_1 _09851_ (.A(_03969_),
    .B(_03972_),
    .C(_03970_),
    .Y(_03976_));
 sky130_fd_sc_hd__nand3b_1 _09852_ (.A_N(_03962_),
    .B(_03975_),
    .C(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand2_1 _09853_ (.A(_03971_),
    .B(_03972_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand3_1 _09854_ (.A(_03969_),
    .B(_03970_),
    .C(_03973_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand3_1 _09855_ (.A(_03978_),
    .B(_03962_),
    .C(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(_03977_),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__nor2_1 _09857_ (.A(_03961_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__inv_2 _09858_ (.A(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _09859_ (.A(_03877_),
    .B(_03872_),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(_03981_),
    .B(_03961_),
    .Y(_03986_));
 sky130_fd_sc_hd__nand3_1 _09861_ (.A(_03983_),
    .B(_03984_),
    .C(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand3_1 _09862_ (.A(_03961_),
    .B(_03977_),
    .C(_03980_),
    .Y(_03988_));
 sky130_fd_sc_hd__inv_2 _09863_ (.A(_03961_),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _09864_ (.A(_03989_),
    .B(_03981_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand3b_1 _09865_ (.A_N(_03984_),
    .B(_03988_),
    .C(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _09866_ (.A(_03987_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__a21oi_2 _09867_ (.A1(_03880_),
    .A2(_03882_),
    .B1(_03879_),
    .Y(_03993_));
 sky130_fd_sc_hd__inv_2 _09868_ (.A(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__nand2_1 _09869_ (.A(_03992_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand3_1 _09870_ (.A(_03987_),
    .B(_03991_),
    .C(_03993_),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_1 _09871_ (.A(_03995_),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__nand2_1 _09872_ (.A(net56),
    .B(_00194_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_1 _09873_ (.A(_03900_),
    .B(_03896_),
    .Y(_04000_));
 sky130_fd_sc_hd__inv_2 _09874_ (.A(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__or4_1 _09875_ (.A(_03643_),
    .B(_03645_),
    .C(_02875_),
    .D(_02309_),
    .X(_04002_));
 sky130_fd_sc_hd__a22o_1 _09876_ (.A1(net52),
    .A2(_00384_),
    .B1(net53),
    .B2(_00381_),
    .X(_04003_));
 sky130_fd_sc_hd__nand2_1 _09877_ (.A(_04002_),
    .B(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand3b_1 _09878_ (.A_N(_04004_),
    .B(net54),
    .C(_05310_),
    .Y(_04005_));
 sky130_fd_sc_hd__o21ai_1 _09879_ (.A1(_03894_),
    .A2(_00187_),
    .B1(_04004_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_1 _09880_ (.A(_04005_),
    .B(_04006_),
    .Y(_04008_));
 sky130_fd_sc_hd__nor2_1 _09881_ (.A(_04001_),
    .B(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__inv_2 _09882_ (.A(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__nand2_1 _09883_ (.A(_04008_),
    .B(_04001_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(_04010_),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__or2_1 _09885_ (.A(_03999_),
    .B(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__nand2_1 _09886_ (.A(_04012_),
    .B(_03999_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_1 _09887_ (.A(_04013_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand2_1 _09888_ (.A(_04015_),
    .B(_03903_),
    .Y(_04016_));
 sky130_fd_sc_hd__nand3b_1 _09889_ (.A_N(_03903_),
    .B(_04013_),
    .C(_04014_),
    .Y(_04017_));
 sky130_fd_sc_hd__nand2_1 _09890_ (.A(_04016_),
    .B(_04017_),
    .Y(_04019_));
 sky130_fd_sc_hd__inv_2 _09891_ (.A(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__nand2_1 _09892_ (.A(_03998_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__nand3_1 _09893_ (.A(_03995_),
    .B(_03997_),
    .C(_04019_),
    .Y(_04022_));
 sky130_fd_sc_hd__nand2_1 _09894_ (.A(_04021_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2_1 _09895_ (.A(_03835_),
    .B(_03838_),
    .Y(_04024_));
 sky130_fd_sc_hd__nor2_1 _09896_ (.A(_03838_),
    .B(_03835_),
    .Y(_04025_));
 sky130_fd_sc_hd__a21oi_2 _09897_ (.A1(_04024_),
    .A2(_03844_),
    .B1(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__inv_2 _09898_ (.A(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__nand2_1 _09899_ (.A(_04023_),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__nand3_1 _09900_ (.A(_04021_),
    .B(_04022_),
    .C(_04026_),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_1 _09901_ (.A(_04028_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__nor2_1 _09902_ (.A(_03889_),
    .B(_03885_),
    .Y(_04032_));
 sky130_fd_sc_hd__inv_2 _09903_ (.A(_03907_),
    .Y(_04033_));
 sky130_fd_sc_hd__nor2_1 _09904_ (.A(_04032_),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__inv_2 _09905_ (.A(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_1 _09906_ (.A(_04031_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__nand3_1 _09907_ (.A(_04028_),
    .B(_04034_),
    .C(_04030_),
    .Y(_04037_));
 sky130_fd_sc_hd__nand2_1 _09908_ (.A(_04036_),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__inv_2 _09909_ (.A(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_1 _09910_ (.A(_02687_),
    .B(_00421_),
    .Y(_04041_));
 sky130_fd_sc_hd__nand2_1 _09911_ (.A(_05096_),
    .B(_00685_),
    .Y(_04042_));
 sky130_fd_sc_hd__or3_1 _09912_ (.A(_02376_),
    .B(_03219_),
    .C(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__o21ai_1 _09913_ (.A1(_02376_),
    .A2(_03219_),
    .B1(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__nand2_1 _09914_ (.A(_04043_),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__or2_1 _09915_ (.A(_04041_),
    .B(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__nand2_1 _09916_ (.A(_04045_),
    .B(_04041_),
    .Y(_04047_));
 sky130_fd_sc_hd__nand2_1 _09917_ (.A(_04046_),
    .B(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__nand2_1 _09918_ (.A(_03694_),
    .B(_03691_),
    .Y(_04049_));
 sky130_fd_sc_hd__inv_2 _09919_ (.A(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__or2_1 _09920_ (.A(_04048_),
    .B(_04050_),
    .X(_04052_));
 sky130_fd_sc_hd__nand2_1 _09921_ (.A(_04050_),
    .B(_04048_),
    .Y(_04053_));
 sky130_fd_sc_hd__nand2_1 _09922_ (.A(_04645_),
    .B(_00520_),
    .Y(_04054_));
 sky130_fd_sc_hd__inv_2 _09923_ (.A(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__and4_1 _09924_ (.A(_03248_),
    .B(_05114_),
    .C(_00311_),
    .D(_00355_),
    .X(_04056_));
 sky130_fd_sc_hd__a22o_1 _09925_ (.A1(_03248_),
    .A2(_00355_),
    .B1(_05114_),
    .B2(_00311_),
    .X(_04057_));
 sky130_fd_sc_hd__or2b_1 _09926_ (.A(_04056_),
    .B_N(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__xor2_1 _09927_ (.A(_04055_),
    .B(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__inv_2 _09928_ (.A(_04059_),
    .Y(_04060_));
 sky130_fd_sc_hd__a21o_1 _09929_ (.A1(_04052_),
    .A2(_04053_),
    .B1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__nand3_1 _09930_ (.A(_04052_),
    .B(_04060_),
    .C(_04053_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2_1 _09931_ (.A(_04061_),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__nand2_1 _09932_ (.A(_03763_),
    .B(_03759_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand2_1 _09933_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__inv_2 _09934_ (.A(_04065_),
    .Y(_04067_));
 sky130_fd_sc_hd__nand3_1 _09935_ (.A(_04061_),
    .B(_04063_),
    .C(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__nand2_1 _09936_ (.A(_03709_),
    .B(_03698_),
    .Y(_04069_));
 sky130_fd_sc_hd__a21bo_1 _09937_ (.A1(_04066_),
    .A2(_04068_),
    .B1_N(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__nand3b_1 _09938_ (.A_N(_04069_),
    .B(_04066_),
    .C(_04068_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_1 _09939_ (.A(_04070_),
    .B(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__inv_2 _09940_ (.A(_04072_),
    .Y(_04074_));
 sky130_fd_sc_hd__nand2_1 _09941_ (.A(_00433_),
    .B(net22),
    .Y(_04075_));
 sky130_fd_sc_hd__inv_2 _09942_ (.A(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__nand2_1 _09943_ (.A(_00232_),
    .B(net21),
    .Y(_04077_));
 sky130_fd_sc_hd__nand2_1 _09944_ (.A(_00234_),
    .B(net20),
    .Y(_04078_));
 sky130_fd_sc_hd__xor2_1 _09945_ (.A(_04077_),
    .B(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__or2_1 _09946_ (.A(_04076_),
    .B(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__nand2_1 _09947_ (.A(_04079_),
    .B(_04076_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand2_1 _09948_ (.A(_04080_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__a31o_1 _09949_ (.A1(_03725_),
    .A2(_00433_),
    .A3(net21),
    .B1(_03724_),
    .X(_04083_));
 sky130_fd_sc_hd__inv_2 _09950_ (.A(_04083_),
    .Y(_04085_));
 sky130_fd_sc_hd__or2_1 _09951_ (.A(_04082_),
    .B(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__nand2_1 _09952_ (.A(_04085_),
    .B(_04082_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand2_1 _09953_ (.A(_00306_),
    .B(net18),
    .Y(_04088_));
 sky130_fd_sc_hd__and4_1 _09954_ (.A(_00303_),
    .B(_00301_),
    .C(net19),
    .D(net24),
    .X(_04089_));
 sky130_fd_sc_hd__inv_2 _09955_ (.A(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__a22o_1 _09956_ (.A1(_00303_),
    .A2(net24),
    .B1(_00301_),
    .B2(net19),
    .X(_04091_));
 sky130_fd_sc_hd__nand2_1 _09957_ (.A(_04090_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__xnor2_1 _09958_ (.A(_04088_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__inv_2 _09959_ (.A(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__a21o_1 _09960_ (.A1(_04086_),
    .A2(_04087_),
    .B1(_04094_),
    .X(_04096_));
 sky130_fd_sc_hd__nand3_1 _09961_ (.A(_04086_),
    .B(_04094_),
    .C(_04087_),
    .Y(_04097_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(_04096_),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__and2_1 _09963_ (.A(_03741_),
    .B(_03731_),
    .X(_04099_));
 sky130_fd_sc_hd__nor2_1 _09964_ (.A(_04098_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__inv_2 _09965_ (.A(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_1 _09966_ (.A(_04099_),
    .B(_04098_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand2_1 _09967_ (.A(_04101_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__nand2_1 _09968_ (.A(_02203_),
    .B(_05049_),
    .Y(_04104_));
 sky130_fd_sc_hd__inv_2 _09969_ (.A(net17),
    .Y(_04105_));
 sky130_fd_sc_hd__nand2_1 _09970_ (.A(_00315_),
    .B(_00526_),
    .Y(_04107_));
 sky130_fd_sc_hd__nor3_1 _09971_ (.A(_00560_),
    .B(_04105_),
    .C(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__inv_2 _09972_ (.A(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__o21ai_1 _09973_ (.A1(_00560_),
    .A2(_04105_),
    .B1(_04107_),
    .Y(_04110_));
 sky130_fd_sc_hd__nand2_1 _09974_ (.A(_04109_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__or2_1 _09975_ (.A(_04104_),
    .B(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__nand2_1 _09976_ (.A(_04111_),
    .B(_04104_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand2_1 _09977_ (.A(_04112_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__o21a_1 _09978_ (.A1(_03734_),
    .A2(_03738_),
    .B1(_03736_),
    .X(_04115_));
 sky130_fd_sc_hd__nor2_1 _09979_ (.A(_04114_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__inv_2 _09980_ (.A(_04116_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand2_1 _09981_ (.A(_04115_),
    .B(_04114_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _09982_ (.A(_03755_),
    .B(_03751_),
    .Y(_04120_));
 sky130_fd_sc_hd__a21o_1 _09983_ (.A1(_04118_),
    .A2(_04119_),
    .B1(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__nand3_1 _09984_ (.A(_04118_),
    .B(_04120_),
    .C(_04119_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _09985_ (.A(_04121_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_1 _09986_ (.A(_04103_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__inv_2 _09987_ (.A(_04123_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand3_1 _09988_ (.A(_04101_),
    .B(_04125_),
    .C(_04102_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_1 _09989_ (.A(_04124_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__nand2_1 _09990_ (.A(_03767_),
    .B(_03746_),
    .Y(_04129_));
 sky130_fd_sc_hd__inv_2 _09991_ (.A(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _09992_ (.A(_04127_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__nand3_1 _09993_ (.A(_04124_),
    .B(_04129_),
    .C(_04126_),
    .Y(_04132_));
 sky130_fd_sc_hd__nand3_1 _09994_ (.A(_04074_),
    .B(_04131_),
    .C(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand2_1 _09995_ (.A(_04131_),
    .B(_04132_),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_04134_),
    .B(_04072_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand2_1 _09997_ (.A(_04133_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__nand2_1 _09998_ (.A(_03772_),
    .B(_03768_),
    .Y(_04137_));
 sky130_fd_sc_hd__inv_2 _09999_ (.A(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand2_1 _10000_ (.A(_04136_),
    .B(_04138_),
    .Y(_04140_));
 sky130_fd_sc_hd__nand3_1 _10001_ (.A(_04137_),
    .B(_04133_),
    .C(_04135_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_1 _10002_ (.A(_04140_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand2_1 _10003_ (.A(_03790_),
    .B(_03786_),
    .Y(_04143_));
 sky130_fd_sc_hd__nand2_1 _10004_ (.A(_02214_),
    .B(_04888_),
    .Y(_04144_));
 sky130_fd_sc_hd__inv_2 _10005_ (.A(_04899_),
    .Y(_04145_));
 sky130_fd_sc_hd__or4_1 _10006_ (.A(_02650_),
    .B(_02377_),
    .C(_00188_),
    .D(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__a22o_1 _10007_ (.A1(_04128_),
    .A2(_04899_),
    .B1(_00960_),
    .B2(_04897_),
    .X(_04147_));
 sky130_fd_sc_hd__nand2_1 _10008_ (.A(_04146_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__or2_1 _10009_ (.A(_04144_),
    .B(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__nand2_1 _10010_ (.A(_04148_),
    .B(_04144_),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_1 _10011_ (.A(_04149_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__inv_2 _10012_ (.A(_03705_),
    .Y(_04153_));
 sky130_fd_sc_hd__o21a_1 _10013_ (.A1(_03702_),
    .A2(_04153_),
    .B1(_03704_),
    .X(_04154_));
 sky130_fd_sc_hd__inv_2 _10014_ (.A(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand2_1 _10015_ (.A(_04152_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand3_1 _10016_ (.A(_04149_),
    .B(_04154_),
    .C(_04151_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand3b_1 _10017_ (.A_N(_04143_),
    .B(_04156_),
    .C(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__nand2_1 _10018_ (.A(_04152_),
    .B(_04154_),
    .Y(_04159_));
 sky130_fd_sc_hd__nand3_1 _10019_ (.A(_04149_),
    .B(_04151_),
    .C(_04155_),
    .Y(_04160_));
 sky130_fd_sc_hd__nand3_1 _10020_ (.A(_04159_),
    .B(_04143_),
    .C(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__nand2_1 _10021_ (.A(_04158_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__nand2_1 _10022_ (.A(_03799_),
    .B(_03794_),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2_1 _10023_ (.A(_04163_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__inv_2 _10024_ (.A(_04164_),
    .Y(_04166_));
 sky130_fd_sc_hd__nand3_1 _10025_ (.A(_04158_),
    .B(_04162_),
    .C(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand2_1 _10026_ (.A(_04165_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__or4_1 _10027_ (.A(_03289_),
    .B(_02437_),
    .C(_05179_),
    .D(_03807_),
    .X(_04169_));
 sky130_fd_sc_hd__a22o_1 _10028_ (.A1(_01532_),
    .A2(_04933_),
    .B1(_01334_),
    .B2(_04936_),
    .X(_04170_));
 sky130_fd_sc_hd__nand2_1 _10029_ (.A(_04169_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand3b_1 _10030_ (.A_N(_04171_),
    .B(_03105_),
    .C(_04941_),
    .Y(_04173_));
 sky130_fd_sc_hd__nand2_1 _10031_ (.A(_03105_),
    .B(_04941_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand2_1 _10032_ (.A(_04171_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_04173_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__inv_2 _10034_ (.A(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_1 _10035_ (.A(_03812_),
    .B(_03808_),
    .Y(_04178_));
 sky130_fd_sc_hd__nand2_1 _10036_ (.A(_04177_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__inv_2 _10037_ (.A(_04178_),
    .Y(_04180_));
 sky130_fd_sc_hd__nand2_1 _10038_ (.A(_04180_),
    .B(_04176_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand2_1 _10039_ (.A(_04179_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2_1 _10040_ (.A(_00682_),
    .B(_00138_),
    .Y(_04184_));
 sky130_fd_sc_hd__inv_2 _10041_ (.A(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__and4_1 _10042_ (.A(net46),
    .B(_05191_),
    .C(_05113_),
    .D(_05278_),
    .X(_04186_));
 sky130_fd_sc_hd__a22o_1 _10043_ (.A1(net46),
    .A2(_05113_),
    .B1(_05191_),
    .B2(_05278_),
    .X(_04187_));
 sky130_fd_sc_hd__or2b_1 _10044_ (.A(_04186_),
    .B_N(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__xor2_1 _10045_ (.A(_04185_),
    .B(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__nand2_1 _10046_ (.A(_04182_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__inv_2 _10047_ (.A(_04189_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand3_1 _10048_ (.A(_04179_),
    .B(_04191_),
    .C(_04181_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand2_1 _10049_ (.A(_04190_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__inv_2 _10050_ (.A(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _10051_ (.A(_04168_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand3_1 _10052_ (.A(_04193_),
    .B(_04165_),
    .C(_04167_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _10053_ (.A(_04196_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__a21oi_1 _10054_ (.A1(_03714_),
    .A2(_03716_),
    .B1(_03713_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _10055_ (.A(_04198_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__inv_2 _10056_ (.A(_04199_),
    .Y(_04201_));
 sky130_fd_sc_hd__nand3_1 _10057_ (.A(_04196_),
    .B(_04197_),
    .C(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__nand2_1 _10058_ (.A(_04200_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__nor2_1 _10059_ (.A(_03800_),
    .B(_03802_),
    .Y(_04204_));
 sky130_fd_sc_hd__inv_2 _10060_ (.A(_03833_),
    .Y(_04206_));
 sky130_fd_sc_hd__nor2_1 _10061_ (.A(_04204_),
    .B(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_1 _10062_ (.A(_04203_),
    .B(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__inv_2 _10063_ (.A(_04207_),
    .Y(_04209_));
 sky130_fd_sc_hd__nand3_1 _10064_ (.A(_04209_),
    .B(_04200_),
    .C(_04202_),
    .Y(_04210_));
 sky130_fd_sc_hd__nand2_1 _10065_ (.A(_04208_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2_1 _10066_ (.A(_04142_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__inv_2 _10067_ (.A(_04211_),
    .Y(_04213_));
 sky130_fd_sc_hd__nand3_1 _10068_ (.A(_04140_),
    .B(_04213_),
    .C(_04141_),
    .Y(_04214_));
 sky130_fd_sc_hd__nand2_1 _10069_ (.A(_04212_),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__nand2_1 _10070_ (.A(_03850_),
    .B(_03780_),
    .Y(_04217_));
 sky130_fd_sc_hd__inv_2 _10071_ (.A(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__nand2_1 _10072_ (.A(_04215_),
    .B(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__nand3_1 _10073_ (.A(_04217_),
    .B(_04212_),
    .C(_04214_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand3_1 _10074_ (.A(_04039_),
    .B(_04219_),
    .C(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__nand2_1 _10075_ (.A(_04219_),
    .B(_04220_),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_1 _10076_ (.A(_04222_),
    .B(_04038_),
    .Y(_04223_));
 sky130_fd_sc_hd__nand2_1 _10077_ (.A(_04221_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__nor2_1 _10078_ (.A(_03960_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__inv_2 _10079_ (.A(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__nand2_1 _10080_ (.A(_04224_),
    .B(_03960_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand2_1 _10081_ (.A(_04226_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nor2_1 _10082_ (.A(_03913_),
    .B(_03910_),
    .Y(_04230_));
 sky130_fd_sc_hd__inv_2 _10083_ (.A(_03923_),
    .Y(_04231_));
 sky130_fd_sc_hd__nor2_1 _10084_ (.A(_04230_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_1 _10085_ (.A(_04229_),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__inv_2 _10086_ (.A(_04232_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand3_2 _10087_ (.A(_04226_),
    .B(_04234_),
    .C(_04228_),
    .Y(_04235_));
 sky130_fd_sc_hd__nand3b_4 _10088_ (.A_N(_03958_),
    .B(_04233_),
    .C(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__nand2_1 _10089_ (.A(_04233_),
    .B(_04235_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_2 _10090_ (.A(_04237_),
    .B(_03958_),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_1 _10091_ (.A(_04236_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_1 _10092_ (.A(_04240_),
    .B(_03946_),
    .Y(_04241_));
 sky130_fd_sc_hd__nand3b_1 _10093_ (.A_N(_03946_),
    .B(_04236_),
    .C(_04239_),
    .Y(_04242_));
 sky130_fd_sc_hd__nand2_1 _10094_ (.A(_04241_),
    .B(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__inv_2 _10095_ (.A(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_1 _10096_ (.A(_03957_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2_1 _10097_ (.A(_04245_),
    .B(_04242_),
    .Y(_04246_));
 sky130_fd_sc_hd__a21boi_1 _10098_ (.A1(_04039_),
    .A2(_04219_),
    .B1_N(_04220_),
    .Y(_04247_));
 sky130_fd_sc_hd__inv_2 _10099_ (.A(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__nand2_1 _10100_ (.A(_04097_),
    .B(_04086_),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2_1 _10101_ (.A(_00306_),
    .B(net19),
    .Y(_04251_));
 sky130_fd_sc_hd__inv_2 _10102_ (.A(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__and4_1 _10103_ (.A(_00303_),
    .B(_00301_),
    .C(net20),
    .D(net25),
    .X(_04253_));
 sky130_fd_sc_hd__a22o_1 _10104_ (.A1(_00303_),
    .A2(net25),
    .B1(_00301_),
    .B2(net20),
    .X(_04254_));
 sky130_fd_sc_hd__or2b_1 _10105_ (.A(_04253_),
    .B_N(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__xor2_1 _10106_ (.A(_04252_),
    .B(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__inv_2 _10107_ (.A(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__and4_1 _10108_ (.A(_00234_),
    .B(_00232_),
    .C(net20),
    .D(net21),
    .X(_04258_));
 sky130_fd_sc_hd__inv_2 _10109_ (.A(_04081_),
    .Y(_04259_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(_04258_),
    .B(_04259_),
    .Y(_04261_));
 sky130_fd_sc_hd__inv_2 _10111_ (.A(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__nand2_1 _10112_ (.A(_00234_),
    .B(net21),
    .Y(_04263_));
 sky130_fd_sc_hd__or3b_1 _10113_ (.A(_02312_),
    .B(_04263_),
    .C_N(net22),
    .X(_04264_));
 sky130_fd_sc_hd__a21bo_1 _10114_ (.A1(_00232_),
    .A2(net22),
    .B1_N(_04263_),
    .X(_04265_));
 sky130_fd_sc_hd__nand2_1 _10115_ (.A(_00433_),
    .B(net24),
    .Y(_04266_));
 sky130_fd_sc_hd__a21bo_1 _10116_ (.A1(_04264_),
    .A2(_04265_),
    .B1_N(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__nand3b_1 _10117_ (.A_N(_04266_),
    .B(_04264_),
    .C(_04265_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_1 _10118_ (.A(_04267_),
    .B(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__or2_1 _10119_ (.A(_04262_),
    .B(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__nand2_1 _10120_ (.A(_04269_),
    .B(_04262_),
    .Y(_04272_));
 sky130_fd_sc_hd__nand2_1 _10121_ (.A(_04270_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__or2_1 _10122_ (.A(_04257_),
    .B(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__nand2_1 _10123_ (.A(_04273_),
    .B(_04257_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand2_1 _10124_ (.A(_04274_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__nor2_1 _10125_ (.A(_04250_),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__and2_1 _10126_ (.A(_04276_),
    .B(_04250_),
    .X(_04278_));
 sky130_fd_sc_hd__nand2_1 _10127_ (.A(_04112_),
    .B(_04109_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _10128_ (.A(_02203_),
    .B(_00526_),
    .Y(_04280_));
 sky130_fd_sc_hd__nand2_1 _10129_ (.A(_00315_),
    .B(net17),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(_05068_),
    .B(net18),
    .Y(_04283_));
 sky130_fd_sc_hd__xnor2_1 _10131_ (.A(_04281_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__xnor2_1 _10132_ (.A(_04280_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__o21a_1 _10133_ (.A1(_04088_),
    .A2(_04092_),
    .B1(_04090_),
    .X(_04286_));
 sky130_fd_sc_hd__xor2_1 _10134_ (.A(_04285_),
    .B(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__or2_1 _10135_ (.A(_04279_),
    .B(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__nand2_1 _10136_ (.A(_04287_),
    .B(_04279_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_1 _10137_ (.A(_04288_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__o21bai_1 _10138_ (.A1(_04277_),
    .A2(_04278_),
    .B1_N(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__or2_1 _10139_ (.A(_04250_),
    .B(_04276_),
    .X(_04292_));
 sky130_fd_sc_hd__nand2_1 _10140_ (.A(_04276_),
    .B(_04250_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand3_1 _10141_ (.A(_04292_),
    .B(_04290_),
    .C(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_1 _10142_ (.A(_04291_),
    .B(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__a21oi_1 _10143_ (.A1(_04102_),
    .A2(_04125_),
    .B1(_04100_),
    .Y(_04297_));
 sky130_fd_sc_hd__inv_2 _10144_ (.A(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__nand2_1 _10145_ (.A(_04296_),
    .B(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__nand3_1 _10146_ (.A(_04291_),
    .B(_04295_),
    .C(_04297_),
    .Y(_04300_));
 sky130_fd_sc_hd__nand2_1 _10147_ (.A(_04299_),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand2_1 _10148_ (.A(_04645_),
    .B(_00311_),
    .Y(_04302_));
 sky130_fd_sc_hd__inv_2 _10149_ (.A(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__nand2_1 _10150_ (.A(_05114_),
    .B(_00355_),
    .Y(_04305_));
 sky130_fd_sc_hd__nand2_1 _10151_ (.A(_03248_),
    .B(_00421_),
    .Y(_04306_));
 sky130_fd_sc_hd__xnor2_1 _10152_ (.A(_04305_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__xor2_1 _10153_ (.A(_04303_),
    .B(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__inv_2 _10154_ (.A(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__and2_1 _10155_ (.A(_04046_),
    .B(_04043_),
    .X(_04310_));
 sky130_fd_sc_hd__nand2_1 _10156_ (.A(_02687_),
    .B(_00685_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand2_1 _10157_ (.A(_05096_),
    .B(_01895_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand2_1 _10158_ (.A(_03039_),
    .B(_05049_),
    .Y(_04313_));
 sky130_fd_sc_hd__xnor2_1 _10159_ (.A(_04312_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__xnor2_1 _10160_ (.A(_04311_),
    .B(_04314_),
    .Y(_04316_));
 sky130_fd_sc_hd__or2b_1 _10161_ (.A(_04310_),
    .B_N(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__or2b_1 _10162_ (.A(_04316_),
    .B_N(_04310_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _10163_ (.A(_04317_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__or2_1 _10164_ (.A(_04309_),
    .B(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__nand2_1 _10165_ (.A(_04319_),
    .B(_04309_),
    .Y(_04321_));
 sky130_fd_sc_hd__nand2_1 _10166_ (.A(_04122_),
    .B(_04118_),
    .Y(_04322_));
 sky130_fd_sc_hd__a21bo_1 _10167_ (.A1(_04320_),
    .A2(_04321_),
    .B1_N(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__nand3b_1 _10168_ (.A_N(_04322_),
    .B(_04320_),
    .C(_04321_),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _10169_ (.A(_04323_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__nand2_1 _10170_ (.A(_04063_),
    .B(_04052_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand2_1 _10171_ (.A(_04325_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__nand3b_1 _10172_ (.A_N(_04327_),
    .B(_04323_),
    .C(_04324_),
    .Y(_04329_));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(_04328_),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__inv_2 _10174_ (.A(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__nand2_1 _10175_ (.A(_04301_),
    .B(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand3_1 _10176_ (.A(_04299_),
    .B(_04330_),
    .C(_04300_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand2_1 _10177_ (.A(_04332_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__a21boi_1 _10178_ (.A1(_04074_),
    .A2(_04131_),
    .B1_N(_04132_),
    .Y(_04335_));
 sky130_fd_sc_hd__inv_2 _10179_ (.A(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(_04334_),
    .B(_04336_),
    .Y(_04338_));
 sky130_fd_sc_hd__nand3_1 _10181_ (.A(_04335_),
    .B(_04332_),
    .C(_04333_),
    .Y(_04339_));
 sky130_fd_sc_hd__nand2_1 _10182_ (.A(_04338_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__nand2_1 _10183_ (.A(_04162_),
    .B(_04160_),
    .Y(_04341_));
 sky130_fd_sc_hd__nand2_1 _10184_ (.A(_04149_),
    .B(_04146_),
    .Y(_04342_));
 sky130_fd_sc_hd__a21oi_1 _10185_ (.A1(_04057_),
    .A2(_04055_),
    .B1(_04056_),
    .Y(_04343_));
 sky130_fd_sc_hd__inv_2 _10186_ (.A(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__nand2_1 _10187_ (.A(_04128_),
    .B(_04888_),
    .Y(_04345_));
 sky130_fd_sc_hd__or4_1 _10188_ (.A(_02377_),
    .B(_00188_),
    .C(_02385_),
    .D(_04145_),
    .X(_04346_));
 sky130_fd_sc_hd__a22o_1 _10189_ (.A1(_00960_),
    .A2(_04899_),
    .B1(_04897_),
    .B2(_00520_),
    .X(_04347_));
 sky130_fd_sc_hd__nand2_1 _10190_ (.A(_04346_),
    .B(_04347_),
    .Y(_04349_));
 sky130_fd_sc_hd__xnor2_1 _10191_ (.A(_04345_),
    .B(_04349_),
    .Y(_04350_));
 sky130_fd_sc_hd__or2_1 _10192_ (.A(_04344_),
    .B(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__nand2_1 _10193_ (.A(_04350_),
    .B(_04344_),
    .Y(_04352_));
 sky130_fd_sc_hd__nand3b_1 _10194_ (.A_N(_04342_),
    .B(_04351_),
    .C(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__nand2_1 _10195_ (.A(_04351_),
    .B(_04352_),
    .Y(_04354_));
 sky130_fd_sc_hd__nand2_1 _10196_ (.A(_04354_),
    .B(_04342_),
    .Y(_04355_));
 sky130_fd_sc_hd__nand3b_1 _10197_ (.A_N(_04341_),
    .B(_04353_),
    .C(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__nand2_1 _10198_ (.A(_04355_),
    .B(_04353_),
    .Y(_04357_));
 sky130_fd_sc_hd__nand2_1 _10199_ (.A(_04357_),
    .B(_04341_),
    .Y(_04358_));
 sky130_fd_sc_hd__nand2_1 _10200_ (.A(_04356_),
    .B(_04358_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand2_1 _10201_ (.A(_01532_),
    .B(_04941_),
    .Y(_04361_));
 sky130_fd_sc_hd__or4_1 _10202_ (.A(_02437_),
    .B(_02369_),
    .C(_05179_),
    .D(_03807_),
    .X(_04362_));
 sky130_fd_sc_hd__a22o_1 _10203_ (.A1(_01334_),
    .A2(_04933_),
    .B1(_02214_),
    .B2(_04936_),
    .X(_04363_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(_04362_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__xnor2_1 _10205_ (.A(_04361_),
    .B(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__nand2_1 _10206_ (.A(_04173_),
    .B(_04169_),
    .Y(_04366_));
 sky130_fd_sc_hd__nor2_1 _10207_ (.A(_04365_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__inv_2 _10208_ (.A(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__nand2_1 _10209_ (.A(_04366_),
    .B(_04365_),
    .Y(_04369_));
 sky130_fd_sc_hd__nand2_1 _10210_ (.A(_00682_),
    .B(_05278_),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_1 _10211_ (.A(_05191_),
    .B(_05113_),
    .Y(_04372_));
 sky130_fd_sc_hd__nand2_1 _10212_ (.A(net46),
    .B(_03105_),
    .Y(_04373_));
 sky130_fd_sc_hd__xnor2_1 _10213_ (.A(_04372_),
    .B(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__xnor2_1 _10214_ (.A(_04371_),
    .B(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__a21o_1 _10215_ (.A1(_04368_),
    .A2(_04369_),
    .B1(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__nand3b_1 _10216_ (.A_N(_04367_),
    .B(_04375_),
    .C(_04369_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand2_1 _10217_ (.A(_04376_),
    .B(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__inv_2 _10218_ (.A(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__nand2_1 _10219_ (.A(_04360_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand3_1 _10220_ (.A(_04356_),
    .B(_04378_),
    .C(_04358_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_1 _10221_ (.A(_04380_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__nand2_1 _10222_ (.A(_04064_),
    .B(_04067_),
    .Y(_04384_));
 sky130_fd_sc_hd__nor2_1 _10223_ (.A(_04067_),
    .B(_04064_),
    .Y(_04385_));
 sky130_fd_sc_hd__a21oi_1 _10224_ (.A1(_04384_),
    .A2(_04069_),
    .B1(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__inv_2 _10225_ (.A(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__nand2_1 _10226_ (.A(_04383_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__nand3_1 _10227_ (.A(_04380_),
    .B(_04382_),
    .C(_04386_),
    .Y(_04389_));
 sky130_fd_sc_hd__nand2_1 _10228_ (.A(_04388_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nor2_1 _10229_ (.A(_04166_),
    .B(_04163_),
    .Y(_04391_));
 sky130_fd_sc_hd__inv_2 _10230_ (.A(_04196_),
    .Y(_04393_));
 sky130_fd_sc_hd__nor2_1 _10231_ (.A(_04391_),
    .B(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__inv_2 _10232_ (.A(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2_1 _10233_ (.A(_04390_),
    .B(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__nand3_1 _10234_ (.A(_04388_),
    .B(_04389_),
    .C(_04394_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _10235_ (.A(_04396_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__inv_2 _10236_ (.A(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2_1 _10237_ (.A(_04340_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand3_1 _10238_ (.A(_04398_),
    .B(_04338_),
    .C(_04339_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _10239_ (.A(_04400_),
    .B(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__a21boi_1 _10240_ (.A1(_04140_),
    .A2(_04213_),
    .B1_N(_04141_),
    .Y(_04404_));
 sky130_fd_sc_hd__inv_2 _10241_ (.A(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__nand2_1 _10242_ (.A(_04402_),
    .B(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__nand3_1 _10243_ (.A(_04404_),
    .B(_04400_),
    .C(_04401_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand2_1 _10244_ (.A(_04406_),
    .B(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21oi_1 _10245_ (.A1(_04187_),
    .A2(_04185_),
    .B1(_04186_),
    .Y(_04409_));
 sky130_fd_sc_hd__inv_2 _10246_ (.A(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nand2_1 _10247_ (.A(net51),
    .B(_05159_),
    .Y(_04411_));
 sky130_fd_sc_hd__or4_1 _10248_ (.A(_03148_),
    .B(_02728_),
    .C(_03965_),
    .D(_02802_),
    .X(_04412_));
 sky130_fd_sc_hd__a22o_1 _10249_ (.A1(net49),
    .A2(_00138_),
    .B1(net50),
    .B2(_00329_),
    .X(_04413_));
 sky130_fd_sc_hd__nand2_1 _10250_ (.A(_04412_),
    .B(_04413_),
    .Y(_04415_));
 sky130_fd_sc_hd__xnor2_1 _10251_ (.A(_04411_),
    .B(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__or2_1 _10252_ (.A(_04410_),
    .B(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__nand2_1 _10253_ (.A(_04416_),
    .B(_04410_),
    .Y(_04418_));
 sky130_fd_sc_hd__nand2_1 _10254_ (.A(_04417_),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__nand2_1 _10255_ (.A(_03969_),
    .B(_03966_),
    .Y(_04420_));
 sky130_fd_sc_hd__nand2_1 _10256_ (.A(_04419_),
    .B(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__nand3b_1 _10257_ (.A_N(_04420_),
    .B(_04417_),
    .C(_04418_),
    .Y(_04422_));
 sky130_fd_sc_hd__nand2_1 _10258_ (.A(_04421_),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__nor2_1 _10259_ (.A(_04176_),
    .B(_04180_),
    .Y(_04424_));
 sky130_fd_sc_hd__a21oi_1 _10260_ (.A1(_04181_),
    .A2(_04191_),
    .B1(_04424_),
    .Y(_04426_));
 sky130_fd_sc_hd__inv_2 _10261_ (.A(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_1 _10262_ (.A(_04423_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__nand3_1 _10263_ (.A(_04421_),
    .B(_04426_),
    .C(_04422_),
    .Y(_04429_));
 sky130_fd_sc_hd__nand2_1 _10264_ (.A(_04428_),
    .B(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__nand2_1 _10265_ (.A(_03980_),
    .B(_03979_),
    .Y(_04431_));
 sky130_fd_sc_hd__nand2_1 _10266_ (.A(_04430_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__nand3b_1 _10267_ (.A_N(_04431_),
    .B(_04428_),
    .C(_04429_),
    .Y(_04433_));
 sky130_fd_sc_hd__nand2_1 _10268_ (.A(_04432_),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__a21oi_1 _10269_ (.A1(_03986_),
    .A2(_03984_),
    .B1(_03982_),
    .Y(_04435_));
 sky130_fd_sc_hd__inv_2 _10270_ (.A(_04435_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _10271_ (.A(_04434_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__nand3_1 _10272_ (.A(_04432_),
    .B(_04433_),
    .C(_04435_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_1 _10273_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__nor2_1 _10274_ (.A(_03999_),
    .B(_04012_),
    .Y(_04441_));
 sky130_fd_sc_hd__nand2_1 _10275_ (.A(net54),
    .B(_00381_),
    .Y(_04442_));
 sky130_fd_sc_hd__or4_1 _10276_ (.A(_03643_),
    .B(_05178_),
    .C(_03645_),
    .D(_02875_),
    .X(_04443_));
 sky130_fd_sc_hd__a22o_1 _10277_ (.A1(net52),
    .A2(_00893_),
    .B1(net53),
    .B2(_00384_),
    .X(_04444_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(_04443_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__xnor2_1 _10279_ (.A(_04442_),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__nand2_1 _10280_ (.A(_04005_),
    .B(_04002_),
    .Y(_04448_));
 sky130_fd_sc_hd__or2_1 _10281_ (.A(_04446_),
    .B(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(_04448_),
    .B(_04446_),
    .Y(_04450_));
 sky130_fd_sc_hd__nand2_1 _10283_ (.A(_04449_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__nand2_1 _10284_ (.A(net56),
    .B(_05310_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_1 _10285_ (.A(_04451_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand3b_1 _10286_ (.A_N(_04452_),
    .B(_04449_),
    .C(_04450_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _10287_ (.A(_04453_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__o21ai_1 _10288_ (.A1(_04009_),
    .A2(_04441_),
    .B1(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__a31oi_1 _10289_ (.A1(_04011_),
    .A2(net56),
    .A3(_00194_),
    .B1(_04009_),
    .Y(_04457_));
 sky130_fd_sc_hd__nand3_1 _10290_ (.A(_04457_),
    .B(_04454_),
    .C(_04453_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(_04456_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_1 _10292_ (.A(net57),
    .B(_00194_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(_04460_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand3b_1 _10294_ (.A_N(_04461_),
    .B(_04456_),
    .C(_04459_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_1 _10295_ (.A(_04462_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__inv_2 _10296_ (.A(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__nand2_1 _10297_ (.A(_04440_),
    .B(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__nand3_1 _10298_ (.A(_04464_),
    .B(_04438_),
    .C(_04439_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _10299_ (.A(_04466_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand2_1 _10300_ (.A(_04210_),
    .B(_04202_),
    .Y(_04470_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(_04468_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__inv_2 _10302_ (.A(_04470_),
    .Y(_04472_));
 sky130_fd_sc_hd__nand3_1 _10303_ (.A(_04472_),
    .B(_04466_),
    .C(_04467_),
    .Y(_04473_));
 sky130_fd_sc_hd__nand2_1 _10304_ (.A(_04471_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__nor2_1 _10305_ (.A(_03993_),
    .B(_03992_),
    .Y(_04475_));
 sky130_fd_sc_hd__inv_2 _10306_ (.A(_04021_),
    .Y(_04476_));
 sky130_fd_sc_hd__nor2_1 _10307_ (.A(_04475_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__inv_2 _10308_ (.A(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__nand2_1 _10309_ (.A(_04474_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__nand3_1 _10310_ (.A(_04471_),
    .B(_04473_),
    .C(_04477_),
    .Y(_04481_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(_04479_),
    .B(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__inv_2 _10312_ (.A(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _10313_ (.A(_04408_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__nand3_1 _10314_ (.A(_04406_),
    .B(_04482_),
    .C(_04407_),
    .Y(_04485_));
 sky130_fd_sc_hd__nand2_1 _10315_ (.A(_04484_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__nand2_1 _10316_ (.A(_04248_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__nand3_1 _10317_ (.A(_04247_),
    .B(_04485_),
    .C(_04484_),
    .Y(_04488_));
 sky130_fd_sc_hd__nand2_1 _10318_ (.A(_04487_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__nor2_1 _10319_ (.A(_04026_),
    .B(_04023_),
    .Y(_04490_));
 sky130_fd_sc_hd__inv_2 _10320_ (.A(_04036_),
    .Y(_04492_));
 sky130_fd_sc_hd__nor2_1 _10321_ (.A(_04490_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__inv_2 _10322_ (.A(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__nand2_1 _10323_ (.A(_04489_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__nand3_1 _10324_ (.A(_04487_),
    .B(_04488_),
    .C(_04493_),
    .Y(_04496_));
 sky130_fd_sc_hd__nand2_1 _10325_ (.A(_04495_),
    .B(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__a21oi_1 _10326_ (.A1(_04228_),
    .A2(_04234_),
    .B1(_04225_),
    .Y(_04498_));
 sky130_fd_sc_hd__inv_2 _10327_ (.A(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__nand2_1 _10328_ (.A(_04497_),
    .B(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__nand3_1 _10329_ (.A(_04495_),
    .B(_04498_),
    .C(_04496_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand2_1 _10330_ (.A(_04500_),
    .B(_04501_),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_1 _10331_ (.A(_04503_),
    .B(_04017_),
    .Y(_04504_));
 sky130_fd_sc_hd__nand3b_1 _10332_ (.A_N(_04017_),
    .B(_04500_),
    .C(_04501_),
    .Y(_04505_));
 sky130_fd_sc_hd__nand2_1 _10333_ (.A(_04504_),
    .B(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__nand2_1 _10334_ (.A(_04506_),
    .B(_04236_),
    .Y(_04507_));
 sky130_fd_sc_hd__nand3b_1 _10335_ (.A_N(_04236_),
    .B(_04504_),
    .C(_04505_),
    .Y(_04508_));
 sky130_fd_sc_hd__nand2_2 _10336_ (.A(_04507_),
    .B(_04508_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _10337_ (.A(_04246_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__inv_2 _10338_ (.A(_04509_),
    .Y(_04511_));
 sky130_fd_sc_hd__nand3_1 _10339_ (.A(_04245_),
    .B(_04511_),
    .C(_04242_),
    .Y(_04512_));
 sky130_fd_sc_hd__nand2_1 _10340_ (.A(_04510_),
    .B(_04512_),
    .Y(_04514_));
 sky130_fd_sc_hd__inv_2 _10341_ (.A(net151),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _10342_ (.A(_04514_),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__nand3_1 _10343_ (.A(_04510_),
    .B(net151),
    .C(_04512_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand2_1 _10344_ (.A(_04516_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__inv_2 _10345_ (.A(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__inv_2 _10346_ (.A(_03687_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _10347_ (.A(_03434_),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand3_1 _10348_ (.A(_03422_),
    .B(_03433_),
    .C(_03687_),
    .Y(_04522_));
 sky130_fd_sc_hd__nand3_1 _10349_ (.A(_04521_),
    .B(_04522_),
    .C(net160),
    .Y(_04523_));
 sky130_fd_sc_hd__nand2_1 _10350_ (.A(_04521_),
    .B(_03686_),
    .Y(_04525_));
 sky130_fd_sc_hd__inv_2 _10351_ (.A(_03950_),
    .Y(_04526_));
 sky130_fd_sc_hd__nand2_1 _10352_ (.A(_04525_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand3_1 _10353_ (.A(_04521_),
    .B(_03950_),
    .C(_03686_),
    .Y(_04528_));
 sky130_fd_sc_hd__nand2_1 _10354_ (.A(_04527_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__inv_2 _10355_ (.A(net140),
    .Y(_04530_));
 sky130_fd_sc_hd__and2_1 _10356_ (.A(_04529_),
    .B(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__nand3_1 _10357_ (.A(_04527_),
    .B(net140),
    .C(_04528_),
    .Y(_04532_));
 sky130_fd_sc_hd__o21a_1 _10358_ (.A1(_04523_),
    .A2(_04531_),
    .B1(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__inv_2 _10359_ (.A(_03420_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _10360_ (.A(_02366_),
    .B(_04534_),
    .Y(_04536_));
 sky130_fd_sc_hd__nand2_1 _10361_ (.A(_04536_),
    .B(_03431_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_2 _10362_ (.A(_04537_),
    .B(_03126_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_1 _10363_ (.A(_04538_),
    .B(_03124_),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _10364_ (.A(_04539_),
    .B(_03394_),
    .Y(_04540_));
 sky130_fd_sc_hd__nand3b_1 _10365_ (.A_N(_03394_),
    .B(_04538_),
    .C(_03124_),
    .Y(_04541_));
 sky130_fd_sc_hd__nand2_1 _10366_ (.A(_04540_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__inv_2 _10367_ (.A(net130),
    .Y(_04543_));
 sky130_fd_sc_hd__nand2_1 _10368_ (.A(_04542_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand3_1 _10369_ (.A(_04540_),
    .B(_04541_),
    .C(net130),
    .Y(_04545_));
 sky130_fd_sc_hd__or2_1 _10370_ (.A(_03126_),
    .B(_04537_),
    .X(_04547_));
 sky130_fd_sc_hd__nand3_2 _10371_ (.A(_04547_),
    .B(net153),
    .C(_04538_),
    .Y(_04548_));
 sky130_fd_sc_hd__inv_2 _10372_ (.A(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__nand3_1 _10373_ (.A(_04544_),
    .B(_04545_),
    .C(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand2_1 _10374_ (.A(_04550_),
    .B(_04545_),
    .Y(_04551_));
 sky130_fd_sc_hd__nand2_1 _10375_ (.A(_04529_),
    .B(_04530_),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_1 _10376_ (.A(_04521_),
    .B(_04522_),
    .Y(_04553_));
 sky130_fd_sc_hd__inv_2 _10377_ (.A(net160),
    .Y(_04554_));
 sky130_fd_sc_hd__nand2_1 _10378_ (.A(_04553_),
    .B(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__nand2_1 _10379_ (.A(_04555_),
    .B(_04523_),
    .Y(_04556_));
 sky130_fd_sc_hd__inv_2 _10380_ (.A(_04556_),
    .Y(_04558_));
 sky130_fd_sc_hd__nand3_1 _10381_ (.A(_04552_),
    .B(_04532_),
    .C(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__inv_2 _10382_ (.A(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_1 _10383_ (.A(_04551_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__nand2_1 _10384_ (.A(_04533_),
    .B(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__nand2_1 _10385_ (.A(_02366_),
    .B(_03419_),
    .Y(_04563_));
 sky130_fd_sc_hd__nand3_1 _10386_ (.A(_01789_),
    .B(_02365_),
    .C(_03418_),
    .Y(_04564_));
 sky130_fd_sc_hd__nand3_1 _10387_ (.A(_04563_),
    .B(net127),
    .C(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _10388_ (.A(_04563_),
    .B(_03417_),
    .Y(_04566_));
 sky130_fd_sc_hd__nand2_1 _10389_ (.A(_04566_),
    .B(_03411_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand3b_1 _10390_ (.A_N(_03411_),
    .B(_04563_),
    .C(_03417_),
    .Y(_04569_));
 sky130_fd_sc_hd__nand2_1 _10391_ (.A(_04567_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__inv_2 _10392_ (.A(net72),
    .Y(_04571_));
 sky130_fd_sc_hd__nand2_1 _10393_ (.A(_04570_),
    .B(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand3_1 _10394_ (.A(_04567_),
    .B(_04569_),
    .C(net72),
    .Y(_04573_));
 sky130_fd_sc_hd__nand2_1 _10395_ (.A(_04572_),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__o21ai_1 _10396_ (.A1(_04565_),
    .A2(_04574_),
    .B1(_04573_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21o_1 _10397_ (.A1(_04563_),
    .A2(_04564_),
    .B1(net127),
    .X(_04576_));
 sky130_fd_sc_hd__nand2_1 _10398_ (.A(_04576_),
    .B(_04565_),
    .Y(_04577_));
 sky130_fd_sc_hd__inv_2 _10399_ (.A(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand3_1 _10400_ (.A(_04578_),
    .B(_04572_),
    .C(_04573_),
    .Y(_04580_));
 sky130_fd_sc_hd__nand2_1 _10401_ (.A(_02364_),
    .B(_02358_),
    .Y(_04581_));
 sky130_fd_sc_hd__nand2_1 _10402_ (.A(_04581_),
    .B(_01780_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_1 _10403_ (.A(_04582_),
    .B(_01786_),
    .Y(_04583_));
 sky130_fd_sc_hd__inv_2 _10404_ (.A(_01148_),
    .Y(_04584_));
 sky130_fd_sc_hd__nand2_1 _10405_ (.A(_04583_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__nand2_1 _10406_ (.A(_04585_),
    .B(_00513_),
    .Y(_04586_));
 sky130_fd_sc_hd__nand2_1 _10407_ (.A(_04586_),
    .B(_00511_),
    .Y(_04587_));
 sky130_fd_sc_hd__nand2_1 _10408_ (.A(_04587_),
    .B(_00770_),
    .Y(_04588_));
 sky130_fd_sc_hd__inv_2 _10409_ (.A(_00770_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand3_1 _10410_ (.A(_04586_),
    .B(_04589_),
    .C(_00511_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand2_1 _10411_ (.A(_04588_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__inv_2 _10412_ (.A(net161),
    .Y(_04593_));
 sky130_fd_sc_hd__nand2_1 _10413_ (.A(_04592_),
    .B(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand3_1 _10414_ (.A(_04583_),
    .B(_00512_),
    .C(_04584_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand2_1 _10415_ (.A(_04586_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__inv_2 _10416_ (.A(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _10417_ (.A(_04597_),
    .B(net135),
    .Y(_04598_));
 sky130_fd_sc_hd__inv_2 _10418_ (.A(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__nand3_1 _10419_ (.A(_04588_),
    .B(net161),
    .C(_04591_),
    .Y(_04600_));
 sky130_fd_sc_hd__inv_2 _10420_ (.A(_04600_),
    .Y(_04602_));
 sky130_fd_sc_hd__a21oi_1 _10421_ (.A1(_04594_),
    .A2(_04599_),
    .B1(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__nor2_1 _10422_ (.A(_04580_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__nor2_1 _10423_ (.A(_04575_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__inv_2 _10424_ (.A(_01783_),
    .Y(_04606_));
 sky130_fd_sc_hd__nand2_1 _10425_ (.A(_04582_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__nand3_1 _10426_ (.A(_04581_),
    .B(_01783_),
    .C(_01780_),
    .Y(_04608_));
 sky130_fd_sc_hd__nand3_1 _10427_ (.A(_04607_),
    .B(net124),
    .C(_04608_),
    .Y(_04609_));
 sky130_fd_sc_hd__nand2_1 _10428_ (.A(_04607_),
    .B(_01138_),
    .Y(_04610_));
 sky130_fd_sc_hd__inv_2 _10429_ (.A(_01784_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_1 _10430_ (.A(_04610_),
    .B(_04611_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand3_1 _10431_ (.A(_04607_),
    .B(_01784_),
    .C(_01138_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2_1 _10432_ (.A(_04613_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__inv_2 _10433_ (.A(net68),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _10434_ (.A(_04615_),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__nand3_1 _10435_ (.A(_04613_),
    .B(_04614_),
    .C(net162),
    .Y(_04618_));
 sky130_fd_sc_hd__nand2_1 _10436_ (.A(_04617_),
    .B(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__o21ai_1 _10437_ (.A1(_04609_),
    .A2(_04619_),
    .B1(_04618_),
    .Y(_04620_));
 sky130_fd_sc_hd__nand2_1 _10438_ (.A(_04607_),
    .B(_04608_),
    .Y(_04621_));
 sky130_fd_sc_hd__inv_2 _10439_ (.A(net124),
    .Y(_04622_));
 sky130_fd_sc_hd__nand2_1 _10440_ (.A(_04621_),
    .B(_04622_),
    .Y(_04624_));
 sky130_fd_sc_hd__nand2_1 _10441_ (.A(_04624_),
    .B(_04609_),
    .Y(_04625_));
 sky130_fd_sc_hd__inv_2 _10442_ (.A(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__nand3_1 _10443_ (.A(_04617_),
    .B(_04618_),
    .C(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__nor2_1 _10444_ (.A(_02361_),
    .B(_02363_),
    .Y(_04628_));
 sky130_fd_sc_hd__nand2_1 _10445_ (.A(_02358_),
    .B(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__nand2_1 _10446_ (.A(_04629_),
    .B(_01778_),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _10447_ (.A(_01485_),
    .B(_01500_),
    .Y(_04631_));
 sky130_fd_sc_hd__inv_2 _10448_ (.A(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand2_1 _10449_ (.A(_04630_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_04633_),
    .B(_01485_),
    .Y(_04635_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_04635_),
    .B(_01497_),
    .Y(_04636_));
 sky130_fd_sc_hd__inv_2 _10452_ (.A(_01497_),
    .Y(_04637_));
 sky130_fd_sc_hd__nand3_1 _10453_ (.A(_04633_),
    .B(_01485_),
    .C(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand2_1 _10454_ (.A(_04636_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__inv_2 _10455_ (.A(net158),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2_1 _10456_ (.A(_04639_),
    .B(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand2b_1 _10457_ (.A_N(_04630_),
    .B(_04631_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand3_1 _10458_ (.A(_04642_),
    .B(net142),
    .C(_04633_),
    .Y(_04643_));
 sky130_fd_sc_hd__inv_2 _10459_ (.A(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__nand3_1 _10460_ (.A(_04636_),
    .B(net158),
    .C(_04638_),
    .Y(_04646_));
 sky130_fd_sc_hd__inv_2 _10461_ (.A(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__a21oi_1 _10462_ (.A1(_04641_),
    .A2(_04644_),
    .B1(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__nor2_1 _10463_ (.A(_04627_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__nor2_1 _10464_ (.A(_04620_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__inv_2 _10465_ (.A(_02361_),
    .Y(_04651_));
 sky130_fd_sc_hd__nand2_1 _10466_ (.A(_02358_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__nand3_1 _10467_ (.A(_02208_),
    .B(_02356_),
    .C(_02361_),
    .Y(_04653_));
 sky130_fd_sc_hd__nand3_1 _10468_ (.A(_04652_),
    .B(_04653_),
    .C(net132),
    .Y(_04654_));
 sky130_fd_sc_hd__nand2_1 _10469_ (.A(_04652_),
    .B(_02359_),
    .Y(_04655_));
 sky130_fd_sc_hd__inv_2 _10470_ (.A(_02363_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _10471_ (.A(_04655_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__nand3_1 _10472_ (.A(_04652_),
    .B(_02363_),
    .C(_02359_),
    .Y(_04659_));
 sky130_fd_sc_hd__nand2_1 _10473_ (.A(_04658_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__inv_2 _10474_ (.A(net95),
    .Y(_04661_));
 sky130_fd_sc_hd__nand2_1 _10475_ (.A(_04660_),
    .B(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__nand3_1 _10476_ (.A(_04658_),
    .B(net156),
    .C(_04659_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand2_1 _10477_ (.A(_04662_),
    .B(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__o21ai_1 _10478_ (.A1(_04654_),
    .A2(_04664_),
    .B1(_04663_),
    .Y(_04665_));
 sky130_fd_sc_hd__nand2_1 _10479_ (.A(_04652_),
    .B(_04653_),
    .Y(_04666_));
 sky130_fd_sc_hd__inv_2 _10480_ (.A(net132),
    .Y(_04668_));
 sky130_fd_sc_hd__nand2_1 _10481_ (.A(_04666_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand2_1 _10482_ (.A(_04669_),
    .B(_04654_),
    .Y(_04670_));
 sky130_fd_sc_hd__inv_2 _10483_ (.A(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__nand3_1 _10484_ (.A(_04662_),
    .B(_04663_),
    .C(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__inv_2 _10485_ (.A(_02354_),
    .Y(_04673_));
 sky130_fd_sc_hd__nand2_1 _10486_ (.A(_02347_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_1 _10487_ (.A(_04674_),
    .B(_02200_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand2_1 _10488_ (.A(_04675_),
    .B(_02205_),
    .Y(_04676_));
 sky130_fd_sc_hd__nand2_1 _10489_ (.A(_04676_),
    .B(_02029_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2_1 _10490_ (.A(_02037_),
    .B(_02033_),
    .Y(_04679_));
 sky130_fd_sc_hd__inv_2 _10491_ (.A(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__nand2_1 _10492_ (.A(_04677_),
    .B(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand3_1 _10493_ (.A(_04676_),
    .B(_02029_),
    .C(_04679_),
    .Y(_04682_));
 sky130_fd_sc_hd__nand2_1 _10494_ (.A(_04681_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__inv_2 _10495_ (.A(net159),
    .Y(_04684_));
 sky130_fd_sc_hd__nand2_1 _10496_ (.A(_04683_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__or2_1 _10497_ (.A(_02205_),
    .B(_04675_),
    .X(_04686_));
 sky130_fd_sc_hd__nand3_1 _10498_ (.A(_04686_),
    .B(net145),
    .C(_04676_),
    .Y(_04687_));
 sky130_fd_sc_hd__inv_2 _10499_ (.A(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__nand3_1 _10500_ (.A(_04681_),
    .B(net159),
    .C(_04682_),
    .Y(_04690_));
 sky130_fd_sc_hd__a21boi_1 _10501_ (.A1(_04685_),
    .A2(_04688_),
    .B1_N(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__nor2_1 _10502_ (.A(_04672_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__nor2_1 _10503_ (.A(_04665_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__nand2_1 _10504_ (.A(_04686_),
    .B(_04676_),
    .Y(_04694_));
 sky130_fd_sc_hd__inv_2 _10505_ (.A(net145),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_1 _10506_ (.A(_04694_),
    .B(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__nand2_1 _10507_ (.A(_04696_),
    .B(_04687_),
    .Y(_04697_));
 sky130_fd_sc_hd__inv_2 _10508_ (.A(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__nand3_1 _10509_ (.A(_04698_),
    .B(_04685_),
    .C(_04690_),
    .Y(_04699_));
 sky130_fd_sc_hd__nor2_1 _10510_ (.A(_04672_),
    .B(_04699_),
    .Y(_04701_));
 sky130_fd_sc_hd__or2_1 _10511_ (.A(_02343_),
    .B(_02337_),
    .X(_04702_));
 sky130_fd_sc_hd__nand2_1 _10512_ (.A(_04702_),
    .B(_02344_),
    .Y(_04703_));
 sky130_fd_sc_hd__inv_2 _10513_ (.A(net122),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2_1 _10514_ (.A(_04703_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__inv_2 _10515_ (.A(net149),
    .Y(_04706_));
 sky130_fd_sc_hd__a21o_1 _10516_ (.A1(_02301_),
    .A2(_02303_),
    .B1(_02334_),
    .X(_04707_));
 sky130_fd_sc_hd__nand2_2 _10517_ (.A(_04707_),
    .B(_02336_),
    .Y(_04708_));
 sky130_fd_sc_hd__or2_1 _10518_ (.A(_04706_),
    .B(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__inv_2 _10519_ (.A(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand3_1 _10520_ (.A(_04702_),
    .B(net122),
    .C(_02344_),
    .Y(_04712_));
 sky130_fd_sc_hd__a21boi_1 _10521_ (.A1(_04705_),
    .A2(_04710_),
    .B1_N(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__nand2_1 _10522_ (.A(_02352_),
    .B(_02353_),
    .Y(_04714_));
 sky130_fd_sc_hd__inv_2 _10523_ (.A(_04714_),
    .Y(_04715_));
 sky130_fd_sc_hd__or2_1 _10524_ (.A(_04715_),
    .B(_02347_),
    .X(_04716_));
 sky130_fd_sc_hd__nand2_1 _10525_ (.A(_02347_),
    .B(_04715_),
    .Y(_04717_));
 sky130_fd_sc_hd__nand2_1 _10526_ (.A(_04716_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__inv_2 _10527_ (.A(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__nor2_1 _10528_ (.A(net150),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__nand2_1 _10529_ (.A(_04719_),
    .B(net150),
    .Y(_04721_));
 sky130_fd_sc_hd__o21ai_1 _10530_ (.A1(_04713_),
    .A2(_04720_),
    .B1(_04721_),
    .Y(_04723_));
 sky130_fd_sc_hd__inv_2 _10531_ (.A(net157),
    .Y(_04724_));
 sky130_fd_sc_hd__nand2_1 _10532_ (.A(_04717_),
    .B(_02352_),
    .Y(_04725_));
 sky130_fd_sc_hd__or2_1 _10533_ (.A(_02351_),
    .B(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__nand2_1 _10534_ (.A(_04725_),
    .B(_02351_),
    .Y(_04727_));
 sky130_fd_sc_hd__nand2_1 _10535_ (.A(_04726_),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__or2_1 _10536_ (.A(_04724_),
    .B(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__nand2_1 _10537_ (.A(_04728_),
    .B(_04724_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand3_1 _10538_ (.A(_04723_),
    .B(_04729_),
    .C(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__nand2_1 _10539_ (.A(_04731_),
    .B(_04729_),
    .Y(_04732_));
 sky130_fd_sc_hd__nand2_1 _10540_ (.A(_04701_),
    .B(_04732_),
    .Y(_04734_));
 sky130_fd_sc_hd__nand2_1 _10541_ (.A(_04693_),
    .B(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_04642_),
    .B(_04633_),
    .Y(_04736_));
 sky130_fd_sc_hd__inv_2 _10543_ (.A(net142),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_1 _10544_ (.A(_04736_),
    .B(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__nand2_1 _10545_ (.A(_04738_),
    .B(_04643_),
    .Y(_04739_));
 sky130_fd_sc_hd__inv_2 _10546_ (.A(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand3_1 _10547_ (.A(_04740_),
    .B(_04641_),
    .C(_04646_),
    .Y(_04741_));
 sky130_fd_sc_hd__nor2_1 _10548_ (.A(_04627_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_1 _10549_ (.A(_04735_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _10550_ (.A(_04650_),
    .B(_04743_),
    .Y(_04745_));
 sky130_fd_sc_hd__a21o_1 _10551_ (.A1(_04586_),
    .A2(_04595_),
    .B1(net135),
    .X(_04746_));
 sky130_fd_sc_hd__nand2_1 _10552_ (.A(_04746_),
    .B(_04598_),
    .Y(_04747_));
 sky130_fd_sc_hd__inv_2 _10553_ (.A(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__nand3_1 _10554_ (.A(_04748_),
    .B(_04594_),
    .C(_04600_),
    .Y(_04749_));
 sky130_fd_sc_hd__nor2_1 _10555_ (.A(_04580_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__nand2_1 _10556_ (.A(_04745_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand2_2 _10557_ (.A(_04605_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _10558_ (.A(_04544_),
    .B(_04545_),
    .Y(_04753_));
 sky130_fd_sc_hd__inv_2 _10559_ (.A(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__nand2_1 _10560_ (.A(_04547_),
    .B(_04538_),
    .Y(_04756_));
 sky130_fd_sc_hd__inv_2 _10561_ (.A(net153),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _10562_ (.A(_04756_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _10563_ (.A(_04758_),
    .B(_04548_),
    .Y(_04759_));
 sky130_fd_sc_hd__inv_2 _10564_ (.A(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_1 _10565_ (.A(_04754_),
    .B(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__nor2_1 _10566_ (.A(_04559_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__nand2_1 _10567_ (.A(_04752_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__nand2b_1 _10568_ (.A_N(_04562_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand3_1 _10569_ (.A(_03953_),
    .B(_03956_),
    .C(_04243_),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _10570_ (.A(_04245_),
    .B(_04765_),
    .Y(_04767_));
 sky130_fd_sc_hd__inv_2 _10571_ (.A(net163),
    .Y(_04768_));
 sky130_fd_sc_hd__nand2_1 _10572_ (.A(_04767_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__nand3_2 _10573_ (.A(_04245_),
    .B(_04765_),
    .C(net163),
    .Y(_04770_));
 sky130_fd_sc_hd__nand2_1 _10574_ (.A(_04769_),
    .B(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__inv_4 _10575_ (.A(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand2_1 _10576_ (.A(_04764_),
    .B(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__nand2_1 _10577_ (.A(_04773_),
    .B(_04770_),
    .Y(_04774_));
 sky130_fd_sc_hd__xor2_1 _10578_ (.A(_04519_),
    .B(_04774_),
    .X(\absum[21] ));
 sky130_fd_sc_hd__nand3_1 _10579_ (.A(_04764_),
    .B(_04772_),
    .C(_04519_),
    .Y(_04775_));
 sky130_fd_sc_hd__inv_2 _10580_ (.A(_04770_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand3_1 _10581_ (.A(_04516_),
    .B(_04777_),
    .C(_04517_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_04778_),
    .B(_04517_),
    .Y(_04779_));
 sky130_fd_sc_hd__inv_2 _10583_ (.A(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _10584_ (.A(_04775_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__xor2_1 _10585_ (.A(net114),
    .B(_04781_),
    .X(\absum[22] ));
 sky130_fd_sc_hd__nand2_1 _10586_ (.A(_04781_),
    .B(net80),
    .Y(_04782_));
 sky130_fd_sc_hd__nand2_1 _10587_ (.A(_04782_),
    .B(net106),
    .Y(_04783_));
 sky130_fd_sc_hd__nand3b_1 _10588_ (.A_N(net106),
    .B(_04781_),
    .C(net80),
    .Y(_04784_));
 sky130_fd_sc_hd__nand2_1 _10589_ (.A(net107),
    .B(_04784_),
    .Y(\absum[23] ));
 sky130_fd_sc_hd__nand2_1 _10590_ (.A(net114),
    .B(net106),
    .Y(_04786_));
 sky130_fd_sc_hd__nand3_1 _10591_ (.A(_04516_),
    .B(_04772_),
    .C(_04517_),
    .Y(_04787_));
 sky130_fd_sc_hd__nor2_1 _10592_ (.A(_04786_),
    .B(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand3_1 _10593_ (.A(_04788_),
    .B(_04752_),
    .C(_04762_),
    .Y(_04789_));
 sky130_fd_sc_hd__inv_2 _10594_ (.A(_04786_),
    .Y(_04790_));
 sky130_fd_sc_hd__nand2_1 _10595_ (.A(_04779_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__nand2_1 _10596_ (.A(_04788_),
    .B(_04562_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand3_2 _10597_ (.A(_04789_),
    .B(_04791_),
    .C(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__or2_1 _10598_ (.A(net148),
    .B(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__nand2_1 _10599_ (.A(_04793_),
    .B(net148),
    .Y(_04795_));
 sky130_fd_sc_hd__and2_1 _10600_ (.A(_04794_),
    .B(_04795_),
    .X(_04797_));
 sky130_fd_sc_hd__clkbuf_1 _10601_ (.A(_04797_),
    .X(\absum[24] ));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(net164),
    .B(net116),
    .Y(_04798_));
 sky130_fd_sc_hd__nand3_1 _10603_ (.A(_04519_),
    .B(_04772_),
    .C(_04790_),
    .Y(_04799_));
 sky130_fd_sc_hd__nor2_1 _10604_ (.A(_04799_),
    .B(_04763_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand2_1 _10605_ (.A(_04792_),
    .B(_04791_),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _10606_ (.A(_04800_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__nor2_1 _10607_ (.A(_04798_),
    .B(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__a21oi_1 _10608_ (.A1(_04793_),
    .A2(net82),
    .B1(net116),
    .Y(_04804_));
 sky130_fd_sc_hd__nor2_1 _10609_ (.A(_04803_),
    .B(net117),
    .Y(\absum[25] ));
 sky130_fd_sc_hd__nor2_1 _10610_ (.A(net119),
    .B(_04803_),
    .Y(_04806_));
 sky130_fd_sc_hd__nand2_1 _10611_ (.A(_04803_),
    .B(net119),
    .Y(_04807_));
 sky130_fd_sc_hd__inv_2 _10612_ (.A(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__nor2_1 _10613_ (.A(net120),
    .B(_04808_),
    .Y(\absum[26] ));
 sky130_fd_sc_hd__inv_2 _10614_ (.A(net111),
    .Y(_04809_));
 sky130_fd_sc_hd__nand2_1 _10615_ (.A(_04808_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__nand2_1 _10616_ (.A(_04807_),
    .B(net111),
    .Y(_04811_));
 sky130_fd_sc_hd__nand2_1 _10617_ (.A(_04810_),
    .B(net112),
    .Y(\absum[27] ));
 sky130_fd_sc_hd__or3b_1 _10618_ (.A(_04809_),
    .B(_04798_),
    .C_N(net119),
    .X(_04812_));
 sky130_fd_sc_hd__nor2_1 _10619_ (.A(_04812_),
    .B(_04802_),
    .Y(_04813_));
 sky130_fd_sc_hd__nor2_1 _10620_ (.A(net138),
    .B(_04813_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _10621_ (.A(_04813_),
    .B(net138),
    .Y(_04816_));
 sky130_fd_sc_hd__nor2b_1 _10622_ (.A(net139),
    .B_N(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_04817_),
    .X(\absum[28] ));
 sky130_fd_sc_hd__nand2_1 _10624_ (.A(_04816_),
    .B(net100),
    .Y(_04818_));
 sky130_fd_sc_hd__nand3b_1 _10625_ (.A_N(net100),
    .B(_04813_),
    .C(net86),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _10626_ (.A(net101),
    .B(_04819_),
    .Y(\absum[29] ));
 sky130_fd_sc_hd__inv_2 _10627_ (.A(_04812_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _10628_ (.A(net86),
    .B(net100),
    .Y(_04821_));
 sky130_fd_sc_hd__inv_2 _10629_ (.A(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand3_1 _10630_ (.A(_04793_),
    .B(_04820_),
    .C(_04822_),
    .Y(_04824_));
 sky130_fd_sc_hd__xnor2_1 _10631_ (.A(net109),
    .B(_04824_),
    .Y(\absum[30] ));
 sky130_fd_sc_hd__nand3_1 _10632_ (.A(_04813_),
    .B(net89),
    .C(_04822_),
    .Y(_04825_));
 sky130_fd_sc_hd__nand2_1 _10633_ (.A(_04825_),
    .B(net103),
    .Y(_04826_));
 sky130_fd_sc_hd__inv_2 _10634_ (.A(_04824_),
    .Y(_04827_));
 sky130_fd_sc_hd__inv_2 _10635_ (.A(net103),
    .Y(_04828_));
 sky130_fd_sc_hd__nand3_1 _10636_ (.A(_04827_),
    .B(net89),
    .C(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(net104),
    .B(_04829_),
    .Y(\absum[31] ));
 sky130_fd_sc_hd__nand2_1 _10638_ (.A(_04708_),
    .B(_04706_),
    .Y(_04830_));
 sky130_fd_sc_hd__and2_1 _10639_ (.A(_04709_),
    .B(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__clkbuf_1 _10640_ (.A(_04831_),
    .X(\absum[0] ));
 sky130_fd_sc_hd__nand2_1 _10641_ (.A(_04705_),
    .B(_04712_),
    .Y(_04833_));
 sky130_fd_sc_hd__xor2_1 _10642_ (.A(_04709_),
    .B(_04833_),
    .X(\absum[1] ));
 sky130_fd_sc_hd__or2b_1 _10643_ (.A(_04720_),
    .B_N(_04721_),
    .X(_04834_));
 sky130_fd_sc_hd__xor2_1 _10644_ (.A(_04713_),
    .B(_04834_),
    .X(\absum[2] ));
 sky130_fd_sc_hd__a21o_1 _10645_ (.A1(_04729_),
    .A2(_04730_),
    .B1(_04723_),
    .X(_04835_));
 sky130_fd_sc_hd__and2_1 _10646_ (.A(_04835_),
    .B(_04731_),
    .X(_04836_));
 sky130_fd_sc_hd__clkbuf_1 _10647_ (.A(_04836_),
    .X(\absum[3] ));
 sky130_fd_sc_hd__or2_1 _10648_ (.A(_04698_),
    .B(_04732_),
    .X(_04837_));
 sky130_fd_sc_hd__nand2_1 _10649_ (.A(_04732_),
    .B(_04698_),
    .Y(_04838_));
 sky130_fd_sc_hd__and2_1 _10650_ (.A(_04837_),
    .B(_04838_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _10651_ (.A(_04840_),
    .X(\absum[4] ));
 sky130_fd_sc_hd__nand2_1 _10652_ (.A(_04685_),
    .B(_04690_),
    .Y(_04841_));
 sky130_fd_sc_hd__nand2_1 _10653_ (.A(_04838_),
    .B(_04687_),
    .Y(_04842_));
 sky130_fd_sc_hd__xnor2_1 _10654_ (.A(_04841_),
    .B(net146),
    .Y(\absum[5] ));
 sky130_fd_sc_hd__o21ai_1 _10655_ (.A1(_04841_),
    .A2(_04838_),
    .B1(_04691_),
    .Y(_04843_));
 sky130_fd_sc_hd__or2_1 _10656_ (.A(_04671_),
    .B(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__nand2_1 _10657_ (.A(_04843_),
    .B(_04671_),
    .Y(_04845_));
 sky130_fd_sc_hd__and2_1 _10658_ (.A(_04844_),
    .B(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__clkbuf_1 _10659_ (.A(_04846_),
    .X(\absum[6] ));
 sky130_fd_sc_hd__nand2_1 _10660_ (.A(_04845_),
    .B(_04654_),
    .Y(_04848_));
 sky130_fd_sc_hd__xnor2_1 _10661_ (.A(_04664_),
    .B(net133),
    .Y(\absum[7] ));
 sky130_fd_sc_hd__inv_2 _10662_ (.A(_04735_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_1 _10663_ (.A(_04849_),
    .B(_04739_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _10664_ (.A(_04735_),
    .B(_04740_),
    .Y(_04851_));
 sky130_fd_sc_hd__and2_1 _10665_ (.A(_04850_),
    .B(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _10666_ (.A(_04852_),
    .X(\absum[8] ));
 sky130_fd_sc_hd__nand2_1 _10667_ (.A(_04641_),
    .B(_04646_),
    .Y(_04853_));
 sky130_fd_sc_hd__nand2_1 _10668_ (.A(_04851_),
    .B(_04643_),
    .Y(_04854_));
 sky130_fd_sc_hd__xnor2_1 _10669_ (.A(_04853_),
    .B(net143),
    .Y(\absum[9] ));
 sky130_fd_sc_hd__o21ai_1 _10670_ (.A1(_04741_),
    .A2(_04849_),
    .B1(_04648_),
    .Y(_04856_));
 sky130_fd_sc_hd__or2_1 _10671_ (.A(_04626_),
    .B(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__nand2_1 _10672_ (.A(_04856_),
    .B(_04626_),
    .Y(_04858_));
 sky130_fd_sc_hd__and2_1 _10673_ (.A(_04857_),
    .B(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__clkbuf_1 _10674_ (.A(_04859_),
    .X(\absum[10] ));
 sky130_fd_sc_hd__nand2_1 _10675_ (.A(_04858_),
    .B(_04609_),
    .Y(_04860_));
 sky130_fd_sc_hd__xnor2_1 _10676_ (.A(_04619_),
    .B(net125),
    .Y(\absum[11] ));
 sky130_fd_sc_hd__or2_1 _10677_ (.A(_04748_),
    .B(_04745_),
    .X(_04861_));
 sky130_fd_sc_hd__nand2_1 _10678_ (.A(_04745_),
    .B(_04748_),
    .Y(_04862_));
 sky130_fd_sc_hd__and2_1 _10679_ (.A(_04861_),
    .B(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__clkbuf_1 _10680_ (.A(_04863_),
    .X(\absum[12] ));
 sky130_fd_sc_hd__nand2_1 _10681_ (.A(_04594_),
    .B(_04600_),
    .Y(_04865_));
 sky130_fd_sc_hd__nand2_1 _10682_ (.A(_04862_),
    .B(_04598_),
    .Y(_04866_));
 sky130_fd_sc_hd__xnor2_1 _10683_ (.A(_04865_),
    .B(net136),
    .Y(\absum[13] ));
 sky130_fd_sc_hd__or2b_1 _10684_ (.A(_04749_),
    .B_N(_04745_),
    .X(_04867_));
 sky130_fd_sc_hd__nand2_1 _10685_ (.A(_04867_),
    .B(_04603_),
    .Y(_04868_));
 sky130_fd_sc_hd__or2_1 _10686_ (.A(_04578_),
    .B(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__nand2_1 _10687_ (.A(_04868_),
    .B(_04578_),
    .Y(_04870_));
 sky130_fd_sc_hd__and2_1 _10688_ (.A(_04869_),
    .B(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_04871_),
    .X(\absum[14] ));
 sky130_fd_sc_hd__nand2_1 _10690_ (.A(_04870_),
    .B(_04565_),
    .Y(_04873_));
 sky130_fd_sc_hd__xnor2_1 _10691_ (.A(_04574_),
    .B(net128),
    .Y(\absum[15] ));
 sky130_fd_sc_hd__inv_2 _10692_ (.A(_04752_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_1 _10693_ (.A(_04874_),
    .B(_04759_),
    .Y(_04875_));
 sky130_fd_sc_hd__nand2_1 _10694_ (.A(_04752_),
    .B(_04760_),
    .Y(_04876_));
 sky130_fd_sc_hd__and2_1 _10695_ (.A(net154),
    .B(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__clkbuf_1 _10696_ (.A(net155),
    .X(\absum[16] ));
 sky130_fd_sc_hd__nand2_1 _10697_ (.A(_04876_),
    .B(_04548_),
    .Y(_04878_));
 sky130_fd_sc_hd__xor2_1 _10698_ (.A(_04754_),
    .B(_04878_),
    .X(\absum[17] ));
 sky130_fd_sc_hd__o21bai_1 _10699_ (.A1(_04761_),
    .A2(_04874_),
    .B1_N(_04551_),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_1 _10700_ (.A(_04558_),
    .B(_04879_),
    .X(_04881_));
 sky130_fd_sc_hd__nand2_1 _10701_ (.A(_04879_),
    .B(_04558_),
    .Y(_04882_));
 sky130_fd_sc_hd__and2_1 _10702_ (.A(_04881_),
    .B(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__clkbuf_1 _10703_ (.A(_04883_),
    .X(\absum[18] ));
 sky130_fd_sc_hd__nand2_1 _10704_ (.A(_04552_),
    .B(_04532_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand2_1 _10705_ (.A(_04882_),
    .B(_04523_),
    .Y(_04885_));
 sky130_fd_sc_hd__xnor2_1 _10706_ (.A(_04884_),
    .B(_04885_),
    .Y(\absum[19] ));
 sky130_fd_sc_hd__or2_1 _10707_ (.A(_04772_),
    .B(_04764_),
    .X(_04886_));
 sky130_fd_sc_hd__and2_1 _10708_ (.A(_04886_),
    .B(_04773_),
    .X(_04887_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(_04887_),
    .X(\absum[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10710_ (.CLK(clknet_2_1__leaf_clk),
    .D(\absum[0] ),
    .RESET_B(net99),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _10711_ (.CLK(clknet_2_1__leaf_clk),
    .D(net123),
    .RESET_B(net99),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _10712_ (.CLK(clknet_2_1__leaf_clk),
    .D(\absum[2] ),
    .RESET_B(net99),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _10713_ (.CLK(clknet_2_1__leaf_clk),
    .D(\absum[3] ),
    .RESET_B(net99),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _10714_ (.CLK(clknet_2_1__leaf_clk),
    .D(\absum[4] ),
    .RESET_B(net99),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _10715_ (.CLK(clknet_2_1__leaf_clk),
    .D(net147),
    .RESET_B(net99),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _10716_ (.CLK(clknet_2_1__leaf_clk),
    .D(\absum[6] ),
    .RESET_B(net99),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_2 _10717_ (.CLK(clknet_2_1__leaf_clk),
    .D(net134),
    .RESET_B(net99),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _10718_ (.CLK(clknet_2_1__leaf_clk),
    .D(\absum[8] ),
    .RESET_B(net99),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _10719_ (.CLK(clknet_2_0__leaf_clk),
    .D(net144),
    .RESET_B(net99),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _10720_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[10] ),
    .RESET_B(net99),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_2 _10721_ (.CLK(clknet_2_0__leaf_clk),
    .D(net126),
    .RESET_B(net99),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _10722_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[12] ),
    .RESET_B(net99),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _10723_ (.CLK(clknet_2_0__leaf_clk),
    .D(net137),
    .RESET_B(net99),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _10724_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[14] ),
    .RESET_B(net99),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_2 _10725_ (.CLK(clknet_2_2__leaf_clk),
    .D(net129),
    .RESET_B(net98),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _10726_ (.CLK(clknet_2_2__leaf_clk),
    .D(\absum[16] ),
    .RESET_B(net98),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _10727_ (.CLK(clknet_2_2__leaf_clk),
    .D(net131),
    .RESET_B(net98),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _10728_ (.CLK(clknet_2_2__leaf_clk),
    .D(\absum[18] ),
    .RESET_B(net98),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _10729_ (.CLK(clknet_2_2__leaf_clk),
    .D(net141),
    .RESET_B(net98),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_2 _10730_ (.CLK(clknet_2_3__leaf_clk),
    .D(\absum[20] ),
    .RESET_B(net98),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_2 _10731_ (.CLK(clknet_2_3__leaf_clk),
    .D(net152),
    .RESET_B(net98),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_2 _10732_ (.CLK(clknet_2_2__leaf_clk),
    .D(net115),
    .RESET_B(net98),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _10733_ (.CLK(clknet_2_2__leaf_clk),
    .D(net108),
    .RESET_B(net98),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_2 _10734_ (.CLK(clknet_2_3__leaf_clk),
    .D(\absum[24] ),
    .RESET_B(net98),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _10735_ (.CLK(clknet_2_3__leaf_clk),
    .D(net118),
    .RESET_B(net98),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _10736_ (.CLK(clknet_2_3__leaf_clk),
    .D(net121),
    .RESET_B(net98),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _10737_ (.CLK(clknet_2_3__leaf_clk),
    .D(net113),
    .RESET_B(net98),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_2 _10738_ (.CLK(clknet_2_3__leaf_clk),
    .D(\absum[28] ),
    .RESET_B(net98),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _10739_ (.CLK(clknet_2_3__leaf_clk),
    .D(net102),
    .RESET_B(net98),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_2 _10740_ (.CLK(clknet_2_3__leaf_clk),
    .D(net110),
    .RESET_B(net98),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _10741_ (.CLK(clknet_2_3__leaf_clk),
    .D(net105),
    .RESET_B(net65),
    .Q(net90));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_8 fanout99 (.A(net65),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net87),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net89),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\absum[30] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net85),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_04811_),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\absum[27] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net80),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\absum[22] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net83),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_04804_),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\absum[25] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_04818_),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net84),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_04806_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\absum[26] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net77),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\absum[1] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net67),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_04860_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\absum[11] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net71),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_04873_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\absum[29] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\absum[15] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net74),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\absum[17] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net94),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_04848_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\absum[7] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net69),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_04866_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\absum[13] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net86),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net90),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_04815_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net76),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\absum[19] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net96),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_04854_),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\absum[9] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net92),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_04842_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\absum[5] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net82),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_04826_),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net66),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net88),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net79),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\absum[21] ),
    .X(net152));
 sky130_fd_sc_hd__buf_1 hold54 (.A(net73),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_04875_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_04877_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net95),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net91),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net97),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\absum[31] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net93),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net75),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net70),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net68),
    .X(net162));
 sky130_fd_sc_hd__buf_1 hold64 (.A(net78),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net82),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net81),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_04783_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\absum[23] ),
    .X(net108));
 sky130_fd_sc_hd__buf_4 input1 (.A(a_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(a_i[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a_i[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(a_i[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(a_i[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a_i[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a_i[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(a_i[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(a_i[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(a_i[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(a_i[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a_i[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(a_i[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(a_i[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(a_i[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(a_i[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(a_i[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(a_i[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(a_i[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(a_i[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a_i[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a_i[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a_i[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(a_i[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(a_i[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a_i[9]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(b_i[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(b_i[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(b_i[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(b_i[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(b_i[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(b_i[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(b_i[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(a_i[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input40 (.A(b_i[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(b_i[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(b_i[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(b_i[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(b_i[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(b_i[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(b_i[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(b_i[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(b_i[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(b_i[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(a_i[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input50 (.A(b_i[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(b_i[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(b_i[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(b_i[28]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(b_i[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input55 (.A(b_i[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(b_i[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(b_i[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(b_i[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(b_i[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input6 (.A(a_i[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b_i[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b_i[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b_i[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(b_i[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(b_i[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(nrst),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input7 (.A(a_i[15]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(a_i[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(a_i[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(y_o[0]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(y_o[10]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(y_o[11]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(y_o[12]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(y_o[13]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(y_o[14]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(y_o[15]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(y_o[16]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(y_o[17]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(y_o[18]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(y_o[19]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(y_o[1]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(y_o[20]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(y_o[21]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(y_o[22]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(y_o[23]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(y_o[24]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(y_o[25]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(y_o[26]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(y_o[27]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(y_o[28]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(y_o[29]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(y_o[2]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(y_o[30]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(y_o[31]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(y_o[3]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(y_o[4]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(y_o[5]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(y_o[6]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(y_o[7]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(y_o[8]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(y_o[9]));
endmodule

