// This is the unpowered netlist.
module busarb_2_2 (clk_i,
    nrst_i,
    mports_i,
    mports_o,
    sports_i,
    sports_o);
 input clk_i;
 input nrst_i;
 input [227:0] mports_i;
 output [135:0] mports_o;
 input [135:0] sports_i;
 output [227:0] sports_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire \arbiter.master_handled[0] ;
 wire \arbiter.master_handled[1] ;
 wire \arbiter.master_handled[2] ;
 wire \arbiter.master_handled[3] ;
 wire \arbiter.master_sel[0][0] ;
 wire \arbiter.master_sel[0][1] ;
 wire \arbiter.slave_handled[0] ;
 wire \arbiter.slave_handled[1] ;
 wire \arbiter.slave_handled[2] ;
 wire \arbiter.slave_handled[3] ;
 wire \arbiter.slave_sel[0][0] ;
 wire \arbiter.slave_sel[0][1] ;
 wire \arbiter.state[0][0] ;
 wire \arbiter.state[0][1] ;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_1_1__leaf_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(mports_i[88]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(mports_i[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(mports_i[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(mports_i[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__A (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__B (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1217__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1220__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__A1 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__B1 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1223__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__B1 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__B2 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__A1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__B2 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1229__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1229__B2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__A1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__B2 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__B2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__B (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1234__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__B1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1240__A2 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1240__B2 (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1241__B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__1242__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1242__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__B1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__A2 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__B2 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__A (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__B2 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__A (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__A (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__B2 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__A (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__A (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1276__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__A (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1280__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1280__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__A (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__A (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__A2 (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__B2 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__A (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__A (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1298__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__A (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1310__A (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1313__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1315__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1321__A (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__B (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1338__A (.DIODE(_1093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__A (.DIODE(_1099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__B (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1341__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1342__A (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__A (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1352__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__A (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__A1 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__A2 (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__A3 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__A (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__B (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1364__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__C (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1377__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__A (.DIODE(_1099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__A (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__A (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__A (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__B (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__A (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__A (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__A2 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A1 (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A2 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1399__B (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__A (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__B (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__C (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1418__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1421__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1426__A (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1426__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__B (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1432__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1433__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1436__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__B (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__A (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__A (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__A (.DIODE(_0018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__A (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1454__B (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A3 (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1456__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__B1 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1460__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__A (.DIODE(_0031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__A (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__A (.DIODE(_0031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__A (.DIODE(_0031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__A (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__A (.DIODE(_0047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__A (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1490__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__A (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__A (.DIODE(_0047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__A (.DIODE(_0047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1508__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__B (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A (.DIODE(_0077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1516__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A (.DIODE(_0091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__B (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A (.DIODE(_0091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A1 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A2 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A2 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A (.DIODE(_0091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__A (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__B (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__B (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__B (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__A (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__B (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__C1 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1564__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1564__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__A (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__B (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__C (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__B1 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__B (.DIODE(_0137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A (.DIODE(_0139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__B (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__B (.DIODE(_0139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__B (.DIODE(_0144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__A (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__A (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__C (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__B (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__C (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__A2 (.DIODE(_0146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__A1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__A2 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__B1 (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__A (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__B (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__A2 (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__C (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__A (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__C (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A2 (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__B (.DIODE(_0173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__C (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__C (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__A (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__A (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__C (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__B (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__C (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__A2 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__B (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__A (.DIODE(_0196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__B (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__A3 (.DIODE(_0196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__A (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__A (.DIODE(_0196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1657__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1657__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1658__B1 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1659__B (.DIODE(_0210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1662__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__B (.DIODE(_0210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__C (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__A (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__A (.DIODE(_0219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__A (.DIODE(_0196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__B (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__B (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__C (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__B (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__A (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__A (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__A (.DIODE(_0254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1711__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__A (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__C (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__A (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__B (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__A (.DIODE(_0285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1739__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__A (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__A (.DIODE(_0296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__A (.DIODE(_0298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__A (.DIODE(_0298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__C (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__A (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__A2 (.DIODE(_0299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__A (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__A (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__A (.DIODE(_0311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__B (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__A (.DIODE(_0298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__A (.DIODE(_0311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1771__A2 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__A (.DIODE(_0311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__A (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__A (.DIODE(_0298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__C (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__A (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__A (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__A (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__B (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__A3 (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1829__C1 (.DIODE(_0372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__C (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__B (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__A (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__A (.DIODE(_0254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (.DIODE(_0254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__A (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__A2 (.DIODE(_0391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__A (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__A (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A1 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A2 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__B2 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__A (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__C (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__B1 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__A (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__A (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__A (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__B (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__C (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__A (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__B (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__A (.DIODE(_0448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__A (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1917__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1917__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1926__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A (.DIODE(_0448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__B (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__C (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__A2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__A (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__A (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__A (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__A (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__A (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__A (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__A (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__B (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__A (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A2 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__B1 (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__A2 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__A (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__A (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__A (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__A2 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__B1 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__B2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__A (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__A (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__B (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1999__C (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2001__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A (.DIODE(_0448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__A (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__C (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__C (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__B (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__B (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__A (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__A (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__C (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__B (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__C1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__A (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__A (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__A (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__A2 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__B (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__A (.DIODE(_0583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__C (.DIODE(_1134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__B (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__A (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__A (.DIODE(_0583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__A (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2073__B (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__B (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A3 (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__C (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__B (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__A (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__A (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__B (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__C1 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__A (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__A (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__A (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__B1 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__A1 (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__A (.DIODE(_0638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__A (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A1 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A2 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__B2 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__A (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__A (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__B (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__B (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__A (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__B (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__B2 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__A (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__B (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__B2 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__A (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__B (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__A (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__A1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__B (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2159__A (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__A (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__A (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__B2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__A1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__A (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__B2 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__A1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__A1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__B2 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__B2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__A1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__B2 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__A2 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__B2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2179__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__C (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__B1 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__B2 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__B (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__B (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__A (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__A (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__A (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__A (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__A (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__A (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__A (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__B (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__B (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__B (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__B1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__A (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__B1 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__A (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A2 (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A3 (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A2 (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__B1 (.DIODE(_0031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__A1 (.DIODE(_0047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__B1 (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__B1 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__C (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__B (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A2 (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__A2 (.DIODE(_0139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A2 (.DIODE(_0146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A2 (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A2 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A2 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A1_N (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__B1 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__A1 (.DIODE(_0196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__B1 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__A1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__A2 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__A2 (.DIODE(_0299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__B1 (.DIODE(_0311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__A (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A2 (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A3 (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A1 (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__B1 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A1 (.DIODE(_0254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__A1 (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__A1 (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__B1 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__B (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A2 (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A3 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__A1_N (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__B1 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__A1 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A2 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A1_N (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__B1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__A2 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__B1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__B1 (.DIODE(_0448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__B (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A2 (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A3 (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__A1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__A (.DIODE(_0583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__B (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A2 (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A3 (.DIODE(_0583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2323__B (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__A1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__A2 (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__A3 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__B1 (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__B (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__B (.DIODE(_0745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__B (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__B (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__A (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__B (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__B (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__B (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2347__A (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__A (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__A (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__A (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__A (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__A (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A2 (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__A (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__A2 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__A3 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A2 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__B1 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__B (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A2 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A3 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__B (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__A (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__A (.DIODE(_0047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__A (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__B (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A2 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A3 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A2 (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__B1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A1 (.DIODE(_0139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__B (.DIODE(_0146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A1 (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__C (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__B (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__A (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__B (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A2 (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__B (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__B (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__B1 (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A (.DIODE(_0219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__C (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A1 (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__C (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__A2 (.DIODE(_0299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__B1 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__A (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__B (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A1 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A3 (.DIODE(_0311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__A (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__B (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__B (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A1 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__B2 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A1 (.DIODE(_0254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__B2 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__C (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__C (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__B1 (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__B (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A1 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A3 (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__B2 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__B (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__C (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__A (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__C (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A1 (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__B1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__A2 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__B1 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A1_N (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__B1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A (.DIODE(_0448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__A (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__A1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__A2 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__A (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__B (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A1 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A3 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__A (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A1 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__B1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__B (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A1 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A3 (.DIODE(_0583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__A2 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__B1 (.DIODE(_0504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__B (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__B2 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__B (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__A (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__B (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__B (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__B (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__B (.DIODE(_0034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__C (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__C (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__A (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__B (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__B (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__B (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__A (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__A (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__A (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__A (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__B (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__B (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__A (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__B (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__B (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__B (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__B (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A2 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__B (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__B (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__A (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__A (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__B (.DIODE(_0139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__B (.DIODE(_0146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__B (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__B (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A (.DIODE(_0219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__B (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__B (.DIODE(_0299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__A (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__B (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A (.DIODE(_0391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__B (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__B (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__A (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__B (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__B (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__B (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__A (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__B (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__A (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__B (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__A (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__B (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__A (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__B (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__B (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__B (.DIODE(_0745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__B (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__A (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__A (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__B (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__B (.DIODE(_1102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A1 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A1 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__B (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__B (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__B (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__B (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__B (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__B (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__C (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A (.DIODE(_1020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__B (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__C (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__C (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__C (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__B (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__C (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__B (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__B (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__C (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_output512_A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_output515_A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_output674_A (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_output686_A (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_output694_A (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_output720_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_output729_A (.DIODE(net729));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _1201_ (.A(net768),
    .Y(_0980_));
 sky130_fd_sc_hd__buf_6 _1202_ (.A(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__buf_8 _1203_ (.A(net765),
    .X(_0982_));
 sky130_fd_sc_hd__buf_8 _1204_ (.A(net769),
    .X(_0983_));
 sky130_fd_sc_hd__nor2_8 _1205_ (.A(_0982_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__clkinv_4 _1206_ (.A(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__nor2_4 _1207_ (.A(_0981_),
    .B(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__clkinv_4 _1208_ (.A(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__buf_8 _1209_ (.A(\arbiter.slave_sel[0][0] ),
    .X(_0988_));
 sky130_fd_sc_hd__inv_2 _1210_ (.A(net770),
    .Y(_0989_));
 sky130_fd_sc_hd__nor2_2 _1211_ (.A(_0988_),
    .B(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__buf_6 _1212_ (.A(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_2 _1213_ (.A(_0989_),
    .B(_0988_),
    .Y(_0992_));
 sky130_fd_sc_hd__inv_2 _1214_ (.A(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__buf_8 _1215_ (.A(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__nand2_8 _1216_ (.A(_0988_),
    .B(\arbiter.slave_sel[0][1] ),
    .Y(_0995_));
 sky130_fd_sc_hd__clkinv_8 _1217_ (.A(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__nand2_1 _1218_ (.A(_0996_),
    .B(net233),
    .Y(_0997_));
 sky130_fd_sc_hd__nor2_8 _1219_ (.A(_0988_),
    .B(\arbiter.slave_sel[0][1] ),
    .Y(_0998_));
 sky130_fd_sc_hd__nand2_1 _1220_ (.A(_0998_),
    .B(net230),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2_1 _1221_ (.A(_0997_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__a221oi_2 _1222_ (.A1(_0991_),
    .A2(net330),
    .B1(_0994_),
    .B2(net293),
    .C1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__nor2_1 _1223_ (.A(_0987_),
    .B(net730),
    .Y(net366));
 sky130_fd_sc_hd__buf_6 _1224_ (.A(_0990_),
    .X(_1002_));
 sky130_fd_sc_hd__a22o_1 _1225_ (.A1(_0998_),
    .A2(net277),
    .B1(_1002_),
    .B2(net331),
    .X(_1003_));
 sky130_fd_sc_hd__a221oi_2 _1226_ (.A1(net294),
    .A2(_0994_),
    .B1(net234),
    .B2(_0996_),
    .C1(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__nor2_1 _1227_ (.A(_0987_),
    .B(net737),
    .Y(net413));
 sky130_fd_sc_hd__a22o_1 _1228_ (.A1(_0996_),
    .A2(net235),
    .B1(net333),
    .B2(_1002_),
    .X(_1005_));
 sky130_fd_sc_hd__a221oi_2 _1229_ (.A1(net295),
    .A2(_0994_),
    .B1(net288),
    .B2(_0998_),
    .C1(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__nor2_2 _1230_ (.A(_0987_),
    .B(net736),
    .Y(net424));
 sky130_fd_sc_hd__a22o_1 _1231_ (.A1(_0996_),
    .A2(net236),
    .B1(net334),
    .B2(_1002_),
    .X(_1007_));
 sky130_fd_sc_hd__a221oi_4 _1232_ (.A1(net296),
    .A2(_0994_),
    .B1(net299),
    .B2(_0998_),
    .C1(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__nor2_2 _1233_ (.A(_0987_),
    .B(_1008_),
    .Y(net435));
 sky130_fd_sc_hd__buf_8 _1234_ (.A(_1002_),
    .X(_1009_));
 sky130_fd_sc_hd__inv_2 _1235_ (.A(_0988_),
    .Y(_1010_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(_1010_),
    .B(net310),
    .Y(_1011_));
 sky130_fd_sc_hd__nand2_1 _1237_ (.A(_0988_),
    .B(net297),
    .Y(_1012_));
 sky130_fd_sc_hd__buf_8 _1238_ (.A(net770),
    .X(_1013_));
 sky130_fd_sc_hd__a21oi_1 _1239_ (.A1(_1011_),
    .A2(_1012_),
    .B1(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__a221oi_2 _1240_ (.A1(net237),
    .A2(_0996_),
    .B1(net335),
    .B2(_1009_),
    .C1(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__nor2_1 _1241_ (.A(_0987_),
    .B(net735),
    .Y(net446));
 sky130_fd_sc_hd__nand2_1 _1242_ (.A(_1010_),
    .B(net321),
    .Y(_1016_));
 sky130_fd_sc_hd__nand2_1 _1243_ (.A(_0988_),
    .B(net298),
    .Y(_1017_));
 sky130_fd_sc_hd__a21oi_1 _1244_ (.A1(_1016_),
    .A2(_1017_),
    .B1(_1013_),
    .Y(_1018_));
 sky130_fd_sc_hd__a221oi_2 _1245_ (.A1(net238),
    .A2(_0996_),
    .B1(net336),
    .B2(_0991_),
    .C1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_2 _1246_ (.A(_0987_),
    .B(net734),
    .Y(net457));
 sky130_fd_sc_hd__buf_8 _1247_ (.A(_0992_),
    .X(_1020_));
 sky130_fd_sc_hd__clkinv_4 _1248_ (.A(_0998_),
    .Y(_1021_));
 sky130_fd_sc_hd__buf_8 _1249_ (.A(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__o22ai_2 _1250_ (.A1(net300),
    .A2(_1020_),
    .B1(net332),
    .B2(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__buf_12 _1251_ (.A(_0995_),
    .X(_1024_));
 sky130_fd_sc_hd__clkinv_4 _1252_ (.A(_0990_),
    .Y(_1025_));
 sky130_fd_sc_hd__buf_8 _1253_ (.A(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__o22ai_4 _1254_ (.A1(net239),
    .A2(_1024_),
    .B1(net337),
    .B2(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_4 _1255_ (.A(_1023_),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__clkbuf_4 _1256_ (.A(_0986_),
    .X(_1029_));
 sky130_fd_sc_hd__and2_1 _1257_ (.A(_1028_),
    .B(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__buf_1 _1258_ (.A(_1030_),
    .X(net468));
 sky130_fd_sc_hd__o22ai_2 _1259_ (.A1(net301),
    .A2(_1020_),
    .B1(net343),
    .B2(_1022_),
    .Y(_1031_));
 sky130_fd_sc_hd__o22ai_4 _1260_ (.A1(net240),
    .A2(_1024_),
    .B1(net338),
    .B2(_1026_),
    .Y(_1032_));
 sky130_fd_sc_hd__nor2_4 _1261_ (.A(_1031_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__and2_1 _1262_ (.A(_1033_),
    .B(_1029_),
    .X(_1034_));
 sky130_fd_sc_hd__buf_1 _1263_ (.A(_1034_),
    .X(net479));
 sky130_fd_sc_hd__o22ai_2 _1264_ (.A1(net302),
    .A2(_1020_),
    .B1(net354),
    .B2(_1022_),
    .Y(_1035_));
 sky130_fd_sc_hd__buf_12 _1265_ (.A(_1025_),
    .X(_1036_));
 sky130_fd_sc_hd__o22ai_4 _1266_ (.A1(net242),
    .A2(_1024_),
    .B1(net339),
    .B2(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__nor2_4 _1267_ (.A(_1035_),
    .B(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__and2_1 _1268_ (.A(_1038_),
    .B(_1029_),
    .X(_1039_));
 sky130_fd_sc_hd__buf_1 _1269_ (.A(_1039_),
    .X(net490));
 sky130_fd_sc_hd__o22ai_2 _1270_ (.A1(net303),
    .A2(_1020_),
    .B1(net365),
    .B2(_1022_),
    .Y(_1040_));
 sky130_fd_sc_hd__o22ai_4 _1271_ (.A1(net243),
    .A2(_1024_),
    .B1(net340),
    .B2(_1036_),
    .Y(_1041_));
 sky130_fd_sc_hd__nor2_4 _1272_ (.A(_1040_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__and2_1 _1273_ (.A(_1042_),
    .B(_1029_),
    .X(_1043_));
 sky130_fd_sc_hd__buf_1 _1274_ (.A(_1043_),
    .X(net501));
 sky130_fd_sc_hd__o22ai_2 _1275_ (.A1(net304),
    .A2(_1020_),
    .B1(net241),
    .B2(_1022_),
    .Y(_1044_));
 sky130_fd_sc_hd__o22ai_4 _1276_ (.A1(net244),
    .A2(_1024_),
    .B1(net341),
    .B2(_1036_),
    .Y(_1045_));
 sky130_fd_sc_hd__nor2_4 _1277_ (.A(_1044_),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__and2_1 _1278_ (.A(_1046_),
    .B(_1029_),
    .X(_1047_));
 sky130_fd_sc_hd__buf_1 _1279_ (.A(_1047_),
    .X(net377));
 sky130_fd_sc_hd__o22ai_2 _1280_ (.A1(net305),
    .A2(_1020_),
    .B1(net252),
    .B2(_1022_),
    .Y(_1048_));
 sky130_fd_sc_hd__o22ai_4 _1281_ (.A1(net245),
    .A2(_1024_),
    .B1(net342),
    .B2(_1036_),
    .Y(_1049_));
 sky130_fd_sc_hd__nor2_4 _1282_ (.A(_1048_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__and2_1 _1283_ (.A(_1050_),
    .B(_1029_),
    .X(_1051_));
 sky130_fd_sc_hd__buf_1 _1284_ (.A(_1051_),
    .X(net388));
 sky130_fd_sc_hd__o22ai_2 _1285_ (.A1(net306),
    .A2(_1020_),
    .B1(net263),
    .B2(_1022_),
    .Y(_1052_));
 sky130_fd_sc_hd__o22ai_4 _1286_ (.A1(net246),
    .A2(_1024_),
    .B1(net344),
    .B2(_1036_),
    .Y(_1053_));
 sky130_fd_sc_hd__nor2_4 _1287_ (.A(_1052_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__and2_1 _1288_ (.A(_1054_),
    .B(_1029_),
    .X(_1055_));
 sky130_fd_sc_hd__buf_1 _1289_ (.A(_1055_),
    .X(net399));
 sky130_fd_sc_hd__o22ai_2 _1290_ (.A1(net307),
    .A2(_1020_),
    .B1(net270),
    .B2(_1022_),
    .Y(_1056_));
 sky130_fd_sc_hd__o22ai_4 _1291_ (.A1(net247),
    .A2(_1024_),
    .B1(net345),
    .B2(_1036_),
    .Y(_1057_));
 sky130_fd_sc_hd__nor2_4 _1292_ (.A(_1056_),
    .B(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__and2_1 _1293_ (.A(_1058_),
    .B(_1029_),
    .X(_1059_));
 sky130_fd_sc_hd__buf_1 _1294_ (.A(_1059_),
    .X(net406));
 sky130_fd_sc_hd__buf_8 _1295_ (.A(_0992_),
    .X(_1060_));
 sky130_fd_sc_hd__buf_8 _1296_ (.A(_1021_),
    .X(_1061_));
 sky130_fd_sc_hd__o22ai_2 _1297_ (.A1(net308),
    .A2(_1060_),
    .B1(net271),
    .B2(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__o22ai_4 _1298_ (.A1(net248),
    .A2(_1024_),
    .B1(net346),
    .B2(_1036_),
    .Y(_1063_));
 sky130_fd_sc_hd__nor2_4 _1299_ (.A(_1062_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__and2_1 _1300_ (.A(_1064_),
    .B(_1029_),
    .X(_1065_));
 sky130_fd_sc_hd__buf_1 _1301_ (.A(_1065_),
    .X(net407));
 sky130_fd_sc_hd__o22ai_2 _1302_ (.A1(net309),
    .A2(_1060_),
    .B1(net272),
    .B2(_1061_),
    .Y(_1066_));
 sky130_fd_sc_hd__o22ai_4 _1303_ (.A1(net249),
    .A2(_1024_),
    .B1(net347),
    .B2(_1036_),
    .Y(_1067_));
 sky130_fd_sc_hd__nor2_4 _1304_ (.A(_1066_),
    .B(_1067_),
    .Y(_1068_));
 sky130_fd_sc_hd__and2_1 _1305_ (.A(_1068_),
    .B(_1029_),
    .X(_1069_));
 sky130_fd_sc_hd__buf_1 _1306_ (.A(_1069_),
    .X(net408));
 sky130_fd_sc_hd__o22ai_2 _1307_ (.A1(net311),
    .A2(_1060_),
    .B1(net273),
    .B2(_1061_),
    .Y(_1070_));
 sky130_fd_sc_hd__o22ai_4 _1308_ (.A1(net250),
    .A2(_1024_),
    .B1(net348),
    .B2(_1036_),
    .Y(_1071_));
 sky130_fd_sc_hd__nor2_4 _1309_ (.A(_1070_),
    .B(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__and2_1 _1310_ (.A(_1072_),
    .B(_1029_),
    .X(_1073_));
 sky130_fd_sc_hd__buf_1 _1311_ (.A(_1073_),
    .X(net409));
 sky130_fd_sc_hd__o22ai_2 _1312_ (.A1(net312),
    .A2(_1060_),
    .B1(net274),
    .B2(_1061_),
    .Y(_1074_));
 sky130_fd_sc_hd__o22ai_4 _1313_ (.A1(net251),
    .A2(_1024_),
    .B1(net349),
    .B2(_1036_),
    .Y(_1075_));
 sky130_fd_sc_hd__nor2_4 _1314_ (.A(_1074_),
    .B(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__and2_1 _1315_ (.A(_1076_),
    .B(_1029_),
    .X(_1077_));
 sky130_fd_sc_hd__buf_1 _1316_ (.A(_1077_),
    .X(net410));
 sky130_fd_sc_hd__inv_2 _1317_ (.A(net759),
    .Y(_1078_));
 sky130_fd_sc_hd__nor2_1 _1318_ (.A(net768),
    .B(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__inv_4 _1319_ (.A(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__nor2_8 _1320_ (.A(\arbiter.slave_handled[1] ),
    .B(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__clkinv_4 _1321_ (.A(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__clkbuf_16 _1322_ (.A(net768),
    .X(_1083_));
 sky130_fd_sc_hd__nand2_4 _1323_ (.A(_0993_),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__nand2_1 _1324_ (.A(_1082_),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__inv_2 _1325_ (.A(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__nand2_4 _1326_ (.A(_0982_),
    .B(_0983_),
    .Y(_1087_));
 sky130_fd_sc_hd__inv_4 _1327_ (.A(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__buf_12 _1328_ (.A(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__inv_4 _1329_ (.A(_0983_),
    .Y(_1090_));
 sky130_fd_sc_hd__nor2_4 _1330_ (.A(_0982_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__buf_12 _1331_ (.A(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__a22oi_4 _1332_ (.A1(_1089_),
    .A2(net80),
    .B1(net17),
    .B2(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__buf_6 _1333_ (.A(_0984_),
    .X(_1094_));
 sky130_fd_sc_hd__inv_6 _1334_ (.A(_0982_),
    .Y(_1095_));
 sky130_fd_sc_hd__nor2_8 _1335_ (.A(_0983_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__buf_8 _1336_ (.A(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__a22oi_1 _1337_ (.A1(_1094_),
    .A2(net1),
    .B1(_1097_),
    .B2(net181),
    .Y(_1098_));
 sky130_fd_sc_hd__nand2_2 _1338_ (.A(_1093_),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__inv_2 _1339_ (.A(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__nor2_1 _1340_ (.A(_1086_),
    .B(_1100_),
    .Y(net682));
 sky130_fd_sc_hd__buf_6 _1341_ (.A(_0988_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_8 _1342_ (.A(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__buf_6 _1343_ (.A(_1095_),
    .X(_1103_));
 sky130_fd_sc_hd__nand2_1 _1344_ (.A(_1103_),
    .B(net112),
    .Y(_1104_));
 sky130_fd_sc_hd__buf_6 _1345_ (.A(_0982_),
    .X(_1105_));
 sky130_fd_sc_hd__nand2_1 _1346_ (.A(_1105_),
    .B(net182),
    .Y(_1106_));
 sky130_fd_sc_hd__nand2_1 _1347_ (.A(_1104_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__clkbuf_8 _1348_ (.A(_1090_),
    .X(_1108_));
 sky130_fd_sc_hd__buf_6 _1349_ (.A(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__nand2_1 _1350_ (.A(_1107_),
    .B(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(_1103_),
    .B(net18),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_1 _1352_ (.A(_1105_),
    .B(net81),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_1 _1353_ (.A(_1111_),
    .B(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__buf_4 _1354_ (.A(_0983_),
    .X(_1114_));
 sky130_fd_sc_hd__nand2_1 _1355_ (.A(_1113_),
    .B(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__nand2_4 _1356_ (.A(_1110_),
    .B(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__inv_2 _1357_ (.A(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__nor2_1 _1358_ (.A(_1082_),
    .B(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__a41o_1 _1359_ (.A1(_1083_),
    .A2(_1102_),
    .A3(_1116_),
    .A4(_0989_),
    .B1(_1118_),
    .X(net683));
 sky130_fd_sc_hd__nand3_1 _1360_ (.A(_1116_),
    .B(_1010_),
    .C(\arbiter.slave_sel[0][1] ),
    .Y(_1119_));
 sky130_fd_sc_hd__buf_6 _1361_ (.A(_1095_),
    .X(_1120_));
 sky130_fd_sc_hd__nand2_1 _1362_ (.A(_1120_),
    .B(net151),
    .Y(_1121_));
 sky130_fd_sc_hd__buf_6 _1363_ (.A(_0982_),
    .X(_1122_));
 sky130_fd_sc_hd__nand2_1 _1364_ (.A(_1122_),
    .B(net183),
    .Y(_1123_));
 sky130_fd_sc_hd__nand2_1 _1365_ (.A(_1121_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__nand2_1 _1366_ (.A(_1124_),
    .B(_1109_),
    .Y(_1125_));
 sky130_fd_sc_hd__nand2_1 _1367_ (.A(_1120_),
    .B(net19),
    .Y(_1126_));
 sky130_fd_sc_hd__nand2_1 _1368_ (.A(_1122_),
    .B(net82),
    .Y(_1127_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(_1126_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__nand2_1 _1370_ (.A(_1128_),
    .B(_1114_),
    .Y(_1129_));
 sky130_fd_sc_hd__nand2_4 _1371_ (.A(_1125_),
    .B(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand3_1 _1372_ (.A(_1130_),
    .B(_1101_),
    .C(_1021_),
    .Y(_1131_));
 sky130_fd_sc_hd__nand2_1 _1373_ (.A(_1119_),
    .B(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__nor2_2 _1374_ (.A(_0998_),
    .B(_0996_),
    .Y(_1133_));
 sky130_fd_sc_hd__buf_4 _1375_ (.A(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_1132_),
    .B(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__clkbuf_8 _1377_ (.A(_0996_),
    .X(_1136_));
 sky130_fd_sc_hd__nand2_1 _1378_ (.A(_1099_),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__a21o_1 _1379_ (.A1(_1135_),
    .A2(_1137_),
    .B1(_1084_),
    .X(_1138_));
 sky130_fd_sc_hd__buf_4 _1380_ (.A(_1081_),
    .X(_1139_));
 sky130_fd_sc_hd__nand2_1 _1381_ (.A(_1130_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_2 _1382_ (.A(_1138_),
    .B(_1140_),
    .Y(net684));
 sky130_fd_sc_hd__nand2_1 _1383_ (.A(_1130_),
    .B(_1061_),
    .Y(_1141_));
 sky130_fd_sc_hd__buf_8 _1384_ (.A(_1010_),
    .X(_1142_));
 sky130_fd_sc_hd__buf_6 _1385_ (.A(_1095_),
    .X(_1143_));
 sky130_fd_sc_hd__nand2_1 _1386_ (.A(_1143_),
    .B(net162),
    .Y(_1144_));
 sky130_fd_sc_hd__buf_6 _1387_ (.A(_0982_),
    .X(_1145_));
 sky130_fd_sc_hd__nand2_1 _1388_ (.A(_1145_),
    .B(net185),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _1389_ (.A(_1144_),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _1390_ (.A(_1147_),
    .B(_1108_),
    .Y(_1148_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(_1143_),
    .B(net20),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _1392_ (.A(_1145_),
    .B(net83),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(_1149_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand2_1 _1394_ (.A(_1151_),
    .B(_0983_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_4 _1395_ (.A(_1148_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__nor2_1 _1396_ (.A(_1020_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__a21oi_1 _1397_ (.A1(_1141_),
    .A2(_1142_),
    .B1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__o21bai_1 _1398_ (.A1(_1010_),
    .A2(_1116_),
    .B1_N(_0989_),
    .Y(_1156_));
 sky130_fd_sc_hd__nand2_1 _1399_ (.A(_1156_),
    .B(_1020_),
    .Y(_1157_));
 sky130_fd_sc_hd__nand2_1 _1400_ (.A(_1155_),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__nand2_1 _1401_ (.A(_1158_),
    .B(_1026_),
    .Y(_1159_));
 sky130_fd_sc_hd__inv_2 _1402_ (.A(_1084_),
    .Y(_1160_));
 sky130_fd_sc_hd__clkbuf_8 _1403_ (.A(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(_1143_),
    .B(net12),
    .Y(_1162_));
 sky130_fd_sc_hd__nand2_1 _1405_ (.A(_1145_),
    .B(net192),
    .Y(_1163_));
 sky130_fd_sc_hd__nand2_1 _1406_ (.A(_1162_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__nand2_1 _1407_ (.A(_1164_),
    .B(_1108_),
    .Y(_1165_));
 sky130_fd_sc_hd__nand2_1 _1408_ (.A(_1143_),
    .B(net28),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _1409_ (.A(_1145_),
    .B(net91),
    .Y(_1167_));
 sky130_fd_sc_hd__nand2_1 _1410_ (.A(_1166_),
    .B(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__nand2_2 _1411_ (.A(_1168_),
    .B(_0983_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand3_1 _1412_ (.A(_1165_),
    .B(_1169_),
    .C(_1002_),
    .Y(_1170_));
 sky130_fd_sc_hd__nand3_1 _1413_ (.A(_1159_),
    .B(_1161_),
    .C(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _1414_ (.A(_1153_),
    .B(_1139_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_2 _1415_ (.A(_1171_),
    .B(_1172_),
    .Y(net686));
 sky130_fd_sc_hd__nand2_2 _1416_ (.A(_1132_),
    .B(_1136_),
    .Y(_1173_));
 sky130_fd_sc_hd__nand2_1 _1417_ (.A(_1143_),
    .B(net173),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_1 _1418_ (.A(_1145_),
    .B(net186),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _1419_ (.A(_1174_),
    .B(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _1420_ (.A(_1176_),
    .B(_1108_),
    .Y(_1177_));
 sky130_fd_sc_hd__nand2_1 _1421_ (.A(_1143_),
    .B(net21),
    .Y(_1178_));
 sky130_fd_sc_hd__nand2_1 _1422_ (.A(_1145_),
    .B(net84),
    .Y(_1179_));
 sky130_fd_sc_hd__nand2_1 _1423_ (.A(_1178_),
    .B(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__nand2_1 _1424_ (.A(_1180_),
    .B(_1114_),
    .Y(_1181_));
 sky130_fd_sc_hd__nand2_4 _1425_ (.A(_1177_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__nand2_1 _1426_ (.A(_1182_),
    .B(_1101_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _1427_ (.A(_1153_),
    .B(_1002_),
    .Y(_1184_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(_1183_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(_1185_),
    .B(_1134_),
    .Y(_1186_));
 sky130_fd_sc_hd__nand3_1 _1430_ (.A(_1173_),
    .B(_1026_),
    .C(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__buf_4 _1431_ (.A(_1160_),
    .X(_1188_));
 sky130_fd_sc_hd__nand2_1 _1432_ (.A(_1103_),
    .B(net23),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _1433_ (.A(_1105_),
    .B(net193),
    .Y(_1190_));
 sky130_fd_sc_hd__nand2_1 _1434_ (.A(_1189_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand2_2 _1435_ (.A(_1191_),
    .B(_1109_),
    .Y(_1192_));
 sky130_fd_sc_hd__nand2_1 _1436_ (.A(_1103_),
    .B(net29),
    .Y(_1193_));
 sky130_fd_sc_hd__nand2_1 _1437_ (.A(_1105_),
    .B(net92),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _1438_ (.A(_1193_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand2_2 _1439_ (.A(_1195_),
    .B(_1114_),
    .Y(_1196_));
 sky130_fd_sc_hd__nand2_2 _1440_ (.A(_1192_),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__inv_2 _1441_ (.A(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__nand2_1 _1442_ (.A(_1198_),
    .B(_1009_),
    .Y(_1199_));
 sky130_fd_sc_hd__nand3_1 _1443_ (.A(_1187_),
    .B(_1188_),
    .C(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nand2_1 _1444_ (.A(_1182_),
    .B(_1139_),
    .Y(_0014_));
 sky130_fd_sc_hd__nand2_2 _1445_ (.A(_1200_),
    .B(_0014_),
    .Y(net687));
 sky130_fd_sc_hd__buf_4 _1446_ (.A(_1083_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_6 _1447_ (.A(_1088_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_12 _1448_ (.A(_1091_),
    .X(_0017_));
 sky130_fd_sc_hd__a22oi_4 _1449_ (.A1(_0016_),
    .A2(net85),
    .B1(net22),
    .B2(_0017_),
    .Y(_0018_));
 sky130_fd_sc_hd__a22oi_2 _1450_ (.A1(_1094_),
    .A2(net184),
    .B1(_1097_),
    .B2(net187),
    .Y(_0019_));
 sky130_fd_sc_hd__nand2_4 _1451_ (.A(_0018_),
    .B(_0019_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_6 _1452_ (.A(_1082_),
    .X(_0021_));
 sky130_fd_sc_hd__clkinv_4 _1453_ (.A(_0020_),
    .Y(_0022_));
 sky130_fd_sc_hd__nor2_1 _1454_ (.A(_0021_),
    .B(_0022_),
    .Y(_0023_));
 sky130_fd_sc_hd__a31o_1 _1455_ (.A1(_0015_),
    .A2(_0994_),
    .A3(_0020_),
    .B1(_0023_),
    .X(net688));
 sky130_fd_sc_hd__nand2_1 _1456_ (.A(_1120_),
    .B(net24),
    .Y(_0024_));
 sky130_fd_sc_hd__nand2_1 _1457_ (.A(_1122_),
    .B(net86),
    .Y(_0025_));
 sky130_fd_sc_hd__a21o_1 _1458_ (.A1(_0024_),
    .A2(_0025_),
    .B1(_1108_),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _1459_ (.A(_1120_),
    .B(net195),
    .Y(_0027_));
 sky130_fd_sc_hd__nand2_1 _1460_ (.A(_1122_),
    .B(net188),
    .Y(_0028_));
 sky130_fd_sc_hd__nand2_1 _1461_ (.A(_0027_),
    .B(_0028_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand2_1 _1462_ (.A(_0029_),
    .B(_1109_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_2 _1463_ (.A(_0026_),
    .B(_0030_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1464_ (.A(_0031_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2_1 _1465_ (.A(_0020_),
    .B(_1009_),
    .Y(_0033_));
 sky130_fd_sc_hd__clkbuf_8 _1466_ (.A(_1133_),
    .X(_0034_));
 sky130_fd_sc_hd__buf_4 _1467_ (.A(_0988_),
    .X(_0035_));
 sky130_fd_sc_hd__nand2_1 _1468_ (.A(_0031_),
    .B(_0035_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand3_1 _1469_ (.A(_0033_),
    .B(_0034_),
    .C(_0036_),
    .Y(_0037_));
 sky130_fd_sc_hd__or2_1 _1470_ (.A(_1024_),
    .B(_1185_),
    .X(_0038_));
 sky130_fd_sc_hd__nand3_1 _1471_ (.A(_0037_),
    .B(_0038_),
    .C(_1188_),
    .Y(_0039_));
 sky130_fd_sc_hd__o21ai_2 _1472_ (.A1(_0021_),
    .A2(_0032_),
    .B1(_0039_),
    .Y(net689));
 sky130_fd_sc_hd__nand2_1 _1473_ (.A(_0031_),
    .B(_0991_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand2_1 _1474_ (.A(_1120_),
    .B(net206),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _1475_ (.A(_1122_),
    .B(net189),
    .Y(_0042_));
 sky130_fd_sc_hd__nand2_1 _1476_ (.A(_0041_),
    .B(_0042_),
    .Y(_0043_));
 sky130_fd_sc_hd__nand2_1 _1477_ (.A(_0043_),
    .B(_1109_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(_1092_),
    .B(net25),
    .Y(_0045_));
 sky130_fd_sc_hd__nand2_1 _1479_ (.A(_1089_),
    .B(net87),
    .Y(_0046_));
 sky130_fd_sc_hd__nand3_4 _1480_ (.A(_0044_),
    .B(_0045_),
    .C(_0046_),
    .Y(_0047_));
 sky130_fd_sc_hd__nand2_1 _1481_ (.A(_0047_),
    .B(_0035_),
    .Y(_0048_));
 sky130_fd_sc_hd__nand2_1 _1482_ (.A(_0040_),
    .B(_0048_),
    .Y(_0049_));
 sky130_fd_sc_hd__nand2_1 _1483_ (.A(_0049_),
    .B(_0034_),
    .Y(_0050_));
 sky130_fd_sc_hd__nand2_1 _1484_ (.A(_0020_),
    .B(_1136_),
    .Y(_0051_));
 sky130_fd_sc_hd__nand3_1 _1485_ (.A(_0050_),
    .B(_1026_),
    .C(_0051_),
    .Y(_0052_));
 sky130_fd_sc_hd__a22oi_2 _1486_ (.A1(_0984_),
    .A2(net56),
    .B1(_1097_),
    .B2(net197),
    .Y(_0053_));
 sky130_fd_sc_hd__nand2_1 _1487_ (.A(_0017_),
    .B(net32),
    .Y(_0054_));
 sky130_fd_sc_hd__nand2_1 _1488_ (.A(_0016_),
    .B(net95),
    .Y(_0055_));
 sky130_fd_sc_hd__and2_2 _1489_ (.A(_0054_),
    .B(_0055_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_4 _1490_ (.A(_0053_),
    .B(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__clkinv_4 _1491_ (.A(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__nand3_1 _1492_ (.A(_0058_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0059_));
 sky130_fd_sc_hd__nand3_1 _1493_ (.A(_0052_),
    .B(_1188_),
    .C(_0059_),
    .Y(_0060_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(_0047_),
    .B(_1139_),
    .Y(_0061_));
 sky130_fd_sc_hd__nand2_2 _1495_ (.A(_0060_),
    .B(_0061_),
    .Y(net690));
 sky130_fd_sc_hd__nand2_1 _1496_ (.A(_1120_),
    .B(net217),
    .Y(_0062_));
 sky130_fd_sc_hd__nand2_1 _1497_ (.A(_1122_),
    .B(net190),
    .Y(_0063_));
 sky130_fd_sc_hd__nand2_1 _1498_ (.A(_0062_),
    .B(_0063_),
    .Y(_0064_));
 sky130_fd_sc_hd__nand2_1 _1499_ (.A(_0064_),
    .B(_1109_),
    .Y(_0065_));
 sky130_fd_sc_hd__nand2_1 _1500_ (.A(_1103_),
    .B(net26),
    .Y(_0066_));
 sky130_fd_sc_hd__nand2_1 _1501_ (.A(_1105_),
    .B(net88),
    .Y(_0067_));
 sky130_fd_sc_hd__nand2_1 _1502_ (.A(_0066_),
    .B(_0067_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand2_1 _1503_ (.A(_0068_),
    .B(_1114_),
    .Y(_0069_));
 sky130_fd_sc_hd__nand2_4 _1504_ (.A(_0065_),
    .B(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1505_ (.A(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__nand2_1 _1506_ (.A(_0047_),
    .B(_0991_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand2_1 _1507_ (.A(_0070_),
    .B(_1101_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand3_1 _1508_ (.A(_0072_),
    .B(_1134_),
    .C(_0073_),
    .Y(_0074_));
 sky130_fd_sc_hd__nand2_1 _1509_ (.A(_0036_),
    .B(_1020_),
    .Y(_0075_));
 sky130_fd_sc_hd__nand2_1 _1510_ (.A(_0074_),
    .B(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__a22oi_4 _1511_ (.A1(_0016_),
    .A2(net96),
    .B1(net33),
    .B2(_0017_),
    .Y(_0077_));
 sky130_fd_sc_hd__a22oi_2 _1512_ (.A1(_1094_),
    .A2(net67),
    .B1(_1097_),
    .B2(net198),
    .Y(_0078_));
 sky130_fd_sc_hd__nand2_4 _1513_ (.A(_0077_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__nand3_2 _1514_ (.A(_0079_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0080_));
 sky130_fd_sc_hd__nand2_1 _1515_ (.A(_0076_),
    .B(_0080_),
    .Y(_0081_));
 sky130_fd_sc_hd__nand2_1 _1516_ (.A(_0081_),
    .B(_1161_),
    .Y(_0082_));
 sky130_fd_sc_hd__o21ai_2 _1517_ (.A1(_0021_),
    .A2(_0071_),
    .B1(_0082_),
    .Y(net691));
 sky130_fd_sc_hd__nand2_1 _1518_ (.A(_1143_),
    .B(net228),
    .Y(_0083_));
 sky130_fd_sc_hd__nand2_1 _1519_ (.A(_1145_),
    .B(net191),
    .Y(_0084_));
 sky130_fd_sc_hd__nand2_1 _1520_ (.A(_0083_),
    .B(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__nand2_1 _1521_ (.A(_0085_),
    .B(_1108_),
    .Y(_0086_));
 sky130_fd_sc_hd__nand2_1 _1522_ (.A(_1143_),
    .B(net27),
    .Y(_0087_));
 sky130_fd_sc_hd__nand2_1 _1523_ (.A(_1145_),
    .B(net90),
    .Y(_0088_));
 sky130_fd_sc_hd__nand2_1 _1524_ (.A(_0087_),
    .B(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__nand2_1 _1525_ (.A(_0089_),
    .B(_1114_),
    .Y(_0090_));
 sky130_fd_sc_hd__nand2_2 _1526_ (.A(_0086_),
    .B(_0090_),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1527_ (.A(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1528_ (.A(_1133_),
    .Y(_0093_));
 sky130_fd_sc_hd__clkbuf_8 _1529_ (.A(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__nand2_1 _1530_ (.A(_0070_),
    .B(_1002_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_1 _1531_ (.A(_0091_),
    .B(_1101_),
    .Y(_0096_));
 sky130_fd_sc_hd__nand2_2 _1532_ (.A(_0095_),
    .B(_0096_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand3_1 _1533_ (.A(_0040_),
    .B(_0048_),
    .C(_0094_),
    .Y(_0098_));
 sky130_fd_sc_hd__o21ai_4 _1534_ (.A1(_0094_),
    .A2(_0097_),
    .B1(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__o22ai_4 _1535_ (.A1(_1082_),
    .A2(_0092_),
    .B1(_1084_),
    .B2(_0099_),
    .Y(net692));
 sky130_fd_sc_hd__o22ai_2 _1536_ (.A1(net313),
    .A2(_1060_),
    .B1(net275),
    .B2(_1061_),
    .Y(_0100_));
 sky130_fd_sc_hd__o22ai_4 _1537_ (.A1(net253),
    .A2(_1024_),
    .B1(net350),
    .B2(_1036_),
    .Y(_0101_));
 sky130_fd_sc_hd__nor2_4 _1538_ (.A(_0100_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__and2_1 _1539_ (.A(_0102_),
    .B(_1029_),
    .X(_0103_));
 sky130_fd_sc_hd__buf_1 _1540_ (.A(_0103_),
    .X(net411));
 sky130_fd_sc_hd__nand2_1 _1541_ (.A(_0091_),
    .B(_1021_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _1542_ (.A(_0104_),
    .B(_1142_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2_1 _1543_ (.A(_1165_),
    .B(_1169_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand2_1 _1544_ (.A(_0106_),
    .B(_1021_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_1 _1545_ (.A(_0107_),
    .B(_1101_),
    .Y(_0108_));
 sky130_fd_sc_hd__nand2_1 _1546_ (.A(_0105_),
    .B(_0108_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(_0109_),
    .B(_1134_),
    .Y(_0110_));
 sky130_fd_sc_hd__nand2_1 _1548_ (.A(_0073_),
    .B(_1020_),
    .Y(_0111_));
 sky130_fd_sc_hd__nand2_1 _1549_ (.A(_0110_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__a22oi_4 _1550_ (.A1(_1089_),
    .A2(net98),
    .B1(net36),
    .B2(_1092_),
    .Y(_0113_));
 sky130_fd_sc_hd__a22oi_2 _1551_ (.A1(_1094_),
    .A2(net89),
    .B1(_1097_),
    .B2(net200),
    .Y(_0114_));
 sky130_fd_sc_hd__nand2_4 _1552_ (.A(_0113_),
    .B(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__nand2_1 _1553_ (.A(_0115_),
    .B(_1009_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand2_1 _1554_ (.A(_0112_),
    .B(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__nand2_1 _1555_ (.A(_0117_),
    .B(_1161_),
    .Y(_0118_));
 sky130_fd_sc_hd__nand2_1 _1556_ (.A(_0106_),
    .B(_1139_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_2 _1557_ (.A(_0118_),
    .B(_0119_),
    .Y(net693));
 sky130_fd_sc_hd__inv_2 _1558_ (.A(net100),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1559_ (.A(net201),
    .Y(_0121_));
 sky130_fd_sc_hd__nand2_4 _1560_ (.A(_1108_),
    .B(_1105_),
    .Y(_0122_));
 sky130_fd_sc_hd__a22oi_4 _1561_ (.A1(_0016_),
    .A2(net99),
    .B1(net37),
    .B2(_0017_),
    .Y(_0123_));
 sky130_fd_sc_hd__o221ai_4 _1562_ (.A1(_0120_),
    .A2(_0985_),
    .B1(_0121_),
    .B2(_0122_),
    .C1(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__buf_6 _1563_ (.A(_0991_),
    .X(_0125_));
 sky130_fd_sc_hd__nand2_1 _1564_ (.A(_0124_),
    .B(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand3_1 _1565_ (.A(_1192_),
    .B(_1196_),
    .C(_0993_),
    .Y(_0127_));
 sky130_fd_sc_hd__nand2_1 _1566_ (.A(_0127_),
    .B(_1170_),
    .Y(_0128_));
 sky130_fd_sc_hd__nand3_1 _1567_ (.A(_0095_),
    .B(_0096_),
    .C(_0093_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand3b_1 _1568_ (.A_N(_0128_),
    .B(_0129_),
    .C(_1026_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_1 _1569_ (.A(_0126_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand2_1 _1570_ (.A(_0131_),
    .B(_1161_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_1 _1571_ (.A(_1197_),
    .B(_1139_),
    .Y(_0133_));
 sky130_fd_sc_hd__nand2_2 _1572_ (.A(_0132_),
    .B(_0133_),
    .Y(net694));
 sky130_fd_sc_hd__a22oi_2 _1573_ (.A1(_1094_),
    .A2(net34),
    .B1(_1097_),
    .B2(net194),
    .Y(_0134_));
 sky130_fd_sc_hd__nand2_1 _1574_ (.A(_1120_),
    .B(net30),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _1575_ (.A(_1122_),
    .B(net93),
    .Y(_0136_));
 sky130_fd_sc_hd__a21o_1 _1576_ (.A1(_0135_),
    .A2(_0136_),
    .B1(_1108_),
    .X(_0137_));
 sky130_fd_sc_hd__nand2_2 _1577_ (.A(_0134_),
    .B(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1578_ (.A(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__nand2_1 _1579_ (.A(_0139_),
    .B(_0994_),
    .Y(_0140_));
 sky130_fd_sc_hd__nor2_1 _1580_ (.A(_0021_),
    .B(_0139_),
    .Y(_0141_));
 sky130_fd_sc_hd__a31o_1 _1581_ (.A1(_0140_),
    .A2(_1160_),
    .A3(_1199_),
    .B1(_0141_),
    .X(net695));
 sky130_fd_sc_hd__a22oi_2 _1582_ (.A1(_1094_),
    .A2(net45),
    .B1(_1097_),
    .B2(net196),
    .Y(_0142_));
 sky130_fd_sc_hd__and2b_1 _1583_ (.A_N(_1087_),
    .B(net94),
    .X(_0143_));
 sky130_fd_sc_hd__a21oi_4 _1584_ (.A1(_0017_),
    .A2(net31),
    .B1(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__nand2_4 _1585_ (.A(_0142_),
    .B(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1586_ (.A(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__nand3_1 _1587_ (.A(_0145_),
    .B(_1102_),
    .C(_1022_),
    .Y(_0147_));
 sky130_fd_sc_hd__nand3_1 _1588_ (.A(_0138_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0148_));
 sky130_fd_sc_hd__nand2_1 _1589_ (.A(_0147_),
    .B(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__nand3_1 _1590_ (.A(_0149_),
    .B(_0015_),
    .C(_0994_),
    .Y(_0150_));
 sky130_fd_sc_hd__o21ai_2 _1591_ (.A1(_0021_),
    .A2(_0146_),
    .B1(_0150_),
    .Y(net697));
 sky130_fd_sc_hd__o21ai_1 _1592_ (.A1(_1013_),
    .A2(_0057_),
    .B1(_1102_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand2_1 _1593_ (.A(_1095_),
    .B(net134),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_1 _1594_ (.A(_0982_),
    .B(net204),
    .Y(_0153_));
 sky130_fd_sc_hd__nand2_1 _1595_ (.A(_0152_),
    .B(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__nand2_1 _1596_ (.A(_0154_),
    .B(_1090_),
    .Y(_0155_));
 sky130_fd_sc_hd__nand2_1 _1597_ (.A(_1095_),
    .B(net40),
    .Y(_0156_));
 sky130_fd_sc_hd__nand2_1 _1598_ (.A(_0982_),
    .B(net103),
    .Y(_0157_));
 sky130_fd_sc_hd__nand2_1 _1599_ (.A(_0156_),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__nand2_1 _1600_ (.A(_0158_),
    .B(_0983_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand2_4 _1601_ (.A(_0155_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _1602_ (.A(_0160_),
    .B(_1002_),
    .Y(_0161_));
 sky130_fd_sc_hd__nand2_1 _1603_ (.A(_0151_),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _1604_ (.A(_0162_),
    .B(_1161_),
    .Y(_0163_));
 sky130_fd_sc_hd__o21ai_2 _1605_ (.A1(_0021_),
    .A2(_0058_),
    .B1(_0163_),
    .Y(net698));
 sky130_fd_sc_hd__nand3_1 _1606_ (.A(_0079_),
    .B(_1102_),
    .C(_1022_),
    .Y(_0164_));
 sky130_fd_sc_hd__nand3_2 _1607_ (.A(_0057_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand3_1 _1608_ (.A(_0164_),
    .B(_0165_),
    .C(_0034_),
    .Y(_0166_));
 sky130_fd_sc_hd__o21a_1 _1609_ (.A1(_1024_),
    .A2(_0145_),
    .B1(_1022_),
    .X(_0167_));
 sky130_fd_sc_hd__nand3_1 _1610_ (.A(_0166_),
    .B(_0167_),
    .C(_1188_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2_1 _1611_ (.A(_0079_),
    .B(_1139_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_2 _1612_ (.A(_0168_),
    .B(_0169_),
    .Y(net699));
 sky130_fd_sc_hd__a22oi_2 _1613_ (.A1(_1094_),
    .A2(net78),
    .B1(_1097_),
    .B2(net199),
    .Y(_0170_));
 sky130_fd_sc_hd__nand2_1 _1614_ (.A(_0017_),
    .B(net35),
    .Y(_0171_));
 sky130_fd_sc_hd__nand2_1 _1615_ (.A(_0016_),
    .B(net97),
    .Y(_0172_));
 sky130_fd_sc_hd__and2_2 _1616_ (.A(_0171_),
    .B(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__nand2_4 _1617_ (.A(_0170_),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand3_1 _1618_ (.A(_0174_),
    .B(_1102_),
    .C(_1022_),
    .Y(_0175_));
 sky130_fd_sc_hd__nand3_1 _1619_ (.A(_0080_),
    .B(_0175_),
    .C(_0034_),
    .Y(_0176_));
 sky130_fd_sc_hd__nand3_2 _1620_ (.A(_0145_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0177_));
 sky130_fd_sc_hd__nand3_1 _1621_ (.A(_0057_),
    .B(_0035_),
    .C(_1021_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand3_1 _1622_ (.A(_0177_),
    .B(_0178_),
    .C(_0094_),
    .Y(_0179_));
 sky130_fd_sc_hd__nand3_1 _1623_ (.A(_0176_),
    .B(_0179_),
    .C(_1188_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_1 _1624_ (.A(_0174_),
    .B(_1139_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_2 _1625_ (.A(_0180_),
    .B(_0181_),
    .Y(net700));
 sky130_fd_sc_hd__nand3_1 _1626_ (.A(_0164_),
    .B(_0165_),
    .C(_0094_),
    .Y(_0182_));
 sky130_fd_sc_hd__nand3_2 _1627_ (.A(_0174_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand2_1 _1628_ (.A(_0115_),
    .B(_0035_),
    .Y(_0184_));
 sky130_fd_sc_hd__nand3_1 _1629_ (.A(_0183_),
    .B(_0034_),
    .C(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__nand3_1 _1630_ (.A(_0182_),
    .B(_0185_),
    .C(_1188_),
    .Y(_0186_));
 sky130_fd_sc_hd__nand2_1 _1631_ (.A(_0115_),
    .B(_1139_),
    .Y(_0187_));
 sky130_fd_sc_hd__nand2_2 _1632_ (.A(_0186_),
    .B(_0187_),
    .Y(net701));
 sky130_fd_sc_hd__inv_2 _1633_ (.A(_0124_),
    .Y(_0188_));
 sky130_fd_sc_hd__nand3_1 _1634_ (.A(_0124_),
    .B(_0015_),
    .C(_0994_),
    .Y(_0189_));
 sky130_fd_sc_hd__o21ai_2 _1635_ (.A1(_0021_),
    .A2(_0188_),
    .B1(_0189_),
    .Y(net702));
 sky130_fd_sc_hd__nand2_1 _1636_ (.A(_1096_),
    .B(net202),
    .Y(_0190_));
 sky130_fd_sc_hd__nand2_1 _1637_ (.A(_0984_),
    .B(net111),
    .Y(_0191_));
 sky130_fd_sc_hd__and2_1 _1638_ (.A(_0190_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _1639_ (.A(_0017_),
    .B(net38),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_1 _1640_ (.A(_0016_),
    .B(net101),
    .Y(_0194_));
 sky130_fd_sc_hd__and2_2 _1641_ (.A(_0193_),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__nand2_4 _1642_ (.A(_0192_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _1643_ (.A(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _1644_ (.A(_0021_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__a31o_1 _1645_ (.A1(_0015_),
    .A2(_0994_),
    .A3(_0196_),
    .B1(_0198_),
    .X(net703));
 sky130_fd_sc_hd__o22ai_2 _1646_ (.A1(net314),
    .A2(_1060_),
    .B1(net276),
    .B2(_1061_),
    .Y(_0199_));
 sky130_fd_sc_hd__o22ai_4 _1647_ (.A1(net254),
    .A2(_0995_),
    .B1(net351),
    .B2(_1036_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_4 _1648_ (.A(_0199_),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__and2_1 _1649_ (.A(_0201_),
    .B(_1029_),
    .X(_0202_));
 sky130_fd_sc_hd__buf_1 _1650_ (.A(_0202_),
    .X(net412));
 sky130_fd_sc_hd__nand2_1 _1651_ (.A(_0124_),
    .B(_1136_),
    .Y(_0203_));
 sky130_fd_sc_hd__nand3_1 _1652_ (.A(_0196_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _1653_ (.A(_1096_),
    .B(net203),
    .Y(_0205_));
 sky130_fd_sc_hd__nand2_1 _1654_ (.A(_0984_),
    .B(net123),
    .Y(_0206_));
 sky130_fd_sc_hd__and2_2 _1655_ (.A(_0205_),
    .B(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _1656_ (.A(_1143_),
    .B(net39),
    .Y(_0208_));
 sky130_fd_sc_hd__nand2_1 _1657_ (.A(_1145_),
    .B(net102),
    .Y(_0209_));
 sky130_fd_sc_hd__a21o_2 _1658_ (.A1(_0208_),
    .A2(_0209_),
    .B1(_1108_),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_4 _1659_ (.A(_0207_),
    .B(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _1660_ (.A(_0211_),
    .B(_0035_),
    .Y(_0212_));
 sky130_fd_sc_hd__nand2_1 _1661_ (.A(_0204_),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__nand2_1 _1662_ (.A(_0213_),
    .B(_0034_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand2_1 _1663_ (.A(_0203_),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__nand2_1 _1664_ (.A(_0215_),
    .B(_1161_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2_1 _1665_ (.A(_0211_),
    .B(_1139_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_2 _1666_ (.A(_0216_),
    .B(_0217_),
    .Y(net704));
 sky130_fd_sc_hd__nand3_1 _1667_ (.A(_0207_),
    .B(_0210_),
    .C(_1002_),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _1668_ (.A(_0160_),
    .Y(_0219_));
 sky130_fd_sc_hd__nand2_1 _1669_ (.A(_0219_),
    .B(_0993_),
    .Y(_0220_));
 sky130_fd_sc_hd__nand2_1 _1670_ (.A(_0218_),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _1671_ (.A(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _1672_ (.A(_0196_),
    .B(_1022_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand2_1 _1673_ (.A(_0223_),
    .B(_0094_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand3_1 _1674_ (.A(_0222_),
    .B(_0224_),
    .C(_1026_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand2_1 _1675_ (.A(_1143_),
    .B(net149),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _1676_ (.A(_1145_),
    .B(net212),
    .Y(_0227_));
 sky130_fd_sc_hd__nand2_1 _1677_ (.A(_0226_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_1 _1678_ (.A(_0228_),
    .B(_1108_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand2_1 _1679_ (.A(_0017_),
    .B(net48),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _1680_ (.A(_0016_),
    .B(net110),
    .Y(_0231_));
 sky130_fd_sc_hd__nand3_4 _1681_ (.A(_0229_),
    .B(_0230_),
    .C(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _1682_ (.A(_0232_),
    .B(_1002_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _1683_ (.A(_0225_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _1684_ (.A(_0234_),
    .B(_1161_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _1685_ (.A(_0160_),
    .B(_1139_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_2 _1686_ (.A(_0235_),
    .B(_0236_),
    .Y(net705));
 sky130_fd_sc_hd__nand2_1 _1687_ (.A(_1143_),
    .B(net148),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_1 _1688_ (.A(_1145_),
    .B(net211),
    .Y(_0238_));
 sky130_fd_sc_hd__a21o_1 _1689_ (.A1(_0237_),
    .A2(_0238_),
    .B1(_0983_),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _1690_ (.A(_1103_),
    .B(net47),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _1691_ (.A(_1105_),
    .B(net109),
    .Y(_0241_));
 sky130_fd_sc_hd__nand2_1 _1692_ (.A(_0240_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2_1 _1693_ (.A(_0242_),
    .B(_1114_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_4 _1694_ (.A(_0239_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__nand2_1 _1695_ (.A(_0244_),
    .B(_0991_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand2_1 _1696_ (.A(_0232_),
    .B(_1101_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand3_1 _1697_ (.A(_0245_),
    .B(_0246_),
    .C(_0094_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_1 _1698_ (.A(_1103_),
    .B(net150),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _1699_ (.A(_1105_),
    .B(net213),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(_0248_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _1701_ (.A(_0250_),
    .B(_1109_),
    .Y(_0251_));
 sky130_fd_sc_hd__nand2_1 _1702_ (.A(_0016_),
    .B(net113),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2_1 _1703_ (.A(_0017_),
    .B(net49),
    .Y(_0253_));
 sky130_fd_sc_hd__nand3_4 _1704_ (.A(_0251_),
    .B(_0252_),
    .C(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _1705_ (.A(_0254_),
    .B(_0991_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand2_1 _1706_ (.A(_1120_),
    .B(net152),
    .Y(_0256_));
 sky130_fd_sc_hd__nand2_1 _1707_ (.A(_1122_),
    .B(net214),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_1 _1708_ (.A(_0256_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__nand2_1 _1709_ (.A(_0258_),
    .B(_1109_),
    .Y(_0259_));
 sky130_fd_sc_hd__nand2_1 _1710_ (.A(_1103_),
    .B(net50),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _1711_ (.A(_1105_),
    .B(net114),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_1 _1712_ (.A(_0260_),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__nand2_1 _1713_ (.A(_0262_),
    .B(_1114_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_4 _1714_ (.A(_0259_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__nand2_1 _1715_ (.A(_0264_),
    .B(_1101_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand3_1 _1716_ (.A(_0255_),
    .B(_0265_),
    .C(_1134_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_2 _1717_ (.A(_0247_),
    .B(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__nand2_1 _1718_ (.A(_0267_),
    .B(_0125_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2_1 _1719_ (.A(_1143_),
    .B(net143),
    .Y(_0269_));
 sky130_fd_sc_hd__nand2_1 _1720_ (.A(_1145_),
    .B(net205),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _1721_ (.A(_0269_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__nand2_1 _1722_ (.A(_0271_),
    .B(_1108_),
    .Y(_0272_));
 sky130_fd_sc_hd__nand2_1 _1723_ (.A(_1143_),
    .B(net41),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _1724_ (.A(_1145_),
    .B(net104),
    .Y(_0274_));
 sky130_fd_sc_hd__nand2_1 _1725_ (.A(_0273_),
    .B(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand2_2 _1726_ (.A(_0275_),
    .B(_0983_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2_4 _1727_ (.A(_0272_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__nand2_1 _1728_ (.A(_0277_),
    .B(_0988_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_1 _1729_ (.A(_0161_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand2_1 _1730_ (.A(_0279_),
    .B(_0034_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_1 _1731_ (.A(_0211_),
    .B(_1136_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand3_1 _1732_ (.A(_0280_),
    .B(_1026_),
    .C(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand3_1 _1733_ (.A(_0268_),
    .B(_0282_),
    .C(_1188_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _1734_ (.A(_0277_),
    .B(_1139_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand2_1 _1735_ (.A(_0283_),
    .B(_0284_),
    .Y(net706));
 sky130_fd_sc_hd__a22oi_4 _1736_ (.A1(_1089_),
    .A2(net105),
    .B1(net42),
    .B2(_1092_),
    .Y(_0285_));
 sky130_fd_sc_hd__a22oi_2 _1737_ (.A1(_1094_),
    .A2(net144),
    .B1(_1097_),
    .B2(net207),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_4 _1738_ (.A(_0285_),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand2_1 _1739_ (.A(_0287_),
    .B(_0035_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _1740_ (.A(_0277_),
    .B(_0991_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _1741_ (.A(_0288_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _1742_ (.A(_0290_),
    .B(_0034_),
    .Y(_0291_));
 sky130_fd_sc_hd__nand2_1 _1743_ (.A(_0160_),
    .B(_1136_),
    .Y(_0292_));
 sky130_fd_sc_hd__nand2_1 _1744_ (.A(_0291_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _1745_ (.A(_0293_),
    .B(_1161_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _1746_ (.A(_0287_),
    .B(_1139_),
    .Y(_0295_));
 sky130_fd_sc_hd__nand2_2 _1747_ (.A(_0294_),
    .B(_0295_),
    .Y(net708));
 sky130_fd_sc_hd__a22oi_4 _1748_ (.A1(_1089_),
    .A2(net106),
    .B1(net43),
    .B2(_1092_),
    .Y(_0296_));
 sky130_fd_sc_hd__a22oi_2 _1749_ (.A1(_1094_),
    .A2(net145),
    .B1(_1097_),
    .B2(net208),
    .Y(_0297_));
 sky130_fd_sc_hd__nand2_4 _1750_ (.A(_0296_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__clkinv_4 _1751_ (.A(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _1752_ (.A(_0287_),
    .B(_1009_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _1753_ (.A(_0298_),
    .B(_1102_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand3_1 _1754_ (.A(_0300_),
    .B(_0301_),
    .C(_0034_),
    .Y(_0302_));
 sky130_fd_sc_hd__or2_1 _1755_ (.A(_1134_),
    .B(_0279_),
    .X(_0303_));
 sky130_fd_sc_hd__nand3_2 _1756_ (.A(_0302_),
    .B(_0303_),
    .C(_1160_),
    .Y(_0304_));
 sky130_fd_sc_hd__o21ai_2 _1757_ (.A1(_0021_),
    .A2(_0299_),
    .B1(_0304_),
    .Y(net709));
 sky130_fd_sc_hd__nand2_1 _1758_ (.A(_1120_),
    .B(net146),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _1759_ (.A(_1122_),
    .B(net209),
    .Y(_0306_));
 sky130_fd_sc_hd__nand2_1 _1760_ (.A(_0305_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__nand2_1 _1761_ (.A(_0307_),
    .B(_1109_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand2_1 _1762_ (.A(_1089_),
    .B(net107),
    .Y(_0309_));
 sky130_fd_sc_hd__nand2_1 _1763_ (.A(_1092_),
    .B(net44),
    .Y(_0310_));
 sky130_fd_sc_hd__nand3_4 _1764_ (.A(_0308_),
    .B(_0309_),
    .C(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _1765_ (.A(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__nand3_1 _1766_ (.A(_0288_),
    .B(_0094_),
    .C(_0289_),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _1767_ (.A(_0298_),
    .B(_1009_),
    .Y(_0314_));
 sky130_fd_sc_hd__nand2_1 _1768_ (.A(_0311_),
    .B(_1102_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand3_1 _1769_ (.A(_0314_),
    .B(_0034_),
    .C(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand3_2 _1770_ (.A(_0313_),
    .B(_0316_),
    .C(_1160_),
    .Y(_0317_));
 sky130_fd_sc_hd__o21ai_2 _1771_ (.A1(_0021_),
    .A2(_0312_),
    .B1(_0317_),
    .Y(net710));
 sky130_fd_sc_hd__nand2_1 _1772_ (.A(_0311_),
    .B(_1009_),
    .Y(_0318_));
 sky130_fd_sc_hd__nand2_1 _1773_ (.A(_1120_),
    .B(net147),
    .Y(_0319_));
 sky130_fd_sc_hd__nand2_1 _1774_ (.A(_1122_),
    .B(net210),
    .Y(_0320_));
 sky130_fd_sc_hd__nand2_1 _1775_ (.A(_0319_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_1 _1776_ (.A(_0321_),
    .B(_1109_),
    .Y(_0322_));
 sky130_fd_sc_hd__nand2_1 _1777_ (.A(_1120_),
    .B(net46),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2_1 _1778_ (.A(_1122_),
    .B(net108),
    .Y(_0324_));
 sky130_fd_sc_hd__nand2_1 _1779_ (.A(_0323_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2_1 _1780_ (.A(_0325_),
    .B(_1114_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_4 _1781_ (.A(_0322_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_1 _1782_ (.A(_0327_),
    .B(_0035_),
    .Y(_0328_));
 sky130_fd_sc_hd__nand2_1 _1783_ (.A(_0318_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_1 _1784_ (.A(_0329_),
    .B(_0034_),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _1785_ (.A(_0298_),
    .B(_1136_),
    .Y(_0331_));
 sky130_fd_sc_hd__nand3_1 _1786_ (.A(_0330_),
    .B(_0331_),
    .C(_1026_),
    .Y(_0332_));
 sky130_fd_sc_hd__nand2_1 _1787_ (.A(_1103_),
    .B(net155),
    .Y(_0333_));
 sky130_fd_sc_hd__nand2_1 _1788_ (.A(_1105_),
    .B(net218),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2_1 _1789_ (.A(_0333_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _1790_ (.A(_0335_),
    .B(_1109_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_1 _1791_ (.A(_1103_),
    .B(net53),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _1792_ (.A(_1105_),
    .B(net117),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _1793_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _1794_ (.A(_0339_),
    .B(_1114_),
    .Y(_0340_));
 sky130_fd_sc_hd__nand2_4 _1795_ (.A(_0336_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand2_1 _1796_ (.A(_0341_),
    .B(_0991_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _1797_ (.A(_1120_),
    .B(net156),
    .Y(_0343_));
 sky130_fd_sc_hd__nand2_1 _1798_ (.A(_1122_),
    .B(net219),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _1799_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_1 _1800_ (.A(_0345_),
    .B(_1109_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand2_1 _1801_ (.A(_1120_),
    .B(net54),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _1802_ (.A(_1122_),
    .B(net118),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _1803_ (.A(_0347_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _1804_ (.A(_0349_),
    .B(_1114_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_4 _1805_ (.A(_0346_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _1806_ (.A(_0351_),
    .B(_0035_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _1807_ (.A(_0342_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _1808_ (.A(_0353_),
    .B(_1134_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _1809_ (.A(_1103_),
    .B(net154),
    .Y(_0355_));
 sky130_fd_sc_hd__nand2_1 _1810_ (.A(_1105_),
    .B(net216),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _1811_ (.A(_0355_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand2_1 _1812_ (.A(_0357_),
    .B(_1109_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _1813_ (.A(_1103_),
    .B(net52),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_1 _1814_ (.A(_1145_),
    .B(net116),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _1815_ (.A(_0359_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _1816_ (.A(_0361_),
    .B(_1114_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2_4 _1817_ (.A(_0358_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__nand2_1 _1818_ (.A(_0363_),
    .B(_1136_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand3_1 _1819_ (.A(_0354_),
    .B(_0125_),
    .C(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__nand3_1 _1820_ (.A(_0332_),
    .B(_1188_),
    .C(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _1821_ (.A(_0327_),
    .B(_1139_),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_2 _1822_ (.A(_0366_),
    .B(_0367_),
    .Y(net711));
 sky130_fd_sc_hd__inv_2 _1823_ (.A(_0244_),
    .Y(_0368_));
 sky130_fd_sc_hd__nor2_1 _1824_ (.A(_0021_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__a31o_1 _1825_ (.A1(_0015_),
    .A2(_0994_),
    .A3(_0244_),
    .B1(_0369_),
    .X(net712));
 sky130_fd_sc_hd__inv_2 _1826_ (.A(net220),
    .Y(_0370_));
 sky130_fd_sc_hd__inv_2 _1827_ (.A(net157),
    .Y(_0371_));
 sky130_fd_sc_hd__a22oi_4 _1828_ (.A1(_0016_),
    .A2(net119),
    .B1(net55),
    .B2(_0017_),
    .Y(_0372_));
 sky130_fd_sc_hd__o221ai_4 _1829_ (.A1(_0370_),
    .A2(_0122_),
    .B1(_0371_),
    .B2(_0985_),
    .C1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_2 _1830_ (.A(_0373_),
    .B(_1009_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand3_1 _1831_ (.A(_0245_),
    .B(_0246_),
    .C(_1134_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _1832_ (.A(_0328_),
    .B(_1020_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _1833_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2_4 _1834_ (.A(_0374_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__nand2_1 _1835_ (.A(_0378_),
    .B(_1161_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _1836_ (.A(_0232_),
    .B(_1139_),
    .Y(_0380_));
 sky130_fd_sc_hd__nand2_1 _1837_ (.A(_0379_),
    .B(_0380_),
    .Y(net713));
 sky130_fd_sc_hd__inv_2 _1838_ (.A(_0254_),
    .Y(_0381_));
 sky130_fd_sc_hd__nand2_1 _1839_ (.A(_0254_),
    .B(_1101_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_2 _1840_ (.A(_0233_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand2_1 _1841_ (.A(_0383_),
    .B(_1134_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_1 _1842_ (.A(_0244_),
    .B(_1136_),
    .Y(_0385_));
 sky130_fd_sc_hd__a21o_1 _1843_ (.A1(_0384_),
    .A2(_0385_),
    .B1(_1084_),
    .X(_0386_));
 sky130_fd_sc_hd__o21ai_2 _1844_ (.A1(_0021_),
    .A2(_0381_),
    .B1(_0386_),
    .Y(net714));
 sky130_fd_sc_hd__o22ai_2 _1845_ (.A1(net315),
    .A2(_1060_),
    .B1(net278),
    .B2(_1061_),
    .Y(_0387_));
 sky130_fd_sc_hd__o22ai_4 _1846_ (.A1(net255),
    .A2(_0995_),
    .B1(net352),
    .B2(_1036_),
    .Y(_0388_));
 sky130_fd_sc_hd__nor2_4 _1847_ (.A(_0387_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__and2_1 _1848_ (.A(_0389_),
    .B(_1029_),
    .X(_0390_));
 sky130_fd_sc_hd__buf_1 _1849_ (.A(_0390_),
    .X(net414));
 sky130_fd_sc_hd__inv_2 _1850_ (.A(_0264_),
    .Y(_0391_));
 sky130_fd_sc_hd__o22ai_4 _1851_ (.A1(_1082_),
    .A2(_0391_),
    .B1(_1084_),
    .B2(_0267_),
    .Y(net715));
 sky130_fd_sc_hd__nand2_1 _1852_ (.A(_1103_),
    .B(net153),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _1853_ (.A(_1105_),
    .B(net215),
    .Y(_0393_));
 sky130_fd_sc_hd__nand2_1 _1854_ (.A(_0392_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__nand2_1 _1855_ (.A(_0394_),
    .B(_1109_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_1 _1856_ (.A(_0017_),
    .B(net51),
    .Y(_0396_));
 sky130_fd_sc_hd__nand2_1 _1857_ (.A(_0016_),
    .B(net115),
    .Y(_0397_));
 sky130_fd_sc_hd__nand3_4 _1858_ (.A(_0395_),
    .B(_0396_),
    .C(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_1 _1859_ (.A(_0398_),
    .B(_0035_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _1860_ (.A(_0264_),
    .B(_0991_),
    .Y(_0400_));
 sky130_fd_sc_hd__nand3_2 _1861_ (.A(_0399_),
    .B(_0034_),
    .C(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__a22o_1 _1862_ (.A1(_1081_),
    .A2(_0398_),
    .B1(_0401_),
    .B2(_1188_),
    .X(net716));
 sky130_fd_sc_hd__nand3_1 _1863_ (.A(_0255_),
    .B(_0265_),
    .C(_0094_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2_1 _1864_ (.A(_0398_),
    .B(_0991_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _1865_ (.A(_0363_),
    .B(_0035_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand3_1 _1866_ (.A(_0403_),
    .B(_0404_),
    .C(_1134_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand2_1 _1867_ (.A(_0402_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _1868_ (.A(_0406_),
    .B(_1026_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _1869_ (.A(_1143_),
    .B(net160),
    .Y(_0408_));
 sky130_fd_sc_hd__nand2_1 _1870_ (.A(_1145_),
    .B(net223),
    .Y(_0409_));
 sky130_fd_sc_hd__a21o_1 _1871_ (.A1(_0408_),
    .A2(_0409_),
    .B1(_0983_),
    .X(_0410_));
 sky130_fd_sc_hd__nand2_1 _1872_ (.A(_1143_),
    .B(net59),
    .Y(_0411_));
 sky130_fd_sc_hd__nand2_1 _1873_ (.A(_0982_),
    .B(net122),
    .Y(_0412_));
 sky130_fd_sc_hd__a21o_1 _1874_ (.A1(_0411_),
    .A2(_0412_),
    .B1(_1108_),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_4 _1875_ (.A(_0410_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__nand2_1 _1876_ (.A(_0414_),
    .B(_0996_),
    .Y(_0415_));
 sky130_fd_sc_hd__nand2_1 _1877_ (.A(_1095_),
    .B(net163),
    .Y(_0416_));
 sky130_fd_sc_hd__nand2_1 _1878_ (.A(_0982_),
    .B(net225),
    .Y(_0417_));
 sky130_fd_sc_hd__nand2_1 _1879_ (.A(_0416_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _1880_ (.A(_0418_),
    .B(_1108_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _1881_ (.A(_1088_),
    .B(net125),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _1882_ (.A(_1091_),
    .B(net61),
    .Y(_0421_));
 sky130_fd_sc_hd__nand3_4 _1883_ (.A(_0419_),
    .B(_0420_),
    .C(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand2_1 _1884_ (.A(_0422_),
    .B(_0993_),
    .Y(_0423_));
 sky130_fd_sc_hd__nand2_1 _1885_ (.A(_0415_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_2 _1886_ (.A(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a22oi_4 _1887_ (.A1(_1089_),
    .A2(net124),
    .B1(net60),
    .B2(_1092_),
    .Y(_0426_));
 sky130_fd_sc_hd__a22oi_2 _1888_ (.A1(_1094_),
    .A2(net161),
    .B1(_1097_),
    .B2(net224),
    .Y(_0427_));
 sky130_fd_sc_hd__nand2_4 _1889_ (.A(_0426_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__nand2_1 _1890_ (.A(_0428_),
    .B(_1009_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand3_1 _1891_ (.A(_0425_),
    .B(_0125_),
    .C(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand3_1 _1892_ (.A(_0407_),
    .B(_0430_),
    .C(_1188_),
    .Y(_0431_));
 sky130_fd_sc_hd__nand2_1 _1893_ (.A(_0363_),
    .B(_1139_),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _1894_ (.A(_0431_),
    .B(_0432_),
    .Y(net717));
 sky130_fd_sc_hd__nand3_1 _1895_ (.A(_0399_),
    .B(_0094_),
    .C(_0400_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2_1 _1896_ (.A(_0363_),
    .B(_0991_),
    .Y(_0434_));
 sky130_fd_sc_hd__nand2_1 _1897_ (.A(_0341_),
    .B(_1101_),
    .Y(_0435_));
 sky130_fd_sc_hd__nand3_1 _1898_ (.A(_0434_),
    .B(_0435_),
    .C(_1134_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand2_1 _1899_ (.A(_0433_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _1900_ (.A(_0437_),
    .B(_1026_),
    .Y(_0438_));
 sky130_fd_sc_hd__nand2_1 _1901_ (.A(_0422_),
    .B(_1002_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(_1103_),
    .B(net164),
    .Y(_0440_));
 sky130_fd_sc_hd__nand2_1 _1903_ (.A(_1105_),
    .B(net226),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_1 _1904_ (.A(_0440_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _1905_ (.A(_0442_),
    .B(_1109_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _1906_ (.A(_1103_),
    .B(net62),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _1907_ (.A(_1105_),
    .B(net126),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _1908_ (.A(_0444_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_1 _1909_ (.A(_0446_),
    .B(_1114_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_4 _1910_ (.A(_0443_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _1911_ (.A(_0448_),
    .B(_1101_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _1912_ (.A(_0439_),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_1 _1913_ (.A(_0450_),
    .B(_1134_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_2 _1914_ (.A(_0428_),
    .B(_0996_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand3_1 _1915_ (.A(_0451_),
    .B(_0125_),
    .C(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand3_1 _1916_ (.A(_0438_),
    .B(_0453_),
    .C(_1188_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand2_1 _1917_ (.A(_0341_),
    .B(_1081_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_2 _1918_ (.A(_0454_),
    .B(_0455_),
    .Y(net719));
 sky130_fd_sc_hd__nand2_1 _1919_ (.A(_1120_),
    .B(net165),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _1920_ (.A(_1122_),
    .B(net227),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _1921_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand2_1 _1922_ (.A(_0458_),
    .B(_1109_),
    .Y(_0459_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(_1089_),
    .B(net127),
    .Y(_0460_));
 sky130_fd_sc_hd__nand2_1 _1924_ (.A(_1092_),
    .B(net63),
    .Y(_0461_));
 sky130_fd_sc_hd__nand3_4 _1925_ (.A(_0459_),
    .B(_0460_),
    .C(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _1926_ (.A(_0462_),
    .B(_0035_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _1927_ (.A(_0448_),
    .B(_0991_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand2_1 _1928_ (.A(_0463_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_1 _1929_ (.A(_0465_),
    .B(_1134_),
    .Y(_0466_));
 sky130_fd_sc_hd__nand2_1 _1930_ (.A(_0422_),
    .B(_1136_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand3_1 _1931_ (.A(_0466_),
    .B(_0125_),
    .C(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand3_1 _1932_ (.A(_0354_),
    .B(_1026_),
    .C(_0364_),
    .Y(_0469_));
 sky130_fd_sc_hd__nand3_1 _1933_ (.A(_0468_),
    .B(_0469_),
    .C(_1188_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _1934_ (.A(_0351_),
    .B(_1081_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_2 _1935_ (.A(_0470_),
    .B(_0471_),
    .Y(net720));
 sky130_fd_sc_hd__inv_2 _1936_ (.A(_0373_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand3_1 _1937_ (.A(_0373_),
    .B(_0015_),
    .C(_0994_),
    .Y(_0473_));
 sky130_fd_sc_hd__o21ai_2 _1938_ (.A1(_0021_),
    .A2(_0472_),
    .B1(_0473_),
    .Y(net721));
 sky130_fd_sc_hd__a22oi_4 _1939_ (.A1(_1089_),
    .A2(net120),
    .B1(net57),
    .B2(_1092_),
    .Y(_0474_));
 sky130_fd_sc_hd__a22oi_2 _1940_ (.A1(_1094_),
    .A2(net158),
    .B1(_1097_),
    .B2(net221),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_4 _1941_ (.A(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _1942_ (.A(_0476_),
    .B(_1102_),
    .Y(_0477_));
 sky130_fd_sc_hd__nand2_2 _1943_ (.A(_0374_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_1 _1944_ (.A(_0478_),
    .B(_1161_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2_1 _1945_ (.A(_0476_),
    .B(_1081_),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_1 _1946_ (.A(_0479_),
    .B(_0480_),
    .Y(net722));
 sky130_fd_sc_hd__a22oi_4 _1947_ (.A1(_1089_),
    .A2(net121),
    .B1(net58),
    .B2(_1092_),
    .Y(_0481_));
 sky130_fd_sc_hd__a22oi_2 _1948_ (.A1(_1094_),
    .A2(net159),
    .B1(_1097_),
    .B2(net222),
    .Y(_0482_));
 sky130_fd_sc_hd__nand2_2 _1949_ (.A(_0481_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__inv_2 _1950_ (.A(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__buf_8 _1951_ (.A(_0981_),
    .X(_0485_));
 sky130_fd_sc_hd__nand2_1 _1952_ (.A(_0476_),
    .B(_1009_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand2_1 _1953_ (.A(_0483_),
    .B(_0035_),
    .Y(_0487_));
 sky130_fd_sc_hd__nand2_1 _1954_ (.A(_0486_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _1955_ (.A(_0488_),
    .B(_0994_),
    .Y(_0489_));
 sky130_fd_sc_hd__o22ai_2 _1956_ (.A1(_1082_),
    .A2(_0484_),
    .B1(_0485_),
    .B2(_0489_),
    .Y(net723));
 sky130_fd_sc_hd__inv_2 _1957_ (.A(_0414_),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _1958_ (.A(_0483_),
    .B(_1009_),
    .Y(_0491_));
 sky130_fd_sc_hd__o211ai_1 _1959_ (.A1(_1142_),
    .A2(_0490_),
    .B1(_0034_),
    .C1(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__nand2_1 _1960_ (.A(_0492_),
    .B(_1161_),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_2 _1961_ (.A1(_0021_),
    .A2(_0490_),
    .B1(_0493_),
    .Y(net724));
 sky130_fd_sc_hd__clkinv_4 _1962_ (.A(_0428_),
    .Y(_0494_));
 sky130_fd_sc_hd__nand3_1 _1963_ (.A(_0486_),
    .B(_0487_),
    .C(_0094_),
    .Y(_0495_));
 sky130_fd_sc_hd__nand2_1 _1964_ (.A(_0428_),
    .B(_1102_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _1965_ (.A(_0414_),
    .B(_1009_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand3_1 _1966_ (.A(_0496_),
    .B(_0034_),
    .C(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand3_1 _1967_ (.A(_0495_),
    .B(_0498_),
    .C(_1160_),
    .Y(_0499_));
 sky130_fd_sc_hd__o21ai_2 _1968_ (.A1(_0021_),
    .A2(_0494_),
    .B1(_0499_),
    .Y(net725));
 sky130_fd_sc_hd__o22ai_2 _1969_ (.A1(net316),
    .A2(_1060_),
    .B1(net279),
    .B2(_1061_),
    .Y(_0500_));
 sky130_fd_sc_hd__o22ai_4 _1970_ (.A1(net256),
    .A2(_0995_),
    .B1(net353),
    .B2(_1036_),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2_4 _1971_ (.A(_0500_),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__and2_1 _1972_ (.A(_0502_),
    .B(_1029_),
    .X(_0503_));
 sky130_fd_sc_hd__buf_1 _1973_ (.A(_0503_),
    .X(net415));
 sky130_fd_sc_hd__buf_6 _1974_ (.A(_0981_),
    .X(_0504_));
 sky130_fd_sc_hd__a2bb2o_1 _1975_ (.A1_N(_0504_),
    .A2_N(_0423_),
    .B1(_1081_),
    .B2(_0422_),
    .X(net726));
 sky130_fd_sc_hd__nand2_1 _1976_ (.A(_1103_),
    .B(net171),
    .Y(_0505_));
 sky130_fd_sc_hd__nand2_1 _1977_ (.A(_1105_),
    .B(net7),
    .Y(_0506_));
 sky130_fd_sc_hd__a21o_1 _1978_ (.A1(_0505_),
    .A2(_0506_),
    .B1(_1114_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _1979_ (.A(_1120_),
    .B(net70),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _1980_ (.A(_1122_),
    .B(net133),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_1 _1981_ (.A(_0508_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _1982_ (.A(_0510_),
    .B(_1114_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_4 _1983_ (.A(_0507_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand2_1 _1984_ (.A(_0512_),
    .B(_0991_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _1985_ (.A(_1143_),
    .B(net172),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_1 _1986_ (.A(_1145_),
    .B(net8),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _1987_ (.A(_0514_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _1988_ (.A(_0516_),
    .B(_1108_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_1 _1989_ (.A(_0016_),
    .B(net135),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _1990_ (.A(_0017_),
    .B(net71),
    .Y(_0519_));
 sky130_fd_sc_hd__nand3_4 _1991_ (.A(_0517_),
    .B(_0518_),
    .C(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _1992_ (.A(_0520_),
    .B(_0035_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _1993_ (.A(_0513_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _1994_ (.A(_0522_),
    .B(_1134_),
    .Y(_0523_));
 sky130_fd_sc_hd__a22oi_4 _1995_ (.A1(_1089_),
    .A2(net132),
    .B1(net69),
    .B2(_1092_),
    .Y(_0524_));
 sky130_fd_sc_hd__a22oi_2 _1996_ (.A1(_1094_),
    .A2(net170),
    .B1(_1097_),
    .B2(net6),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_4 _1997_ (.A(_0524_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_2 _1998_ (.A(_0526_),
    .B(_1136_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand3_1 _1999_ (.A(_0523_),
    .B(_0527_),
    .C(_0125_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand3_1 _2000_ (.A(_0451_),
    .B(_1026_),
    .C(_0452_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand3_1 _2001_ (.A(_0528_),
    .B(_0529_),
    .C(_1188_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _2002_ (.A(_0448_),
    .B(_1081_),
    .Y(_0531_));
 sky130_fd_sc_hd__nand2_2 _2003_ (.A(_0530_),
    .B(_0531_),
    .Y(net727));
 sky130_fd_sc_hd__nand3_1 _2004_ (.A(_0466_),
    .B(_1026_),
    .C(_0467_),
    .Y(_0532_));
 sky130_fd_sc_hd__or3_1 _2005_ (.A(_1101_),
    .B(_0989_),
    .C(_0520_),
    .X(_0533_));
 sky130_fd_sc_hd__nand3_1 _2006_ (.A(_0532_),
    .B(_0533_),
    .C(_1188_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _2007_ (.A(_0462_),
    .B(_1081_),
    .Y(_0535_));
 sky130_fd_sc_hd__nand2_2 _2008_ (.A(_0534_),
    .B(_0535_),
    .Y(net728));
 sky130_fd_sc_hd__nand2_1 _2009_ (.A(_1096_),
    .B(net2),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _2010_ (.A(_0984_),
    .B(net166),
    .Y(_0537_));
 sky130_fd_sc_hd__and2_1 _2011_ (.A(_0536_),
    .B(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__nand2_1 _2012_ (.A(_0017_),
    .B(net64),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _2013_ (.A(_0016_),
    .B(net128),
    .Y(_0540_));
 sky130_fd_sc_hd__and2_2 _2014_ (.A(_0539_),
    .B(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__nand2_2 _2015_ (.A(_0538_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _2016_ (.A(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__nor2_1 _2017_ (.A(_1086_),
    .B(_0543_),
    .Y(net503));
 sky130_fd_sc_hd__nand2_1 _2018_ (.A(_1091_),
    .B(net65),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _2019_ (.A(_1088_),
    .B(net129),
    .Y(_0545_));
 sky130_fd_sc_hd__and2_2 _2020_ (.A(_0544_),
    .B(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__nand2_1 _2021_ (.A(_1096_),
    .B(net3),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _2022_ (.A(_0984_),
    .B(net167),
    .Y(_0548_));
 sky130_fd_sc_hd__and2_1 _2023_ (.A(_0547_),
    .B(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_4 _2024_ (.A(_0546_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__nand2_1 _2025_ (.A(_0550_),
    .B(_0035_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _2026_ (.A(_0542_),
    .B(_0991_),
    .Y(_0552_));
 sky130_fd_sc_hd__nand3_1 _2027_ (.A(_0551_),
    .B(_0552_),
    .C(_1134_),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_1 _2028_ (.A(_0463_),
    .B(_1020_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _2029_ (.A(_0553_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_2 _2030_ (.A(net10),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_2 _2031_ (.A(net175),
    .Y(_0557_));
 sky130_fd_sc_hd__a22oi_4 _2032_ (.A1(_1089_),
    .A2(net137),
    .B1(net73),
    .B2(_1092_),
    .Y(_0558_));
 sky130_fd_sc_hd__o221ai_4 _2033_ (.A1(_0556_),
    .A2(_0122_),
    .B1(_0557_),
    .B2(_0985_),
    .C1(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _2034_ (.A(_0559_),
    .B(_1009_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_2 _2035_ (.A(_0555_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _2036_ (.A(_0561_),
    .B(_1161_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _2037_ (.A(_0550_),
    .B(_1081_),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2_1 _2038_ (.A(_0562_),
    .B(_0563_),
    .Y(net504));
 sky130_fd_sc_hd__nand2_1 _2039_ (.A(_0017_),
    .B(net66),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _2040_ (.A(_0016_),
    .B(net130),
    .Y(_0565_));
 sky130_fd_sc_hd__and2_2 _2041_ (.A(_0564_),
    .B(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__nand2_1 _2042_ (.A(_1096_),
    .B(net4),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _2043_ (.A(_0984_),
    .B(net168),
    .Y(_0568_));
 sky130_fd_sc_hd__and2_1 _2044_ (.A(_0567_),
    .B(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_4 _2045_ (.A(_0566_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_1 _2047_ (.A(_0550_),
    .B(_1009_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2_1 _2048_ (.A(_0570_),
    .B(_0035_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_1 _2049_ (.A(_0572_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand3_2 _2050_ (.A(_0574_),
    .B(_1102_),
    .C(_0989_),
    .Y(_0575_));
 sky130_fd_sc_hd__o22ai_2 _2051_ (.A1(_1082_),
    .A2(_0571_),
    .B1(_0485_),
    .B2(_0575_),
    .Y(net505));
 sky130_fd_sc_hd__nand2_1 _2052_ (.A(_0570_),
    .B(_0991_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _2053_ (.A(_1096_),
    .B(net5),
    .Y(_0577_));
 sky130_fd_sc_hd__nand2_1 _2054_ (.A(_0984_),
    .B(net169),
    .Y(_0578_));
 sky130_fd_sc_hd__and2_1 _2055_ (.A(_0577_),
    .B(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__nand2_1 _2056_ (.A(_1091_),
    .B(net68),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_1 _2057_ (.A(_0016_),
    .B(net131),
    .Y(_0581_));
 sky130_fd_sc_hd__and2_2 _2058_ (.A(_0580_),
    .B(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_4 _2059_ (.A(_0579_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_1 _2060_ (.A(_0583_),
    .B(_0035_),
    .Y(_0584_));
 sky130_fd_sc_hd__nand3_1 _2061_ (.A(_0576_),
    .B(_0584_),
    .C(_1134_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_1 _2062_ (.A(_0551_),
    .B(_1020_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _2063_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__a22oi_4 _2064_ (.A1(_1089_),
    .A2(net139),
    .B1(net75),
    .B2(_1092_),
    .Y(_0588_));
 sky130_fd_sc_hd__a22oi_2 _2065_ (.A1(_1094_),
    .A2(net177),
    .B1(_1097_),
    .B2(net13),
    .Y(_0589_));
 sky130_fd_sc_hd__nand2_2 _2066_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _2067_ (.A(_0590_),
    .B(_1009_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _2068_ (.A(_0587_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _2069_ (.A(_0592_),
    .B(_1161_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _2070_ (.A(_0583_),
    .B(_1081_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_2 _2071_ (.A(_0593_),
    .B(_0594_),
    .Y(net506));
 sky130_fd_sc_hd__clkinv_4 _2072_ (.A(_0526_),
    .Y(_0595_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(_1086_),
    .B(_0595_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _2074_ (.A(_0512_),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_1 _2075_ (.A(_0021_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__a31o_1 _2076_ (.A1(_0015_),
    .A2(_0994_),
    .A3(_0512_),
    .B1(_0597_),
    .X(net508));
 sky130_fd_sc_hd__nand3_1 _2077_ (.A(_0523_),
    .B(_0527_),
    .C(_1026_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2_1 _2078_ (.A(_1096_),
    .B(net16),
    .Y(_0599_));
 sky130_fd_sc_hd__nand2_1 _2079_ (.A(_0984_),
    .B(net180),
    .Y(_0600_));
 sky130_fd_sc_hd__and2_1 _2080_ (.A(_0599_),
    .B(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__nand2_1 _2081_ (.A(_0017_),
    .B(net79),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _2082_ (.A(_0016_),
    .B(net142),
    .Y(_0603_));
 sky130_fd_sc_hd__and2_2 _2083_ (.A(_0602_),
    .B(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_2 _2084_ (.A(_0601_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__clkinv_4 _2085_ (.A(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _2086_ (.A(_0606_),
    .B(_0125_),
    .Y(_0607_));
 sky130_fd_sc_hd__nand3_2 _2087_ (.A(_0598_),
    .B(_1188_),
    .C(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _2088_ (.A(_0520_),
    .B(_1081_),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _2089_ (.A(_0608_),
    .B(_0609_),
    .Y(net509));
 sky130_fd_sc_hd__o22ai_2 _2090_ (.A1(net317),
    .A2(_1060_),
    .B1(net280),
    .B2(_1061_),
    .Y(_0610_));
 sky130_fd_sc_hd__o22ai_4 _2091_ (.A1(net257),
    .A2(_0995_),
    .B1(net355),
    .B2(_1036_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_4 _2092_ (.A(_0610_),
    .B(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__and2_1 _2093_ (.A(_0612_),
    .B(_0986_),
    .X(_0613_));
 sky130_fd_sc_hd__buf_1 _2094_ (.A(_0613_),
    .X(net416));
 sky130_fd_sc_hd__inv_2 _2095_ (.A(net174),
    .Y(_0614_));
 sky130_fd_sc_hd__inv_2 _2096_ (.A(net9),
    .Y(_0615_));
 sky130_fd_sc_hd__a22oi_4 _2097_ (.A1(_1089_),
    .A2(net136),
    .B1(net72),
    .B2(_1092_),
    .Y(_0616_));
 sky130_fd_sc_hd__o221ai_4 _2098_ (.A1(_0614_),
    .A2(_0985_),
    .B1(_0615_),
    .B2(_0122_),
    .C1(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand2_1 _2099_ (.A(_0617_),
    .B(_1102_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _2100_ (.A(_0520_),
    .B(_1009_),
    .Y(_0619_));
 sky130_fd_sc_hd__nand2_1 _2101_ (.A(_0618_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nand2_1 _2102_ (.A(_0620_),
    .B(_1161_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand2_1 _2103_ (.A(_0617_),
    .B(_1081_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_2 _2104_ (.A(_0621_),
    .B(_0622_),
    .Y(net510));
 sky130_fd_sc_hd__nand2_1 _2105_ (.A(_0617_),
    .B(_0125_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _2106_ (.A(_0559_),
    .B(_1102_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _2107_ (.A(_0623_),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _2108_ (.A(_0625_),
    .B(_1161_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _2109_ (.A(_0559_),
    .B(_1081_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_4 _2110_ (.A(_0626_),
    .B(_0627_),
    .Y(net511));
 sky130_fd_sc_hd__a22oi_2 _2111_ (.A1(_0984_),
    .A2(net176),
    .B1(_1096_),
    .B2(net11),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _2112_ (.A(_1095_),
    .B(net74),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _2113_ (.A(_0982_),
    .B(net138),
    .Y(_0630_));
 sky130_fd_sc_hd__a21o_1 _2114_ (.A1(_0629_),
    .A2(_0630_),
    .B1(_1108_),
    .X(_0631_));
 sky130_fd_sc_hd__nand2_4 _2115_ (.A(_0628_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand2_1 _2116_ (.A(_0632_),
    .B(_1102_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand2_1 _2117_ (.A(_0560_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _2118_ (.A(_0634_),
    .B(_1161_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2_1 _2119_ (.A(_0632_),
    .B(_1081_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_2 _2120_ (.A(_0635_),
    .B(_0636_),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _2121_ (.A(_0590_),
    .Y(_0637_));
 sky130_fd_sc_hd__nor2_1 _2122_ (.A(_1086_),
    .B(_0637_),
    .Y(net514));
 sky130_fd_sc_hd__a22oi_4 _2123_ (.A1(_1089_),
    .A2(net140),
    .B1(net76),
    .B2(_1092_),
    .Y(_0638_));
 sky130_fd_sc_hd__a22oi_2 _2124_ (.A1(_1094_),
    .A2(net178),
    .B1(_1097_),
    .B2(net14),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_2 _2125_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nand2_1 _2126_ (.A(_0640_),
    .B(_1102_),
    .Y(_0641_));
 sky130_fd_sc_hd__nand2_1 _2127_ (.A(_0591_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__a22o_2 _2128_ (.A1(_1081_),
    .A2(_0640_),
    .B1(_0642_),
    .B2(_1188_),
    .X(net515));
 sky130_fd_sc_hd__nand2_1 _2129_ (.A(_0017_),
    .B(net77),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _2130_ (.A(_0016_),
    .B(net141),
    .Y(_0644_));
 sky130_fd_sc_hd__and2_2 _2131_ (.A(_0643_),
    .B(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nand2_1 _2132_ (.A(_1096_),
    .B(net15),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _2133_ (.A(_0984_),
    .B(net179),
    .Y(_0647_));
 sky130_fd_sc_hd__and2_1 _2134_ (.A(_0646_),
    .B(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__nand2_2 _2135_ (.A(_0645_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__inv_2 _2136_ (.A(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _2137_ (.A(_1086_),
    .B(_0650_),
    .Y(net516));
 sky130_fd_sc_hd__nor2_1 _2138_ (.A(_1086_),
    .B(_0606_),
    .Y(net517));
 sky130_fd_sc_hd__o22ai_2 _2139_ (.A1(net318),
    .A2(_1060_),
    .B1(net281),
    .B2(_1061_),
    .Y(_0651_));
 sky130_fd_sc_hd__o22ai_4 _2140_ (.A1(net258),
    .A2(_0995_),
    .B1(net356),
    .B2(_1036_),
    .Y(_0652_));
 sky130_fd_sc_hd__nor2_4 _2141_ (.A(_0651_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__and2_1 _2142_ (.A(_0653_),
    .B(_0986_),
    .X(_0654_));
 sky130_fd_sc_hd__buf_1 _2143_ (.A(_0654_),
    .X(net417));
 sky130_fd_sc_hd__o22ai_2 _2144_ (.A1(net319),
    .A2(_1060_),
    .B1(net282),
    .B2(_1061_),
    .Y(_0655_));
 sky130_fd_sc_hd__o22ai_4 _2145_ (.A1(net259),
    .A2(_0995_),
    .B1(net357),
    .B2(_1025_),
    .Y(_0656_));
 sky130_fd_sc_hd__nor2_4 _2146_ (.A(_0655_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__and2_1 _2147_ (.A(_0657_),
    .B(_0986_),
    .X(_0658_));
 sky130_fd_sc_hd__buf_1 _2148_ (.A(_0658_),
    .X(net418));
 sky130_fd_sc_hd__o22ai_2 _2149_ (.A1(net320),
    .A2(_1060_),
    .B1(net283),
    .B2(_1061_),
    .Y(_0659_));
 sky130_fd_sc_hd__o22ai_4 _2150_ (.A1(net260),
    .A2(_0995_),
    .B1(net358),
    .B2(_1025_),
    .Y(_0660_));
 sky130_fd_sc_hd__nor2_4 _2151_ (.A(_0659_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__and2_1 _2152_ (.A(_0661_),
    .B(_0986_),
    .X(_0662_));
 sky130_fd_sc_hd__buf_1 _2153_ (.A(_0662_),
    .X(net419));
 sky130_fd_sc_hd__nand2_1 _2154_ (.A(_1142_),
    .B(net359),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _2155_ (.A(_1101_),
    .B(net261),
    .Y(_0664_));
 sky130_fd_sc_hd__o22ai_2 _2156_ (.A1(net322),
    .A2(_1060_),
    .B1(net284),
    .B2(_1061_),
    .Y(_0665_));
 sky130_fd_sc_hd__a31o_4 _2157_ (.A1(_1013_),
    .A2(_0663_),
    .A3(_0664_),
    .B1(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__nor2_1 _2158_ (.A(_0987_),
    .B(_0666_),
    .Y(net420));
 sky130_fd_sc_hd__nand2_1 _2159_ (.A(_1142_),
    .B(net360),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2_1 _2160_ (.A(_1101_),
    .B(net262),
    .Y(_0668_));
 sky130_fd_sc_hd__o22ai_2 _2161_ (.A1(net323),
    .A2(_1060_),
    .B1(net285),
    .B2(_1061_),
    .Y(_0669_));
 sky130_fd_sc_hd__a31o_4 _2162_ (.A1(_1013_),
    .A2(_0667_),
    .A3(_0668_),
    .B1(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__nor2_1 _2163_ (.A(_0987_),
    .B(_0670_),
    .Y(net421));
 sky130_fd_sc_hd__nand2_1 _2164_ (.A(_1142_),
    .B(net361),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _2165_ (.A(_1101_),
    .B(net264),
    .Y(_0672_));
 sky130_fd_sc_hd__o22ai_2 _2166_ (.A1(net324),
    .A2(_1060_),
    .B1(net286),
    .B2(_1061_),
    .Y(_0673_));
 sky130_fd_sc_hd__a31o_4 _2167_ (.A1(_1013_),
    .A2(_0671_),
    .A3(_0672_),
    .B1(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_1 _2168_ (.A(_0987_),
    .B(_0674_),
    .Y(net422));
 sky130_fd_sc_hd__nand2_1 _2169_ (.A(_1142_),
    .B(net362),
    .Y(_0675_));
 sky130_fd_sc_hd__nand2_1 _2170_ (.A(_1101_),
    .B(net265),
    .Y(_0676_));
 sky130_fd_sc_hd__o22ai_2 _2171_ (.A1(net325),
    .A2(_1060_),
    .B1(net287),
    .B2(_1021_),
    .Y(_0677_));
 sky130_fd_sc_hd__a31o_4 _2172_ (.A1(_1013_),
    .A2(_0675_),
    .A3(_0676_),
    .B1(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__nor2_1 _2173_ (.A(_0987_),
    .B(_0678_),
    .Y(net423));
 sky130_fd_sc_hd__a22o_1 _2174_ (.A1(_0996_),
    .A2(net266),
    .B1(net363),
    .B2(_1002_),
    .X(_0679_));
 sky130_fd_sc_hd__a221oi_2 _2175_ (.A1(net326),
    .A2(_0994_),
    .B1(net289),
    .B2(_0998_),
    .C1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nor2_1 _2176_ (.A(_0987_),
    .B(net733),
    .Y(net425));
 sky130_fd_sc_hd__a22o_1 _2177_ (.A1(_0996_),
    .A2(net267),
    .B1(net364),
    .B2(_1002_),
    .X(_0681_));
 sky130_fd_sc_hd__a221oi_2 _2178_ (.A1(net290),
    .A2(_0998_),
    .B1(net327),
    .B2(_0994_),
    .C1(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nor2_1 _2179_ (.A(_0987_),
    .B(net732),
    .Y(net426));
 sky130_fd_sc_hd__nand2_1 _2180_ (.A(_0993_),
    .B(net328),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _2181_ (.A(_0998_),
    .B(net291),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_2 _2182_ (.A(_0683_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__and3_1 _2183_ (.A(_0988_),
    .B(\arbiter.slave_sel[0][1] ),
    .C(net268),
    .X(_0686_));
 sky130_fd_sc_hd__nand2_1 _2184_ (.A(_0990_),
    .B(net231),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2b_2 _2185_ (.A_N(_0686_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nor2_4 _2186_ (.A(_0685_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__nor2_1 _2187_ (.A(_0987_),
    .B(_0689_),
    .Y(net427));
 sky130_fd_sc_hd__a22o_1 _2188_ (.A1(_0998_),
    .A2(net292),
    .B1(_1002_),
    .B2(net232),
    .X(_0690_));
 sky130_fd_sc_hd__a221oi_2 _2189_ (.A1(net329),
    .A2(_0994_),
    .B1(net269),
    .B2(_0996_),
    .C1(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__nor2_1 _2190_ (.A(_0987_),
    .B(net731),
    .Y(net428));
 sky130_fd_sc_hd__nand2_8 _2191_ (.A(_1096_),
    .B(_1083_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2_1 _2192_ (.A(_0692_),
    .B(net730),
    .Y(net429));
 sky130_fd_sc_hd__nor2_1 _2193_ (.A(_0692_),
    .B(net737),
    .Y(net430));
 sky130_fd_sc_hd__nor2_1 _2194_ (.A(_0692_),
    .B(net736),
    .Y(net431));
 sky130_fd_sc_hd__nor2_1 _2195_ (.A(_0692_),
    .B(_1008_),
    .Y(net432));
 sky130_fd_sc_hd__nor2_1 _2196_ (.A(_0692_),
    .B(net735),
    .Y(net433));
 sky130_fd_sc_hd__nor2_1 _2197_ (.A(_0692_),
    .B(net734),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _2198_ (.A(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__buf_4 _2199_ (.A(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__and2_1 _2200_ (.A(_1028_),
    .B(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__buf_1 _2201_ (.A(_0695_),
    .X(net436));
 sky130_fd_sc_hd__and2_1 _2202_ (.A(_1033_),
    .B(_0694_),
    .X(_0696_));
 sky130_fd_sc_hd__buf_1 _2203_ (.A(_0696_),
    .X(net437));
 sky130_fd_sc_hd__and2_1 _2204_ (.A(_1038_),
    .B(_0694_),
    .X(_0697_));
 sky130_fd_sc_hd__buf_1 _2205_ (.A(_0697_),
    .X(net438));
 sky130_fd_sc_hd__and2_1 _2206_ (.A(_1042_),
    .B(_0694_),
    .X(_0698_));
 sky130_fd_sc_hd__buf_1 _2207_ (.A(_0698_),
    .X(net439));
 sky130_fd_sc_hd__and2_1 _2208_ (.A(_1046_),
    .B(_0694_),
    .X(_0699_));
 sky130_fd_sc_hd__buf_1 _2209_ (.A(_0699_),
    .X(net440));
 sky130_fd_sc_hd__and2_1 _2210_ (.A(_1050_),
    .B(_0694_),
    .X(_0700_));
 sky130_fd_sc_hd__buf_1 _2211_ (.A(_0700_),
    .X(net441));
 sky130_fd_sc_hd__and2_1 _2212_ (.A(_1054_),
    .B(_0694_),
    .X(_0701_));
 sky130_fd_sc_hd__buf_1 _2213_ (.A(_0701_),
    .X(net442));
 sky130_fd_sc_hd__and2_1 _2214_ (.A(_1058_),
    .B(_0694_),
    .X(_0702_));
 sky130_fd_sc_hd__buf_1 _2215_ (.A(_0702_),
    .X(net443));
 sky130_fd_sc_hd__and2_1 _2216_ (.A(_1064_),
    .B(_0694_),
    .X(_0703_));
 sky130_fd_sc_hd__buf_1 _2217_ (.A(_0703_),
    .X(net444));
 sky130_fd_sc_hd__and2_1 _2218_ (.A(_1068_),
    .B(_0694_),
    .X(_0704_));
 sky130_fd_sc_hd__buf_1 _2219_ (.A(_0704_),
    .X(net445));
 sky130_fd_sc_hd__and2_1 _2220_ (.A(_1072_),
    .B(_0694_),
    .X(_0705_));
 sky130_fd_sc_hd__buf_1 _2221_ (.A(_0705_),
    .X(net447));
 sky130_fd_sc_hd__and2_1 _2222_ (.A(_1076_),
    .B(_0694_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_1 _2223_ (.A(_0706_),
    .X(net448));
 sky130_fd_sc_hd__and2_1 _2224_ (.A(_0102_),
    .B(_0694_),
    .X(_0707_));
 sky130_fd_sc_hd__buf_1 _2225_ (.A(_0707_),
    .X(net449));
 sky130_fd_sc_hd__and2_1 _2226_ (.A(_0201_),
    .B(_0694_),
    .X(_0708_));
 sky130_fd_sc_hd__buf_1 _2227_ (.A(_0708_),
    .X(net450));
 sky130_fd_sc_hd__and2_1 _2228_ (.A(_0389_),
    .B(_0694_),
    .X(_0709_));
 sky130_fd_sc_hd__buf_1 _2229_ (.A(_0709_),
    .X(net451));
 sky130_fd_sc_hd__and2_1 _2230_ (.A(_0502_),
    .B(_0694_),
    .X(_0710_));
 sky130_fd_sc_hd__buf_1 _2231_ (.A(_0710_),
    .X(net452));
 sky130_fd_sc_hd__and2_1 _2232_ (.A(_0612_),
    .B(_0693_),
    .X(_0711_));
 sky130_fd_sc_hd__buf_1 _2233_ (.A(_0711_),
    .X(net453));
 sky130_fd_sc_hd__and2_1 _2234_ (.A(_0653_),
    .B(_0693_),
    .X(_0712_));
 sky130_fd_sc_hd__buf_1 _2235_ (.A(_0712_),
    .X(net454));
 sky130_fd_sc_hd__and2_1 _2236_ (.A(_0657_),
    .B(_0693_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_1 _2237_ (.A(_0713_),
    .X(net455));
 sky130_fd_sc_hd__and2_1 _2238_ (.A(_0661_),
    .B(_0693_),
    .X(_0714_));
 sky130_fd_sc_hd__buf_1 _2239_ (.A(_0714_),
    .X(net456));
 sky130_fd_sc_hd__nor2_1 _2240_ (.A(_0692_),
    .B(_0666_),
    .Y(net458));
 sky130_fd_sc_hd__nor2_1 _2241_ (.A(_0692_),
    .B(_0670_),
    .Y(net459));
 sky130_fd_sc_hd__nor2_1 _2242_ (.A(_0692_),
    .B(_0674_),
    .Y(net460));
 sky130_fd_sc_hd__nor2_8 _2243_ (.A(\arbiter.slave_handled[2] ),
    .B(_1080_),
    .Y(_0715_));
 sky130_fd_sc_hd__clkinv_4 _2244_ (.A(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nand2_2 _2245_ (.A(_1002_),
    .B(_1083_),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_1 _2246_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__inv_2 _2247_ (.A(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_1 _2248_ (.A(_0719_),
    .B(_1100_),
    .Y(net518));
 sky130_fd_sc_hd__buf_4 _2249_ (.A(_0715_),
    .X(_0720_));
 sky130_fd_sc_hd__a2bb2o_1 _2250_ (.A1_N(_0504_),
    .A2_N(_1119_),
    .B1(_1116_),
    .B2(_0720_),
    .X(net519));
 sky130_fd_sc_hd__inv_2 _2251_ (.A(_1130_),
    .Y(_0721_));
 sky130_fd_sc_hd__buf_8 _2252_ (.A(_0716_),
    .X(_0722_));
 sky130_fd_sc_hd__o22ai_2 _2253_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0717_),
    .B2(_1158_),
    .Y(net520));
 sky130_fd_sc_hd__a2bb2o_1 _2254_ (.A1_N(_0504_),
    .A2_N(_1184_),
    .B1(_1153_),
    .B2(_0720_),
    .X(net521));
 sky130_fd_sc_hd__nor2_1 _2255_ (.A(_0692_),
    .B(_0678_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _2256_ (.A(_1182_),
    .Y(_0723_));
 sky130_fd_sc_hd__nor2_1 _2257_ (.A(_0722_),
    .B(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__a31o_1 _2258_ (.A1(_0015_),
    .A2(_0125_),
    .A3(_1182_),
    .B1(_0724_),
    .X(net522));
 sky130_fd_sc_hd__o22ai_2 _2259_ (.A1(_0722_),
    .A2(_0022_),
    .B1(_0485_),
    .B2(_0033_),
    .Y(net523));
 sky130_fd_sc_hd__a2bb2o_1 _2260_ (.A1_N(_0504_),
    .A2_N(_0040_),
    .B1(_0031_),
    .B2(_0720_),
    .X(net525));
 sky130_fd_sc_hd__clkinv_4 _2261_ (.A(_0717_),
    .Y(_0725_));
 sky130_fd_sc_hd__a22o_1 _2262_ (.A1(_0047_),
    .A2(_0715_),
    .B1(_0074_),
    .B2(_0725_),
    .X(net526));
 sky130_fd_sc_hd__a2bb2o_1 _2263_ (.A1_N(_0504_),
    .A2_N(_0095_),
    .B1(_0070_),
    .B2(_0720_),
    .X(net527));
 sky130_fd_sc_hd__o2bb2ai_2 _2264_ (.A1_N(_0110_),
    .A2_N(_0725_),
    .B1(_0092_),
    .B2(_0722_),
    .Y(net528));
 sky130_fd_sc_hd__inv_2 _2265_ (.A(_0106_),
    .Y(_0726_));
 sky130_fd_sc_hd__or3_1 _2266_ (.A(_0981_),
    .B(_1026_),
    .C(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__o21ai_2 _2267_ (.A1(_0726_),
    .A2(_0722_),
    .B1(_0727_),
    .Y(net529));
 sky130_fd_sc_hd__nand3_1 _2268_ (.A(_0140_),
    .B(_0125_),
    .C(_1197_),
    .Y(_0728_));
 sky130_fd_sc_hd__o22ai_4 _2269_ (.A1(_0722_),
    .A2(_1198_),
    .B1(_0485_),
    .B2(_0728_),
    .Y(net530));
 sky130_fd_sc_hd__o22ai_2 _2270_ (.A1(_0722_),
    .A2(_0139_),
    .B1(_0485_),
    .B2(_0148_),
    .Y(net531));
 sky130_fd_sc_hd__o22ai_2 _2271_ (.A1(_0722_),
    .A2(_0146_),
    .B1(_0485_),
    .B2(_0177_),
    .Y(net532));
 sky130_fd_sc_hd__nor2_1 _2272_ (.A(_0692_),
    .B(net733),
    .Y(net462));
 sky130_fd_sc_hd__o22ai_4 _2273_ (.A1(_0722_),
    .A2(_0058_),
    .B1(_0485_),
    .B2(_0165_),
    .Y(net533));
 sky130_fd_sc_hd__inv_2 _2274_ (.A(_0079_),
    .Y(_0729_));
 sky130_fd_sc_hd__o22ai_4 _2275_ (.A1(_0722_),
    .A2(_0729_),
    .B1(_0485_),
    .B2(_0080_),
    .Y(net534));
 sky130_fd_sc_hd__inv_2 _2276_ (.A(_0174_),
    .Y(_0730_));
 sky130_fd_sc_hd__o22ai_2 _2277_ (.A1(_0722_),
    .A2(_0730_),
    .B1(_0485_),
    .B2(_0183_),
    .Y(net536));
 sky130_fd_sc_hd__inv_2 _2278_ (.A(_0115_),
    .Y(_0731_));
 sky130_fd_sc_hd__o22ai_2 _2279_ (.A1(_0716_),
    .A2(_0731_),
    .B1(_0485_),
    .B2(_0116_),
    .Y(net537));
 sky130_fd_sc_hd__o2bb2ai_2 _2280_ (.A1_N(_0124_),
    .A2_N(_0720_),
    .B1(_0504_),
    .B2(_0126_),
    .Y(net538));
 sky130_fd_sc_hd__a22o_1 _2281_ (.A1(_0196_),
    .A2(_0715_),
    .B1(_0213_),
    .B2(_0725_),
    .X(net539));
 sky130_fd_sc_hd__inv_2 _2282_ (.A(_0211_),
    .Y(_0732_));
 sky130_fd_sc_hd__nand3_1 _2283_ (.A(_0211_),
    .B(_1142_),
    .C(_1013_),
    .Y(_0733_));
 sky130_fd_sc_hd__o22ai_2 _2284_ (.A1(_0716_),
    .A2(_0732_),
    .B1(_0485_),
    .B2(_0733_),
    .Y(net540));
 sky130_fd_sc_hd__a2bb2o_1 _2285_ (.A1_N(_0504_),
    .A2_N(_0161_),
    .B1(_0160_),
    .B2(_0720_),
    .X(net541));
 sky130_fd_sc_hd__a22o_1 _2286_ (.A1(_0277_),
    .A2(_0715_),
    .B1(_0290_),
    .B2(_0725_),
    .X(net542));
 sky130_fd_sc_hd__inv_2 _2287_ (.A(_0287_),
    .Y(_0734_));
 sky130_fd_sc_hd__o22ai_2 _2288_ (.A1(_0716_),
    .A2(_0734_),
    .B1(_0485_),
    .B2(_0300_),
    .Y(net543));
 sky130_fd_sc_hd__nor2_1 _2289_ (.A(_0692_),
    .B(net732),
    .Y(net463));
 sky130_fd_sc_hd__o22ai_2 _2290_ (.A1(_0716_),
    .A2(_0299_),
    .B1(_0485_),
    .B2(_0314_),
    .Y(net544));
 sky130_fd_sc_hd__a2bb2o_1 _2291_ (.A1_N(_0504_),
    .A2_N(_0318_),
    .B1(_0311_),
    .B2(_0720_),
    .X(net545));
 sky130_fd_sc_hd__inv_2 _2292_ (.A(_0327_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _2293_ (.A(_0722_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__a31o_1 _2294_ (.A1(_0015_),
    .A2(_0125_),
    .A3(_0327_),
    .B1(_0736_),
    .X(net547));
 sky130_fd_sc_hd__a22o_1 _2295_ (.A1(_0244_),
    .A2(_0715_),
    .B1(_0375_),
    .B2(_0725_),
    .X(net548));
 sky130_fd_sc_hd__a2bb2o_1 _2296_ (.A1_N(_0504_),
    .A2_N(_0233_),
    .B1(_0232_),
    .B2(_0720_),
    .X(net549));
 sky130_fd_sc_hd__a22o_1 _2297_ (.A1(_0254_),
    .A2(_0715_),
    .B1(_0266_),
    .B2(_0725_),
    .X(net550));
 sky130_fd_sc_hd__a22o_1 _2298_ (.A1(_0264_),
    .A2(_0715_),
    .B1(_0401_),
    .B2(_0725_),
    .X(net551));
 sky130_fd_sc_hd__a22o_1 _2299_ (.A1(_0398_),
    .A2(_0715_),
    .B1(_0405_),
    .B2(_0725_),
    .X(net552));
 sky130_fd_sc_hd__a22o_1 _2300_ (.A1(_0363_),
    .A2(_0715_),
    .B1(_0436_),
    .B2(_0725_),
    .X(net553));
 sky130_fd_sc_hd__a2bb2o_1 _2301_ (.A1_N(_0504_),
    .A2_N(_0342_),
    .B1(_0341_),
    .B2(_0720_),
    .X(net554));
 sky130_fd_sc_hd__nor2_1 _2302_ (.A(_0692_),
    .B(_0689_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _2303_ (.A(_0351_),
    .Y(_0737_));
 sky130_fd_sc_hd__nor2_1 _2304_ (.A(_0722_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__a31o_1 _2305_ (.A1(_0015_),
    .A2(_0125_),
    .A3(_0351_),
    .B1(_0738_),
    .X(net555));
 sky130_fd_sc_hd__o2bb2ai_2 _2306_ (.A1_N(_0373_),
    .A2_N(_0720_),
    .B1(_0504_),
    .B2(_0374_),
    .Y(net556));
 sky130_fd_sc_hd__a22o_1 _2307_ (.A1(_0476_),
    .A2(_0715_),
    .B1(_0488_),
    .B2(_0725_),
    .X(net558));
 sky130_fd_sc_hd__o22ai_2 _2308_ (.A1(_0716_),
    .A2(_0484_),
    .B1(_0485_),
    .B2(_0491_),
    .Y(net559));
 sky130_fd_sc_hd__a2bb2o_1 _2309_ (.A1_N(_0504_),
    .A2_N(_0497_),
    .B1(_0414_),
    .B2(_0720_),
    .X(net560));
 sky130_fd_sc_hd__o22ai_4 _2310_ (.A1(_0716_),
    .A2(_0494_),
    .B1(_0485_),
    .B2(_0429_),
    .Y(net561));
 sky130_fd_sc_hd__a2bb2o_1 _2311_ (.A1_N(_0981_),
    .A2_N(_0439_),
    .B1(_0422_),
    .B2(_0720_),
    .X(net562));
 sky130_fd_sc_hd__a2bb2o_1 _2312_ (.A1_N(_0981_),
    .A2_N(_0464_),
    .B1(_0448_),
    .B2(_0720_),
    .X(net563));
 sky130_fd_sc_hd__inv_2 _2313_ (.A(_0462_),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2_1 _2314_ (.A(_0722_),
    .B(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__a31o_1 _2315_ (.A1(_0015_),
    .A2(_0125_),
    .A3(_0462_),
    .B1(_0740_),
    .X(net564));
 sky130_fd_sc_hd__a22o_1 _2316_ (.A1(_0542_),
    .A2(_0715_),
    .B1(_0553_),
    .B2(_0725_),
    .X(net565));
 sky130_fd_sc_hd__nor2_1 _2317_ (.A(_0692_),
    .B(net731),
    .Y(net465));
 sky130_fd_sc_hd__a2bb2o_1 _2318_ (.A1_N(_0981_),
    .A2_N(_0572_),
    .B1(_0550_),
    .B2(_0720_),
    .X(net566));
 sky130_fd_sc_hd__a22o_1 _2319_ (.A1(_0570_),
    .A2(_0715_),
    .B1(_0585_),
    .B2(_0725_),
    .X(net567));
 sky130_fd_sc_hd__inv_2 _2320_ (.A(_0583_),
    .Y(_0741_));
 sky130_fd_sc_hd__nor2_1 _2321_ (.A(_0722_),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__a31o_1 _2322_ (.A1(_0015_),
    .A2(_0125_),
    .A3(_0583_),
    .B1(_0742_),
    .X(net569));
 sky130_fd_sc_hd__nor2_1 _2323_ (.A(_0722_),
    .B(_0595_),
    .Y(_0743_));
 sky130_fd_sc_hd__a31o_1 _2324_ (.A1(_0015_),
    .A2(_0125_),
    .A3(_0526_),
    .B1(_0743_),
    .X(net570));
 sky130_fd_sc_hd__a2bb2o_1 _2325_ (.A1_N(_0981_),
    .A2_N(_0513_),
    .B1(_0512_),
    .B2(_0720_),
    .X(net571));
 sky130_fd_sc_hd__a2bb2o_1 _2326_ (.A1_N(_0981_),
    .A2_N(_0619_),
    .B1(_0520_),
    .B2(_0720_),
    .X(net572));
 sky130_fd_sc_hd__inv_2 _2327_ (.A(_0617_),
    .Y(_0744_));
 sky130_fd_sc_hd__nor2_1 _2328_ (.A(_0719_),
    .B(_0744_),
    .Y(net573));
 sky130_fd_sc_hd__inv_2 _2329_ (.A(_0559_),
    .Y(_0745_));
 sky130_fd_sc_hd__nor2_1 _2330_ (.A(_0719_),
    .B(_0745_),
    .Y(net574));
 sky130_fd_sc_hd__inv_2 _2331_ (.A(_0632_),
    .Y(_0746_));
 sky130_fd_sc_hd__nor2_1 _2332_ (.A(_0719_),
    .B(_0746_),
    .Y(net575));
 sky130_fd_sc_hd__nor2_1 _2333_ (.A(_0719_),
    .B(_0637_),
    .Y(net576));
 sky130_fd_sc_hd__nand2_8 _2334_ (.A(_1091_),
    .B(_1083_),
    .Y(_0747_));
 sky130_fd_sc_hd__nor2_1 _2335_ (.A(_0747_),
    .B(net730),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _2336_ (.A(_0640_),
    .Y(_0748_));
 sky130_fd_sc_hd__nor2_1 _2337_ (.A(_0719_),
    .B(_0748_),
    .Y(net577));
 sky130_fd_sc_hd__nor2_1 _2338_ (.A(_0719_),
    .B(_0650_),
    .Y(net578));
 sky130_fd_sc_hd__nor2_1 _2339_ (.A(_0719_),
    .B(_0606_),
    .Y(net580));
 sky130_fd_sc_hd__nor2_1 _2340_ (.A(_0747_),
    .B(net737),
    .Y(net467));
 sky130_fd_sc_hd__nor2_1 _2341_ (.A(_0747_),
    .B(net736),
    .Y(net469));
 sky130_fd_sc_hd__nor2_1 _2342_ (.A(_0747_),
    .B(_1008_),
    .Y(net470));
 sky130_fd_sc_hd__nor2_1 _2343_ (.A(_0747_),
    .B(net735),
    .Y(net471));
 sky130_fd_sc_hd__nor2_1 _2344_ (.A(_0747_),
    .B(net734),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _2345_ (.A(_0747_),
    .Y(_0749_));
 sky130_fd_sc_hd__clkbuf_4 _2346_ (.A(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__and2_1 _2347_ (.A(_1028_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__buf_1 _2348_ (.A(_0751_),
    .X(net473));
 sky130_fd_sc_hd__and2_1 _2349_ (.A(_1033_),
    .B(_0750_),
    .X(_0752_));
 sky130_fd_sc_hd__buf_1 _2350_ (.A(_0752_),
    .X(net474));
 sky130_fd_sc_hd__and2_1 _2351_ (.A(_1038_),
    .B(_0750_),
    .X(_0753_));
 sky130_fd_sc_hd__buf_1 _2352_ (.A(_0753_),
    .X(net475));
 sky130_fd_sc_hd__and2_1 _2353_ (.A(_1042_),
    .B(_0750_),
    .X(_0754_));
 sky130_fd_sc_hd__buf_1 _2354_ (.A(_0754_),
    .X(net476));
 sky130_fd_sc_hd__and2_1 _2355_ (.A(_1046_),
    .B(_0750_),
    .X(_0755_));
 sky130_fd_sc_hd__buf_1 _2356_ (.A(_0755_),
    .X(net477));
 sky130_fd_sc_hd__and2_1 _2357_ (.A(_1050_),
    .B(_0750_),
    .X(_0756_));
 sky130_fd_sc_hd__buf_1 _2358_ (.A(_0756_),
    .X(net478));
 sky130_fd_sc_hd__and2_1 _2359_ (.A(_1054_),
    .B(_0750_),
    .X(_0757_));
 sky130_fd_sc_hd__buf_1 _2360_ (.A(_0757_),
    .X(net480));
 sky130_fd_sc_hd__and2_1 _2361_ (.A(_1058_),
    .B(_0750_),
    .X(_0758_));
 sky130_fd_sc_hd__buf_1 _2362_ (.A(_0758_),
    .X(net481));
 sky130_fd_sc_hd__and2_1 _2363_ (.A(_1064_),
    .B(_0750_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_1 _2364_ (.A(_0759_),
    .X(net482));
 sky130_fd_sc_hd__and2_1 _2365_ (.A(_1068_),
    .B(_0750_),
    .X(_0760_));
 sky130_fd_sc_hd__buf_1 _2366_ (.A(_0760_),
    .X(net483));
 sky130_fd_sc_hd__and2_1 _2367_ (.A(_1072_),
    .B(_0750_),
    .X(_0761_));
 sky130_fd_sc_hd__buf_1 _2368_ (.A(_0761_),
    .X(net484));
 sky130_fd_sc_hd__and2_1 _2369_ (.A(_1076_),
    .B(_0750_),
    .X(_0762_));
 sky130_fd_sc_hd__buf_1 _2370_ (.A(_0762_),
    .X(net485));
 sky130_fd_sc_hd__and2_1 _2371_ (.A(_0102_),
    .B(_0750_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_1 _2372_ (.A(_0763_),
    .X(net486));
 sky130_fd_sc_hd__and2_1 _2373_ (.A(_0201_),
    .B(_0750_),
    .X(_0764_));
 sky130_fd_sc_hd__buf_1 _2374_ (.A(_0764_),
    .X(net487));
 sky130_fd_sc_hd__and2_1 _2375_ (.A(_0389_),
    .B(_0750_),
    .X(_0765_));
 sky130_fd_sc_hd__buf_1 _2376_ (.A(_0765_),
    .X(net488));
 sky130_fd_sc_hd__and2_1 _2377_ (.A(_0502_),
    .B(_0750_),
    .X(_0766_));
 sky130_fd_sc_hd__buf_1 _2378_ (.A(_0766_),
    .X(net489));
 sky130_fd_sc_hd__and2_1 _2379_ (.A(_0612_),
    .B(_0749_),
    .X(_0767_));
 sky130_fd_sc_hd__buf_1 _2380_ (.A(_0767_),
    .X(net491));
 sky130_fd_sc_hd__and2_1 _2381_ (.A(_0653_),
    .B(_0749_),
    .X(_0768_));
 sky130_fd_sc_hd__buf_1 _2382_ (.A(_0768_),
    .X(net492));
 sky130_fd_sc_hd__nor2_4 _2383_ (.A(\arbiter.slave_handled[3] ),
    .B(_1080_),
    .Y(_0769_));
 sky130_fd_sc_hd__inv_4 _2384_ (.A(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__o22ai_2 _2385_ (.A1(_0770_),
    .A2(_1100_),
    .B1(_0485_),
    .B2(_1137_),
    .Y(net581));
 sky130_fd_sc_hd__buf_8 _2386_ (.A(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_1 _2387_ (.A(_0771_),
    .B(_1117_),
    .Y(_0772_));
 sky130_fd_sc_hd__a31o_1 _2388_ (.A1(_1157_),
    .A2(_1083_),
    .A3(_0094_),
    .B1(_0772_),
    .X(net582));
 sky130_fd_sc_hd__o22ai_4 _2389_ (.A1(_0770_),
    .A2(_0721_),
    .B1(_0504_),
    .B2(_1173_),
    .Y(net583));
 sky130_fd_sc_hd__inv_2 _2390_ (.A(_1153_),
    .Y(_0773_));
 sky130_fd_sc_hd__nor2_4 _2391_ (.A(_0981_),
    .B(_0995_),
    .Y(_0774_));
 sky130_fd_sc_hd__clkinv_4 _2392_ (.A(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_1 _2393_ (.A(_0770_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__clkinv_4 _2394_ (.A(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__nor2_1 _2395_ (.A(_0773_),
    .B(_0777_),
    .Y(net584));
 sky130_fd_sc_hd__nor2_1 _2396_ (.A(_0771_),
    .B(_0723_),
    .Y(_0778_));
 sky130_fd_sc_hd__a31o_2 _2397_ (.A1(_1185_),
    .A2(_1083_),
    .A3(_0094_),
    .B1(_0778_),
    .X(net585));
 sky130_fd_sc_hd__nor2_1 _2398_ (.A(_0777_),
    .B(_0022_),
    .Y(net586));
 sky130_fd_sc_hd__buf_4 _2399_ (.A(_0774_),
    .X(_0779_));
 sky130_fd_sc_hd__nand2_1 _2400_ (.A(_0081_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__o21ai_4 _2401_ (.A1(_0032_),
    .A2(_0771_),
    .B1(_0780_),
    .Y(net587));
 sky130_fd_sc_hd__and2_1 _2402_ (.A(_0657_),
    .B(_0749_),
    .X(_0781_));
 sky130_fd_sc_hd__buf_1 _2403_ (.A(_0781_),
    .X(net493));
 sky130_fd_sc_hd__inv_2 _2404_ (.A(_0047_),
    .Y(_0782_));
 sky130_fd_sc_hd__o22ai_4 _2405_ (.A1(_0782_),
    .A2(_0771_),
    .B1(_0775_),
    .B2(_0099_),
    .Y(net588));
 sky130_fd_sc_hd__nand2_1 _2406_ (.A(_0117_),
    .B(_0779_),
    .Y(_0783_));
 sky130_fd_sc_hd__clkbuf_4 _2407_ (.A(_0769_),
    .X(_0784_));
 sky130_fd_sc_hd__nand2_1 _2408_ (.A(_0070_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__nand2_1 _2409_ (.A(_0783_),
    .B(_0785_),
    .Y(net589));
 sky130_fd_sc_hd__nor2_1 _2410_ (.A(_0771_),
    .B(_0092_),
    .Y(_0786_));
 sky130_fd_sc_hd__a31o_2 _2411_ (.A1(_0097_),
    .A2(_1083_),
    .A3(_0094_),
    .B1(_0786_),
    .X(net591));
 sky130_fd_sc_hd__nor2_1 _2412_ (.A(_0726_),
    .B(_0777_),
    .Y(net592));
 sky130_fd_sc_hd__nor2_1 _2413_ (.A(_1198_),
    .B(_0777_),
    .Y(net593));
 sky130_fd_sc_hd__o21ai_2 _2414_ (.A1(_1024_),
    .A2(_0138_),
    .B1(_1022_),
    .Y(_0787_));
 sky130_fd_sc_hd__o22ai_4 _2415_ (.A1(_0139_),
    .A2(_0771_),
    .B1(_0775_),
    .B2(_0787_),
    .Y(net594));
 sky130_fd_sc_hd__nor2_1 _2416_ (.A(_0777_),
    .B(_0146_),
    .Y(net595));
 sky130_fd_sc_hd__and2_1 _2417_ (.A(_0177_),
    .B(_0178_),
    .X(_0788_));
 sky130_fd_sc_hd__o22ai_4 _2418_ (.A1(_0058_),
    .A2(_0771_),
    .B1(_0775_),
    .B2(_0788_),
    .Y(net596));
 sky130_fd_sc_hd__nand3_1 _2419_ (.A(_0182_),
    .B(_0185_),
    .C(_0779_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2_1 _2420_ (.A(_0079_),
    .B(_0784_),
    .Y(_0790_));
 sky130_fd_sc_hd__nand2_1 _2421_ (.A(_0789_),
    .B(_0790_),
    .Y(net597));
 sky130_fd_sc_hd__nand2_1 _2422_ (.A(_0080_),
    .B(_0175_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand3_1 _2423_ (.A(_0791_),
    .B(_0015_),
    .C(_0094_),
    .Y(_0792_));
 sky130_fd_sc_hd__o21ai_4 _2424_ (.A1(_0730_),
    .A2(_0771_),
    .B1(_0792_),
    .Y(net598));
 sky130_fd_sc_hd__and2_1 _2425_ (.A(_0661_),
    .B(_0749_),
    .X(_0793_));
 sky130_fd_sc_hd__buf_1 _2426_ (.A(_0793_),
    .X(net494));
 sky130_fd_sc_hd__nand2_1 _2427_ (.A(_0183_),
    .B(_0184_),
    .Y(_0794_));
 sky130_fd_sc_hd__nand3_1 _2428_ (.A(_0794_),
    .B(_0015_),
    .C(_0094_),
    .Y(_0795_));
 sky130_fd_sc_hd__o21ai_2 _2429_ (.A1(_0771_),
    .A2(_0731_),
    .B1(_0795_),
    .Y(net599));
 sky130_fd_sc_hd__nor2_1 _2430_ (.A(_0777_),
    .B(_0188_),
    .Y(net600));
 sky130_fd_sc_hd__nor2_1 _2431_ (.A(_0777_),
    .B(_0197_),
    .Y(net602));
 sky130_fd_sc_hd__a2bb2o_1 _2432_ (.A1_N(_0981_),
    .A2_N(_0281_),
    .B1(_0211_),
    .B2(_0784_),
    .X(net603));
 sky130_fd_sc_hd__nor2_1 _2433_ (.A(_0219_),
    .B(_0777_),
    .Y(net604));
 sky130_fd_sc_hd__inv_2 _2434_ (.A(_0277_),
    .Y(_0796_));
 sky130_fd_sc_hd__nand3_1 _2435_ (.A(_0302_),
    .B(_0303_),
    .C(_0774_),
    .Y(_0797_));
 sky130_fd_sc_hd__o21ai_2 _2436_ (.A1(_0796_),
    .A2(_0771_),
    .B1(_0797_),
    .Y(net605));
 sky130_fd_sc_hd__nand3_1 _2437_ (.A(_0316_),
    .B(_0313_),
    .C(_0774_),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_2 _2438_ (.A1(_0734_),
    .A2(_0771_),
    .B1(_0798_),
    .Y(net606));
 sky130_fd_sc_hd__o22ai_4 _2439_ (.A1(_0770_),
    .A2(_0299_),
    .B1(_0504_),
    .B2(_0331_),
    .Y(net607));
 sky130_fd_sc_hd__nor2_1 _2440_ (.A(_0771_),
    .B(_0312_),
    .Y(_0799_));
 sky130_fd_sc_hd__a31o_1 _2441_ (.A1(_1083_),
    .A2(_1136_),
    .A3(_0311_),
    .B1(_0799_),
    .X(net608));
 sky130_fd_sc_hd__nand2_1 _2442_ (.A(_0378_),
    .B(_0779_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _2443_ (.A(_0327_),
    .B(_0784_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_1 _2444_ (.A(_0800_),
    .B(_0801_),
    .Y(net609));
 sky130_fd_sc_hd__nor2_1 _2445_ (.A(_0747_),
    .B(_0666_),
    .Y(net495));
 sky130_fd_sc_hd__nor2_1 _2446_ (.A(_0777_),
    .B(_0368_),
    .Y(net610));
 sky130_fd_sc_hd__nand2_1 _2447_ (.A(_0245_),
    .B(_0246_),
    .Y(_0802_));
 sky130_fd_sc_hd__a22o_1 _2448_ (.A1(_0232_),
    .A2(_0769_),
    .B1(_0802_),
    .B2(_0779_),
    .X(net611));
 sky130_fd_sc_hd__a22o_1 _2449_ (.A1(_0254_),
    .A2(_0769_),
    .B1(_0383_),
    .B2(_0779_),
    .X(net614));
 sky130_fd_sc_hd__nand3_1 _2450_ (.A(_0407_),
    .B(_0430_),
    .C(_0779_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_1 _2451_ (.A(_0264_),
    .B(_0784_),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_1 _2452_ (.A(_0803_),
    .B(_0804_),
    .Y(net615));
 sky130_fd_sc_hd__nand3_1 _2453_ (.A(_0438_),
    .B(_0453_),
    .C(_0779_),
    .Y(_0805_));
 sky130_fd_sc_hd__nand2_1 _2454_ (.A(_0398_),
    .B(_0784_),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2_1 _2455_ (.A(_0805_),
    .B(_0806_),
    .Y(net616));
 sky130_fd_sc_hd__a2bb2o_1 _2456_ (.A1_N(_0981_),
    .A2_N(_0364_),
    .B1(_0363_),
    .B2(_0784_),
    .X(net617));
 sky130_fd_sc_hd__inv_2 _2457_ (.A(_0341_),
    .Y(_0807_));
 sky130_fd_sc_hd__nor2_1 _2458_ (.A(_0771_),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__a31o_1 _2459_ (.A1(_1083_),
    .A2(_1136_),
    .A3(_0341_),
    .B1(_0808_),
    .X(net618));
 sky130_fd_sc_hd__a22o_1 _2460_ (.A1(_0351_),
    .A2(_0769_),
    .B1(_0353_),
    .B2(_0779_),
    .X(net619));
 sky130_fd_sc_hd__nand3_1 _2461_ (.A(_0373_),
    .B(_0015_),
    .C(_1136_),
    .Y(_0809_));
 sky130_fd_sc_hd__o21ai_2 _2462_ (.A1(_0771_),
    .A2(_0472_),
    .B1(_0809_),
    .Y(net620));
 sky130_fd_sc_hd__nand2_1 _2463_ (.A(_0478_),
    .B(_0779_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _2464_ (.A(_0476_),
    .B(_0784_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _2465_ (.A(_0810_),
    .B(_0811_),
    .Y(net621));
 sky130_fd_sc_hd__nor2_1 _2466_ (.A(_0747_),
    .B(_0670_),
    .Y(net496));
 sky130_fd_sc_hd__nand3_1 _2467_ (.A(_0495_),
    .B(_0498_),
    .C(_0774_),
    .Y(_0812_));
 sky130_fd_sc_hd__o21ai_2 _2468_ (.A1(_0484_),
    .A2(_0771_),
    .B1(_0812_),
    .Y(net622));
 sky130_fd_sc_hd__a2bb2o_1 _2469_ (.A1_N(_0981_),
    .A2_N(_0415_),
    .B1(_0414_),
    .B2(_0784_),
    .X(net623));
 sky130_fd_sc_hd__o22ai_4 _2470_ (.A1(_0770_),
    .A2(_0494_),
    .B1(_0504_),
    .B2(_0452_),
    .Y(net625));
 sky130_fd_sc_hd__a2bb2o_1 _2471_ (.A1_N(_0981_),
    .A2_N(_0467_),
    .B1(_0422_),
    .B2(_0784_),
    .X(net626));
 sky130_fd_sc_hd__inv_2 _2472_ (.A(_0448_),
    .Y(_0813_));
 sky130_fd_sc_hd__nor2_1 _2473_ (.A(_0034_),
    .B(_0450_),
    .Y(_0814_));
 sky130_fd_sc_hd__o22ai_4 _2474_ (.A1(_0813_),
    .A2(_0771_),
    .B1(_0775_),
    .B2(_0814_),
    .Y(net627));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(_0561_),
    .B(_0779_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_1 _2476_ (.A(_0462_),
    .B(_0784_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand2_1 _2477_ (.A(_0815_),
    .B(_0816_),
    .Y(net628));
 sky130_fd_sc_hd__nor2_1 _2478_ (.A(_0770_),
    .B(_0543_),
    .Y(_0817_));
 sky130_fd_sc_hd__a31o_1 _2479_ (.A1(_1083_),
    .A2(_1136_),
    .A3(_0542_),
    .B1(_0817_),
    .X(net629));
 sky130_fd_sc_hd__nand2_1 _2480_ (.A(_0592_),
    .B(_0779_),
    .Y(_0818_));
 sky130_fd_sc_hd__nand2_1 _2481_ (.A(_0550_),
    .B(_0784_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _2482_ (.A(_0818_),
    .B(_0819_),
    .Y(net630));
 sky130_fd_sc_hd__o21a_1 _2483_ (.A1(_0774_),
    .A2(_0784_),
    .B1(_0570_),
    .X(net631));
 sky130_fd_sc_hd__nor2_1 _2484_ (.A(_0770_),
    .B(_0741_),
    .Y(_0820_));
 sky130_fd_sc_hd__a31o_1 _2485_ (.A1(_1083_),
    .A2(_1136_),
    .A3(_0583_),
    .B1(_0820_),
    .X(net632));
 sky130_fd_sc_hd__nor2_1 _2486_ (.A(_0747_),
    .B(_0674_),
    .Y(net497));
 sky130_fd_sc_hd__o22ai_4 _2487_ (.A1(_0770_),
    .A2(_0595_),
    .B1(_0504_),
    .B2(_0527_),
    .Y(net633));
 sky130_fd_sc_hd__nor2_1 _2488_ (.A(_0777_),
    .B(_0596_),
    .Y(net634));
 sky130_fd_sc_hd__a22o_1 _2489_ (.A1(_0520_),
    .A2(_0769_),
    .B1(_0522_),
    .B2(_0779_),
    .X(net636));
 sky130_fd_sc_hd__nand2_1 _2490_ (.A(_0620_),
    .B(_0779_),
    .Y(_0821_));
 sky130_fd_sc_hd__nand2_1 _2491_ (.A(_0617_),
    .B(_0784_),
    .Y(_0822_));
 sky130_fd_sc_hd__nand2_1 _2492_ (.A(_0821_),
    .B(_0822_),
    .Y(net637));
 sky130_fd_sc_hd__nand2_1 _2493_ (.A(_0625_),
    .B(_0779_),
    .Y(_0823_));
 sky130_fd_sc_hd__nand2_1 _2494_ (.A(_0559_),
    .B(_0784_),
    .Y(_0824_));
 sky130_fd_sc_hd__nand2_2 _2495_ (.A(_0823_),
    .B(_0824_),
    .Y(net638));
 sky130_fd_sc_hd__nor2_1 _2496_ (.A(_0777_),
    .B(_0746_),
    .Y(net639));
 sky130_fd_sc_hd__nor2_1 _2497_ (.A(_0777_),
    .B(_0637_),
    .Y(net640));
 sky130_fd_sc_hd__nand2_1 _2498_ (.A(_0649_),
    .B(_1022_),
    .Y(_0825_));
 sky130_fd_sc_hd__nand2_1 _2499_ (.A(_0825_),
    .B(_1142_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand2_1 _2500_ (.A(_0605_),
    .B(_1022_),
    .Y(_0827_));
 sky130_fd_sc_hd__nand2_1 _2501_ (.A(_0827_),
    .B(_1102_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _2502_ (.A(_0826_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__nand2_1 _2503_ (.A(_0829_),
    .B(_0034_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand3_1 _2504_ (.A(_0591_),
    .B(_0641_),
    .C(_0094_),
    .Y(_0831_));
 sky130_fd_sc_hd__nand3_1 _2505_ (.A(_0830_),
    .B(_0831_),
    .C(_0779_),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_1 _2506_ (.A(_0640_),
    .B(_0784_),
    .Y(_0833_));
 sky130_fd_sc_hd__nand2_2 _2507_ (.A(_0832_),
    .B(_0833_),
    .Y(net641));
 sky130_fd_sc_hd__nor2_1 _2508_ (.A(_0777_),
    .B(_0650_),
    .Y(net642));
 sky130_fd_sc_hd__nor2_1 _2509_ (.A(_0777_),
    .B(_0606_),
    .Y(net643));
 sky130_fd_sc_hd__nor2_1 _2510_ (.A(_0747_),
    .B(_0678_),
    .Y(net498));
 sky130_fd_sc_hd__nor2_1 _2511_ (.A(_0747_),
    .B(net733),
    .Y(net499));
 sky130_fd_sc_hd__nor2_1 _2512_ (.A(_0747_),
    .B(net732),
    .Y(net500));
 sky130_fd_sc_hd__nor2_1 _2513_ (.A(_0747_),
    .B(_0689_),
    .Y(net367));
 sky130_fd_sc_hd__nor2_1 _2514_ (.A(_0747_),
    .B(net731),
    .Y(net368));
 sky130_fd_sc_hd__nor2_4 _2515_ (.A(_0981_),
    .B(_1087_),
    .Y(_0834_));
 sky130_fd_sc_hd__clkinv_4 _2516_ (.A(_0834_),
    .Y(_0835_));
 sky130_fd_sc_hd__nor2_1 _2517_ (.A(_0835_),
    .B(net730),
    .Y(net369));
 sky130_fd_sc_hd__nor2_1 _2518_ (.A(_0835_),
    .B(net737),
    .Y(net370));
 sky130_fd_sc_hd__nor2_1 _2519_ (.A(_0835_),
    .B(net736),
    .Y(net371));
 sky130_fd_sc_hd__nor2_1 _2520_ (.A(_0835_),
    .B(_1008_),
    .Y(net372));
 sky130_fd_sc_hd__nor2_1 _2521_ (.A(_0835_),
    .B(net735),
    .Y(net373));
 sky130_fd_sc_hd__nor2_1 _2522_ (.A(_0835_),
    .B(net734),
    .Y(net374));
 sky130_fd_sc_hd__clkbuf_4 _2523_ (.A(_0834_),
    .X(_0836_));
 sky130_fd_sc_hd__and2_1 _2524_ (.A(_1028_),
    .B(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__buf_1 _2525_ (.A(_0837_),
    .X(net375));
 sky130_fd_sc_hd__and2_1 _2526_ (.A(_1033_),
    .B(_0836_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_1 _2527_ (.A(_0838_),
    .X(net376));
 sky130_fd_sc_hd__and2_1 _2528_ (.A(_1038_),
    .B(_0836_),
    .X(_0839_));
 sky130_fd_sc_hd__buf_1 _2529_ (.A(_0839_),
    .X(net378));
 sky130_fd_sc_hd__and2_1 _2530_ (.A(_1042_),
    .B(_0836_),
    .X(_0840_));
 sky130_fd_sc_hd__buf_1 _2531_ (.A(_0840_),
    .X(net379));
 sky130_fd_sc_hd__and2_1 _2532_ (.A(_1046_),
    .B(_0836_),
    .X(_0841_));
 sky130_fd_sc_hd__buf_1 _2533_ (.A(_0841_),
    .X(net380));
 sky130_fd_sc_hd__and2_1 _2534_ (.A(_1050_),
    .B(_0836_),
    .X(_0842_));
 sky130_fd_sc_hd__buf_1 _2535_ (.A(_0842_),
    .X(net381));
 sky130_fd_sc_hd__and2_1 _2536_ (.A(_1054_),
    .B(_0836_),
    .X(_0843_));
 sky130_fd_sc_hd__buf_1 _2537_ (.A(_0843_),
    .X(net382));
 sky130_fd_sc_hd__and2_1 _2538_ (.A(_1058_),
    .B(_0836_),
    .X(_0844_));
 sky130_fd_sc_hd__buf_1 _2539_ (.A(_0844_),
    .X(net383));
 sky130_fd_sc_hd__and2_1 _2540_ (.A(_1064_),
    .B(_0836_),
    .X(_0845_));
 sky130_fd_sc_hd__buf_1 _2541_ (.A(_0845_),
    .X(net384));
 sky130_fd_sc_hd__and2_1 _2542_ (.A(_1068_),
    .B(_0836_),
    .X(_0846_));
 sky130_fd_sc_hd__buf_1 _2543_ (.A(_0846_),
    .X(net385));
 sky130_fd_sc_hd__and2_1 _2544_ (.A(_1072_),
    .B(_0836_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_1 _2545_ (.A(_0847_),
    .X(net386));
 sky130_fd_sc_hd__and2_1 _2546_ (.A(_1076_),
    .B(_0836_),
    .X(_0848_));
 sky130_fd_sc_hd__buf_1 _2547_ (.A(_0848_),
    .X(net387));
 sky130_fd_sc_hd__and2_1 _2548_ (.A(_0102_),
    .B(_0836_),
    .X(_0849_));
 sky130_fd_sc_hd__buf_1 _2549_ (.A(_0849_),
    .X(net389));
 sky130_fd_sc_hd__and2_1 _2550_ (.A(_0201_),
    .B(_0836_),
    .X(_0850_));
 sky130_fd_sc_hd__buf_1 _2551_ (.A(_0850_),
    .X(net390));
 sky130_fd_sc_hd__and2_1 _2552_ (.A(_0389_),
    .B(_0836_),
    .X(_0851_));
 sky130_fd_sc_hd__buf_1 _2553_ (.A(_0851_),
    .X(net391));
 sky130_fd_sc_hd__and2_1 _2554_ (.A(_0502_),
    .B(_0836_),
    .X(_0852_));
 sky130_fd_sc_hd__buf_1 _2555_ (.A(_0852_),
    .X(net392));
 sky130_fd_sc_hd__and2_1 _2556_ (.A(_0612_),
    .B(_0834_),
    .X(_0853_));
 sky130_fd_sc_hd__buf_1 _2557_ (.A(_0853_),
    .X(net393));
 sky130_fd_sc_hd__and2_1 _2558_ (.A(_0653_),
    .B(_0834_),
    .X(_0854_));
 sky130_fd_sc_hd__buf_1 _2559_ (.A(_0854_),
    .X(net394));
 sky130_fd_sc_hd__and2_1 _2560_ (.A(_0657_),
    .B(_0834_),
    .X(_0855_));
 sky130_fd_sc_hd__buf_1 _2561_ (.A(_0855_),
    .X(net395));
 sky130_fd_sc_hd__and2_1 _2562_ (.A(_0661_),
    .B(_0834_),
    .X(_0856_));
 sky130_fd_sc_hd__buf_1 _2563_ (.A(_0856_),
    .X(net396));
 sky130_fd_sc_hd__nor2_1 _2564_ (.A(_0835_),
    .B(_0666_),
    .Y(net397));
 sky130_fd_sc_hd__nor2_1 _2565_ (.A(_0835_),
    .B(_0670_),
    .Y(net398));
 sky130_fd_sc_hd__nor2_1 _2566_ (.A(_0835_),
    .B(_0674_),
    .Y(net400));
 sky130_fd_sc_hd__nor2_1 _2567_ (.A(_0835_),
    .B(_0678_),
    .Y(net401));
 sky130_fd_sc_hd__nor2_1 _2568_ (.A(_0835_),
    .B(net733),
    .Y(net402));
 sky130_fd_sc_hd__nor2_1 _2569_ (.A(_0835_),
    .B(net732),
    .Y(net403));
 sky130_fd_sc_hd__nor2_2 _2570_ (.A(_0835_),
    .B(_0689_),
    .Y(net404));
 sky130_fd_sc_hd__nor2_1 _2571_ (.A(_0835_),
    .B(net731),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _2572_ (.A(net744),
    .Y(_0857_));
 sky130_fd_sc_hd__a22o_2 _2573_ (.A1(_0998_),
    .A2(_1083_),
    .B1(_1079_),
    .B2(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__inv_2 _2574_ (.A(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__buf_4 _2575_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _2576_ (.A(_0860_),
    .B(_1100_),
    .Y(net502));
 sky130_fd_sc_hd__clkbuf_8 _2577_ (.A(_0859_),
    .X(_0861_));
 sky130_fd_sc_hd__nor2_2 _2578_ (.A(_1117_),
    .B(_0861_),
    .Y(net613));
 sky130_fd_sc_hd__nor2_2 _2579_ (.A(_0721_),
    .B(_0861_),
    .Y(net652));
 sky130_fd_sc_hd__nor2_2 _2580_ (.A(_0773_),
    .B(_0861_),
    .Y(net663));
 sky130_fd_sc_hd__nor2_2 _2581_ (.A(_0723_),
    .B(_0861_),
    .Y(net674));
 sky130_fd_sc_hd__nor2_1 _2582_ (.A(_0860_),
    .B(_0022_),
    .Y(net685));
 sky130_fd_sc_hd__nor2_2 _2583_ (.A(_0032_),
    .B(_0861_),
    .Y(net696));
 sky130_fd_sc_hd__nor2_2 _2584_ (.A(_0782_),
    .B(_0861_),
    .Y(net707));
 sky130_fd_sc_hd__nor2_2 _2585_ (.A(_0071_),
    .B(_0861_),
    .Y(net718));
 sky130_fd_sc_hd__nor2_2 _2586_ (.A(_0092_),
    .B(_0861_),
    .Y(net729));
 sky130_fd_sc_hd__nor2_1 _2587_ (.A(_0726_),
    .B(_0861_),
    .Y(net513));
 sky130_fd_sc_hd__nor2_2 _2588_ (.A(_1198_),
    .B(_0861_),
    .Y(net524));
 sky130_fd_sc_hd__buf_4 _2589_ (.A(_0859_),
    .X(_0862_));
 sky130_fd_sc_hd__nor2_1 _2590_ (.A(_0862_),
    .B(_0139_),
    .Y(net535));
 sky130_fd_sc_hd__nor2_1 _2591_ (.A(_0862_),
    .B(_0146_),
    .Y(net546));
 sky130_fd_sc_hd__nor2_1 _2592_ (.A(_0862_),
    .B(_0058_),
    .Y(net557));
 sky130_fd_sc_hd__nor2_1 _2593_ (.A(_0862_),
    .B(_0729_),
    .Y(net568));
 sky130_fd_sc_hd__nor2_1 _2594_ (.A(_0862_),
    .B(_0730_),
    .Y(net579));
 sky130_fd_sc_hd__nor2_1 _2595_ (.A(_0862_),
    .B(_0731_),
    .Y(net590));
 sky130_fd_sc_hd__nor2_1 _2596_ (.A(_0862_),
    .B(_0188_),
    .Y(net601));
 sky130_fd_sc_hd__nor2_2 _2597_ (.A(_0197_),
    .B(_0861_),
    .Y(net612));
 sky130_fd_sc_hd__nor2_2 _2598_ (.A(_0732_),
    .B(_0861_),
    .Y(net624));
 sky130_fd_sc_hd__nor2_2 _2599_ (.A(_0219_),
    .B(_0861_),
    .Y(net635));
 sky130_fd_sc_hd__nor2_1 _2600_ (.A(_0796_),
    .B(_0861_),
    .Y(net644));
 sky130_fd_sc_hd__nor2_1 _2601_ (.A(_0862_),
    .B(_0734_),
    .Y(net645));
 sky130_fd_sc_hd__nor2_1 _2602_ (.A(_0862_),
    .B(_0299_),
    .Y(net646));
 sky130_fd_sc_hd__nor2_1 _2603_ (.A(_0312_),
    .B(_0861_),
    .Y(net647));
 sky130_fd_sc_hd__nor2_1 _2604_ (.A(_0735_),
    .B(_0861_),
    .Y(net648));
 sky130_fd_sc_hd__nor2_1 _2605_ (.A(_0368_),
    .B(_0860_),
    .Y(net649));
 sky130_fd_sc_hd__and2_1 _2606_ (.A(_0858_),
    .B(_0232_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_2 _2607_ (.A(_0863_),
    .X(net650));
 sky130_fd_sc_hd__nor2_1 _2608_ (.A(_0381_),
    .B(_0860_),
    .Y(net651));
 sky130_fd_sc_hd__nor2_1 _2609_ (.A(_0391_),
    .B(_0860_),
    .Y(net653));
 sky130_fd_sc_hd__and2_1 _2610_ (.A(_0858_),
    .B(_0398_),
    .X(_0864_));
 sky130_fd_sc_hd__clkbuf_2 _2611_ (.A(_0864_),
    .X(net654));
 sky130_fd_sc_hd__and2_1 _2612_ (.A(_0858_),
    .B(_0363_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_2 _2613_ (.A(_0865_),
    .X(net655));
 sky130_fd_sc_hd__nor2_1 _2614_ (.A(_0807_),
    .B(_0860_),
    .Y(net656));
 sky130_fd_sc_hd__nor2_1 _2615_ (.A(_0737_),
    .B(_0860_),
    .Y(net657));
 sky130_fd_sc_hd__nor2_1 _2616_ (.A(_0862_),
    .B(_0472_),
    .Y(net658));
 sky130_fd_sc_hd__and2_1 _2617_ (.A(_0476_),
    .B(_0858_),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_2 _2618_ (.A(_0866_),
    .X(net659));
 sky130_fd_sc_hd__nor2_1 _2619_ (.A(_0862_),
    .B(_0484_),
    .Y(net660));
 sky130_fd_sc_hd__nor2_1 _2620_ (.A(_0490_),
    .B(_0860_),
    .Y(net661));
 sky130_fd_sc_hd__nor2_1 _2621_ (.A(_0862_),
    .B(_0494_),
    .Y(net662));
 sky130_fd_sc_hd__and2_1 _2622_ (.A(_0858_),
    .B(_0422_),
    .X(_0867_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2623_ (.A(_0867_),
    .X(net664));
 sky130_fd_sc_hd__nor2_1 _2624_ (.A(_0813_),
    .B(_0860_),
    .Y(net665));
 sky130_fd_sc_hd__nor2_1 _2625_ (.A(_0739_),
    .B(_0860_),
    .Y(net666));
 sky130_fd_sc_hd__nor2_1 _2626_ (.A(_0543_),
    .B(_0860_),
    .Y(net667));
 sky130_fd_sc_hd__and2_1 _2627_ (.A(_0858_),
    .B(_0550_),
    .X(_0868_));
 sky130_fd_sc_hd__clkbuf_2 _2628_ (.A(_0868_),
    .X(net668));
 sky130_fd_sc_hd__nor2_1 _2629_ (.A(_0571_),
    .B(_0860_),
    .Y(net669));
 sky130_fd_sc_hd__nor2_1 _2630_ (.A(_0741_),
    .B(_0860_),
    .Y(net670));
 sky130_fd_sc_hd__nor2_1 _2631_ (.A(_0862_),
    .B(_0595_),
    .Y(net671));
 sky130_fd_sc_hd__nor2_1 _2632_ (.A(_0596_),
    .B(_0860_),
    .Y(net672));
 sky130_fd_sc_hd__and2_1 _2633_ (.A(_0858_),
    .B(_0520_),
    .X(_0869_));
 sky130_fd_sc_hd__clkbuf_2 _2634_ (.A(_0869_),
    .X(net673));
 sky130_fd_sc_hd__nor2_1 _2635_ (.A(_0862_),
    .B(_0744_),
    .Y(net675));
 sky130_fd_sc_hd__nor2_1 _2636_ (.A(_0862_),
    .B(_0745_),
    .Y(net676));
 sky130_fd_sc_hd__nor2_1 _2637_ (.A(_0862_),
    .B(_0746_),
    .Y(net677));
 sky130_fd_sc_hd__nor2_1 _2638_ (.A(_0859_),
    .B(_0637_),
    .Y(net678));
 sky130_fd_sc_hd__nor2_1 _2639_ (.A(_0859_),
    .B(_0748_),
    .Y(net679));
 sky130_fd_sc_hd__nor2_1 _2640_ (.A(_0650_),
    .B(_0860_),
    .Y(net680));
 sky130_fd_sc_hd__nor2_1 _2641_ (.A(_0606_),
    .B(_0860_),
    .Y(net681));
 sky130_fd_sc_hd__inv_2 _2642_ (.A(net753),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_1 _2643_ (.A(_0870_),
    .B(net268),
    .Y(_0871_));
 sky130_fd_sc_hd__nand2_1 _2644_ (.A(_0871_),
    .B(_1010_),
    .Y(_0872_));
 sky130_fd_sc_hd__inv_2 _2645_ (.A(net756),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _2646_ (.A(_0873_),
    .B(net231),
    .Y(_0874_));
 sky130_fd_sc_hd__inv_2 _2647_ (.A(net762),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _2648_ (.A(_0875_),
    .B(net328),
    .Y(_0876_));
 sky130_fd_sc_hd__a21bo_1 _2649_ (.A1(_0872_),
    .A2(_0874_),
    .B1_N(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _2650_ (.A(_0857_),
    .B(net291),
    .Y(_0878_));
 sky130_fd_sc_hd__nand2_1 _2651_ (.A(_0877_),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nand2_1 _2652_ (.A(_1080_),
    .B(_1102_),
    .Y(_0880_));
 sky130_fd_sc_hd__o21ai_1 _2653_ (.A1(_1080_),
    .A2(_0879_),
    .B1(_0880_),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2_1 _2654_ (.A(_0871_),
    .B(_0874_),
    .Y(_0881_));
 sky130_fd_sc_hd__inv_2 _2655_ (.A(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand2_1 _2656_ (.A(_0882_),
    .B(_0989_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand2_1 _2657_ (.A(_0878_),
    .B(_0876_),
    .Y(_0884_));
 sky130_fd_sc_hd__inv_2 _2658_ (.A(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__nand2_1 _2659_ (.A(_0883_),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__inv_2 _2660_ (.A(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(_0887_),
    .A1(_1013_),
    .S(_1080_),
    .X(_0888_));
 sky130_fd_sc_hd__clkbuf_1 _2662_ (.A(_0888_),
    .X(_0001_));
 sky130_fd_sc_hd__nor3_1 _2663_ (.A(_1083_),
    .B(_0881_),
    .C(_0884_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_1 _2664_ (.A(_0889_),
    .B(net759),
    .Y(_0890_));
 sky130_fd_sc_hd__inv_2 _2665_ (.A(net738),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_1 _2666_ (.A(_0891_),
    .B(net176),
    .Y(_0892_));
 sky130_fd_sc_hd__inv_2 _2667_ (.A(net750),
    .Y(_0893_));
 sky130_fd_sc_hd__nand2_1 _2668_ (.A(_0893_),
    .B(net11),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_1 _2669_ (.A(_0892_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__inv_2 _2670_ (.A(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__inv_2 _2671_ (.A(net747),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2_1 _2672_ (.A(_0897_),
    .B(net74),
    .Y(_0898_));
 sky130_fd_sc_hd__inv_2 _2673_ (.A(net741),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _2674_ (.A(_0899_),
    .B(net138),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_1 _2675_ (.A(_0898_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__inv_2 _2676_ (.A(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__nand2_1 _2677_ (.A(_0896_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__o21ai_1 _2678_ (.A1(_1083_),
    .A2(_0903_),
    .B1(_1078_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor2_2 _2679_ (.A(net759),
    .B(_0980_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand3_2 _2680_ (.A(_0689_),
    .B(_0632_),
    .C(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__o21ai_2 _2681_ (.A1(_0685_),
    .A2(_0688_),
    .B1(_0905_),
    .Y(_0907_));
 sky130_fd_sc_hd__nand2_1 _2682_ (.A(_0906_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21oi_1 _2683_ (.A1(net760),
    .A2(_0904_),
    .B1(_0908_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _2684_ (.A(_0905_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21oi_1 _2685_ (.A1(_1080_),
    .A2(_0909_),
    .B1(_0889_),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_1 _2686_ (.A(_1078_),
    .B(_0981_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2_1 _2687_ (.A(_0900_),
    .B(_1120_),
    .Y(_0911_));
 sky130_fd_sc_hd__a21bo_1 _2688_ (.A1(_0911_),
    .A2(_0898_),
    .B1_N(_0894_),
    .X(_0912_));
 sky130_fd_sc_hd__nand2_1 _2689_ (.A(_0912_),
    .B(_0892_),
    .Y(_0913_));
 sky130_fd_sc_hd__nand2_1 _2690_ (.A(_0910_),
    .B(_1122_),
    .Y(_0914_));
 sky130_fd_sc_hd__o21ai_1 _2691_ (.A1(_0910_),
    .A2(_0913_),
    .B1(net766),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_1 _2692_ (.A(_0902_),
    .B(_1108_),
    .Y(_0915_));
 sky130_fd_sc_hd__nand2_1 _2693_ (.A(_0915_),
    .B(_0896_),
    .Y(_0916_));
 sky130_fd_sc_hd__inv_2 _2694_ (.A(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__mux2_1 _2695_ (.A0(_0917_),
    .A1(_1114_),
    .S(_0910_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_1 _2696_ (.A(_0918_),
    .X(_0005_));
 sky130_fd_sc_hd__nand2_1 _2697_ (.A(_0879_),
    .B(_0886_),
    .Y(_0919_));
 sky130_fd_sc_hd__nand2_1 _2698_ (.A(_0919_),
    .B(_0857_),
    .Y(_0920_));
 sky130_fd_sc_hd__buf_4 _2699_ (.A(_0909_),
    .X(_0921_));
 sky130_fd_sc_hd__nand2_1 _2700_ (.A(_0920_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__or3_1 _2701_ (.A(_0857_),
    .B(_0998_),
    .C(_0921_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _2702_ (.A(_0922_),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__nand3_2 _2703_ (.A(_0906_),
    .B(_0907_),
    .C(_0003_),
    .Y(_0925_));
 sky130_fd_sc_hd__inv_2 _2704_ (.A(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__nand2_1 _2705_ (.A(_0924_),
    .B(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__nand2_1 _2706_ (.A(_0925_),
    .B(net744),
    .Y(_0928_));
 sky130_fd_sc_hd__nand2_1 _2707_ (.A(_0927_),
    .B(net745),
    .Y(_0006_));
 sky130_fd_sc_hd__nand2_1 _2708_ (.A(_1020_),
    .B(net762),
    .Y(_0929_));
 sky130_fd_sc_hd__nand3_1 _2709_ (.A(_0877_),
    .B(_0886_),
    .C(_0878_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_1 _2710_ (.A(_0930_),
    .B(_0875_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _2711_ (.A(_0931_),
    .B(_0921_),
    .Y(_0932_));
 sky130_fd_sc_hd__o21ai_1 _2712_ (.A1(_0921_),
    .A2(_0929_),
    .B1(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_1 _2713_ (.A(_0933_),
    .B(_0926_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _2714_ (.A(_0925_),
    .B(net762),
    .Y(_0935_));
 sky130_fd_sc_hd__nand2_1 _2715_ (.A(_0934_),
    .B(net763),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_1 _2716_ (.A(_0879_),
    .B(_0887_),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2_1 _2717_ (.A(_0936_),
    .B(_0873_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _2718_ (.A(_0937_),
    .B(_0921_),
    .Y(_0938_));
 sky130_fd_sc_hd__or3_1 _2719_ (.A(_0873_),
    .B(_1002_),
    .C(_0921_),
    .X(_0939_));
 sky130_fd_sc_hd__nand2_1 _2720_ (.A(_0938_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand2_1 _2721_ (.A(_0940_),
    .B(_0926_),
    .Y(_0941_));
 sky130_fd_sc_hd__nand2_1 _2722_ (.A(_0925_),
    .B(net756),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _2723_ (.A(_0941_),
    .B(net757),
    .Y(_0008_));
 sky130_fd_sc_hd__nand3_1 _2724_ (.A(_0887_),
    .B(_0878_),
    .C(_0877_),
    .Y(_0943_));
 sky130_fd_sc_hd__nand2_1 _2725_ (.A(_0943_),
    .B(_0870_),
    .Y(_0944_));
 sky130_fd_sc_hd__nand2_1 _2726_ (.A(_0944_),
    .B(_0921_),
    .Y(_0945_));
 sky130_fd_sc_hd__or3_1 _2727_ (.A(_0870_),
    .B(_0996_),
    .C(_0921_),
    .X(_0946_));
 sky130_fd_sc_hd__nand2_1 _2728_ (.A(_0945_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _2729_ (.A(_0947_),
    .B(_0926_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand2_1 _2730_ (.A(_0925_),
    .B(net753),
    .Y(_0949_));
 sky130_fd_sc_hd__nand2_1 _2731_ (.A(_0948_),
    .B(net754),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_1 _2732_ (.A(_0913_),
    .B(_0916_),
    .Y(_0950_));
 sky130_fd_sc_hd__nand2_1 _2733_ (.A(_0950_),
    .B(_0891_),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _2734_ (.A(_0951_),
    .B(_0921_),
    .Y(_0952_));
 sky130_fd_sc_hd__or3_1 _2735_ (.A(_0891_),
    .B(_1094_),
    .C(_0921_),
    .X(_0953_));
 sky130_fd_sc_hd__nand2_1 _2736_ (.A(_0952_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__nor2_1 _2737_ (.A(_0904_),
    .B(_0908_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _2738_ (.A(_0954_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__nand3b_2 _2739_ (.A_N(_0904_),
    .B(_0906_),
    .C(_0907_),
    .Y(_0957_));
 sky130_fd_sc_hd__nand2_1 _2740_ (.A(_0957_),
    .B(net738),
    .Y(_0958_));
 sky130_fd_sc_hd__nand2_1 _2741_ (.A(_0956_),
    .B(net739),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _2742_ (.A(_0122_),
    .B(net750),
    .Y(_0959_));
 sky130_fd_sc_hd__nand3_1 _2743_ (.A(_0912_),
    .B(_0916_),
    .C(_0892_),
    .Y(_0960_));
 sky130_fd_sc_hd__nand2_1 _2744_ (.A(_0960_),
    .B(_0893_),
    .Y(_0961_));
 sky130_fd_sc_hd__nand2_1 _2745_ (.A(_0961_),
    .B(_0921_),
    .Y(_0962_));
 sky130_fd_sc_hd__o21ai_1 _2746_ (.A1(_0921_),
    .A2(_0959_),
    .B1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__nand2_1 _2747_ (.A(_0963_),
    .B(_0955_),
    .Y(_0964_));
 sky130_fd_sc_hd__nand2_1 _2748_ (.A(_0957_),
    .B(net750),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _2749_ (.A(_0964_),
    .B(net751),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2_1 _2750_ (.A(_0913_),
    .B(_0917_),
    .Y(_0966_));
 sky130_fd_sc_hd__nand2_1 _2751_ (.A(_0966_),
    .B(_0897_),
    .Y(_0967_));
 sky130_fd_sc_hd__nand2_1 _2752_ (.A(_0967_),
    .B(_0921_),
    .Y(_0968_));
 sky130_fd_sc_hd__or3_1 _2753_ (.A(_0897_),
    .B(_1092_),
    .C(_0921_),
    .X(_0969_));
 sky130_fd_sc_hd__nand2_1 _2754_ (.A(_0968_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__nand2_1 _2755_ (.A(_0970_),
    .B(_0955_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand2_1 _2756_ (.A(_0957_),
    .B(net747),
    .Y(_0972_));
 sky130_fd_sc_hd__nand2_1 _2757_ (.A(_0971_),
    .B(net748),
    .Y(_0012_));
 sky130_fd_sc_hd__nand3_1 _2758_ (.A(_0917_),
    .B(_0892_),
    .C(_0912_),
    .Y(_0973_));
 sky130_fd_sc_hd__nand2_1 _2759_ (.A(_0973_),
    .B(_0899_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_1 _2760_ (.A(_0974_),
    .B(_0921_),
    .Y(_0975_));
 sky130_fd_sc_hd__or3_1 _2761_ (.A(_0899_),
    .B(_1089_),
    .C(_0921_),
    .X(_0976_));
 sky130_fd_sc_hd__nand2_1 _2762_ (.A(_0975_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__nand2_1 _2763_ (.A(_0955_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__nand2_1 _2764_ (.A(_0957_),
    .B(net741),
    .Y(_0979_));
 sky130_fd_sc_hd__nand2_1 _2765_ (.A(_0978_),
    .B(net742),
    .Y(_0013_));
 sky130_fd_sc_hd__dfrtp_1 _2766_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_0000_),
    .RESET_B(net229),
    .Q(\arbiter.slave_sel[0][0] ));
 sky130_fd_sc_hd__dfrtp_4 _2767_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_0001_),
    .RESET_B(net229),
    .Q(\arbiter.slave_sel[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _2768_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(net761),
    .RESET_B(net229),
    .Q(\arbiter.state[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _2769_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(_0003_),
    .RESET_B(net229),
    .Q(\arbiter.state[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _2770_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(net767),
    .RESET_B(net229),
    .Q(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _2771_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(_0005_),
    .RESET_B(net229),
    .Q(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _2772_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(net746),
    .RESET_B(net229),
    .Q(\arbiter.slave_handled[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2773_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(net764),
    .RESET_B(net229),
    .Q(\arbiter.slave_handled[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2774_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(net758),
    .RESET_B(net229),
    .Q(\arbiter.slave_handled[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2775_ (.CLK(clknet_1_0__leaf_clk_i),
    .D(net755),
    .RESET_B(net229),
    .Q(\arbiter.slave_handled[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2776_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(net740),
    .RESET_B(net229),
    .Q(\arbiter.master_handled[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2777_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(net752),
    .RESET_B(net229),
    .Q(\arbiter.master_handled[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2778_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(net749),
    .RESET_B(net229),
    .Q(\arbiter.master_handled[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2779_ (.CLK(clknet_1_1__leaf_clk_i),
    .D(net743),
    .RESET_B(net229),
    .Q(\arbiter.master_handled[3] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_1__leaf_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\arbiter.master_handled[0] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\arbiter.master_handled[2] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0972_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0012_),
    .X(net749));
 sky130_fd_sc_hd__buf_1 hold13 (.A(\arbiter.master_handled[1] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0965_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0011_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\arbiter.slave_handled[3] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0949_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0009_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\arbiter.slave_handled[2] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0958_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0942_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0008_),
    .X(net758));
 sky130_fd_sc_hd__buf_1 hold22 (.A(\arbiter.state[0][0] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0890_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0002_),
    .X(net761));
 sky130_fd_sc_hd__buf_1 hold25 (.A(\arbiter.slave_handled[1] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0935_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0007_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\arbiter.master_sel[0][0] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0914_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0010_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0004_),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_2 hold31 (.A(\arbiter.state[0][1] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\arbiter.master_sel[0][1] ),
    .X(net769));
 sky130_fd_sc_hd__buf_1 hold33 (.A(\arbiter.slave_sel[0][1] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\arbiter.master_handled[3] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0979_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0013_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\arbiter.slave_handled[0] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0928_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0006_),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(mports_i[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(mports_i[108]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(mports_i[18]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(mports_i[190]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(mports_i[191]),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 input103 (.A(mports_i[192]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(mports_i[193]),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 input105 (.A(mports_i[194]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(mports_i[195]),
    .X(net106));
 sky130_fd_sc_hd__dlymetal6s2s_1 input107 (.A(mports_i[196]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(mports_i[197]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(mports_i[198]),
    .X(net109));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(mports_i[109]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input110 (.A(mports_i[199]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(mports_i[19]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(mports_i[1]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(mports_i[200]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(mports_i[201]),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(mports_i[202]),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(mports_i[203]),
    .X(net116));
 sky130_fd_sc_hd__buf_1 input117 (.A(mports_i[204]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(mports_i[205]),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 input119 (.A(mports_i[206]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(mports_i[10]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input120 (.A(mports_i[207]),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s2s_1 input121 (.A(mports_i[208]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(mports_i[209]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(mports_i[20]),
    .X(net123));
 sky130_fd_sc_hd__dlymetal6s2s_1 input124 (.A(mports_i[210]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(mports_i[211]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(mports_i[212]),
    .X(net126));
 sky130_fd_sc_hd__dlymetal6s2s_1 input127 (.A(mports_i[213]),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input128 (.A(mports_i[214]),
    .X(net128));
 sky130_fd_sc_hd__buf_1 input129 (.A(mports_i[215]),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input13 (.A(mports_i[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input130 (.A(mports_i[216]),
    .X(net130));
 sky130_fd_sc_hd__buf_1 input131 (.A(mports_i[217]),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 input132 (.A(mports_i[218]),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 input133 (.A(mports_i[219]),
    .X(net133));
 sky130_fd_sc_hd__buf_1 input134 (.A(mports_i[21]),
    .X(net134));
 sky130_fd_sc_hd__buf_1 input135 (.A(mports_i[220]),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input136 (.A(mports_i[221]),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 input137 (.A(mports_i[222]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(mports_i[223]),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 input139 (.A(mports_i[224]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input14 (.A(mports_i[111]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input140 (.A(mports_i[225]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(mports_i[226]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(mports_i[227]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(mports_i[22]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(mports_i[23]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(mports_i[24]),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(mports_i[25]),
    .X(net146));
 sky130_fd_sc_hd__buf_1 input147 (.A(mports_i[26]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(mports_i[27]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(mports_i[28]),
    .X(net149));
 sky130_fd_sc_hd__buf_1 input15 (.A(mports_i[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input150 (.A(mports_i[29]),
    .X(net150));
 sky130_fd_sc_hd__buf_1 input151 (.A(mports_i[2]),
    .X(net151));
 sky130_fd_sc_hd__buf_1 input152 (.A(mports_i[30]),
    .X(net152));
 sky130_fd_sc_hd__buf_1 input153 (.A(mports_i[31]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(mports_i[32]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(mports_i[33]),
    .X(net155));
 sky130_fd_sc_hd__buf_1 input156 (.A(mports_i[34]),
    .X(net156));
 sky130_fd_sc_hd__buf_1 input157 (.A(mports_i[35]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(mports_i[36]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(mports_i[37]),
    .X(net159));
 sky130_fd_sc_hd__buf_1 input16 (.A(mports_i[113]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(mports_i[38]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(mports_i[39]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(mports_i[3]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 input163 (.A(mports_i[40]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(mports_i[41]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 input165 (.A(mports_i[42]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(mports_i[43]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(mports_i[44]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(mports_i[45]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(mports_i[46]),
    .X(net169));
 sky130_fd_sc_hd__buf_1 input17 (.A(mports_i[114]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(mports_i[47]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(mports_i[48]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(mports_i[49]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(mports_i[4]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(mports_i[50]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(mports_i[51]),
    .X(net175));
 sky130_fd_sc_hd__buf_1 input176 (.A(mports_i[52]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(mports_i[53]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(mports_i[54]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(mports_i[55]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(mports_i[115]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(mports_i[56]),
    .X(net180));
 sky130_fd_sc_hd__buf_1 input181 (.A(mports_i[57]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(mports_i[58]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(mports_i[59]),
    .X(net183));
 sky130_fd_sc_hd__buf_1 input184 (.A(mports_i[5]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(mports_i[60]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(mports_i[61]),
    .X(net186));
 sky130_fd_sc_hd__buf_1 input187 (.A(mports_i[62]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(mports_i[63]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(mports_i[64]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(mports_i[116]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(mports_i[65]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(mports_i[66]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(mports_i[67]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(mports_i[68]),
    .X(net193));
 sky130_fd_sc_hd__buf_1 input194 (.A(mports_i[69]),
    .X(net194));
 sky130_fd_sc_hd__buf_1 input195 (.A(mports_i[6]),
    .X(net195));
 sky130_fd_sc_hd__buf_1 input196 (.A(mports_i[70]),
    .X(net196));
 sky130_fd_sc_hd__buf_1 input197 (.A(mports_i[71]),
    .X(net197));
 sky130_fd_sc_hd__buf_1 input198 (.A(mports_i[72]),
    .X(net198));
 sky130_fd_sc_hd__buf_1 input199 (.A(mports_i[73]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(mports_i[100]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(mports_i[117]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input200 (.A(mports_i[74]),
    .X(net200));
 sky130_fd_sc_hd__buf_1 input201 (.A(mports_i[75]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(mports_i[76]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(mports_i[77]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(mports_i[78]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(mports_i[79]),
    .X(net205));
 sky130_fd_sc_hd__buf_1 input206 (.A(mports_i[7]),
    .X(net206));
 sky130_fd_sc_hd__buf_1 input207 (.A(mports_i[80]),
    .X(net207));
 sky130_fd_sc_hd__buf_1 input208 (.A(mports_i[81]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(mports_i[82]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(mports_i[118]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(mports_i[83]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(mports_i[84]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(mports_i[85]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(mports_i[86]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(mports_i[87]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(mports_i[88]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(mports_i[89]),
    .X(net216));
 sky130_fd_sc_hd__buf_1 input217 (.A(mports_i[8]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(mports_i[90]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(mports_i[91]),
    .X(net219));
 sky130_fd_sc_hd__buf_1 input22 (.A(mports_i[119]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input220 (.A(mports_i[92]),
    .X(net220));
 sky130_fd_sc_hd__buf_1 input221 (.A(mports_i[93]),
    .X(net221));
 sky130_fd_sc_hd__buf_1 input222 (.A(mports_i[94]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(mports_i[95]),
    .X(net223));
 sky130_fd_sc_hd__buf_1 input224 (.A(mports_i[96]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(mports_i[97]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(mports_i[98]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(mports_i[99]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(mports_i[9]),
    .X(net228));
 sky130_fd_sc_hd__buf_6 input229 (.A(nrst_i),
    .X(net229));
 sky130_fd_sc_hd__buf_1 input23 (.A(mports_i[11]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input230 (.A(sports_i[0]),
    .X(net230));
 sky130_fd_sc_hd__buf_2 input231 (.A(sports_i[100]),
    .X(net231));
 sky130_fd_sc_hd__buf_1 input232 (.A(sports_i[101]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(sports_i[102]),
    .X(net233));
 sky130_fd_sc_hd__buf_1 input234 (.A(sports_i[103]),
    .X(net234));
 sky130_fd_sc_hd__buf_1 input235 (.A(sports_i[104]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(sports_i[105]),
    .X(net236));
 sky130_fd_sc_hd__buf_1 input237 (.A(sports_i[106]),
    .X(net237));
 sky130_fd_sc_hd__buf_1 input238 (.A(sports_i[107]),
    .X(net238));
 sky130_fd_sc_hd__buf_1 input239 (.A(sports_i[108]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(mports_i[120]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input240 (.A(sports_i[109]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(sports_i[10]),
    .X(net241));
 sky130_fd_sc_hd__dlymetal6s2s_1 input242 (.A(sports_i[110]),
    .X(net242));
 sky130_fd_sc_hd__buf_1 input243 (.A(sports_i[111]),
    .X(net243));
 sky130_fd_sc_hd__dlymetal6s2s_1 input244 (.A(sports_i[112]),
    .X(net244));
 sky130_fd_sc_hd__buf_1 input245 (.A(sports_i[113]),
    .X(net245));
 sky130_fd_sc_hd__buf_1 input246 (.A(sports_i[114]),
    .X(net246));
 sky130_fd_sc_hd__buf_1 input247 (.A(sports_i[115]),
    .X(net247));
 sky130_fd_sc_hd__buf_1 input248 (.A(sports_i[116]),
    .X(net248));
 sky130_fd_sc_hd__buf_1 input249 (.A(sports_i[117]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(mports_i[121]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input250 (.A(sports_i[118]),
    .X(net250));
 sky130_fd_sc_hd__buf_1 input251 (.A(sports_i[119]),
    .X(net251));
 sky130_fd_sc_hd__buf_1 input252 (.A(sports_i[11]),
    .X(net252));
 sky130_fd_sc_hd__dlymetal6s2s_1 input253 (.A(sports_i[120]),
    .X(net253));
 sky130_fd_sc_hd__buf_1 input254 (.A(sports_i[121]),
    .X(net254));
 sky130_fd_sc_hd__dlymetal6s2s_1 input255 (.A(sports_i[122]),
    .X(net255));
 sky130_fd_sc_hd__dlymetal6s2s_1 input256 (.A(sports_i[123]),
    .X(net256));
 sky130_fd_sc_hd__buf_1 input257 (.A(sports_i[124]),
    .X(net257));
 sky130_fd_sc_hd__buf_1 input258 (.A(sports_i[125]),
    .X(net258));
 sky130_fd_sc_hd__buf_1 input259 (.A(sports_i[126]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(mports_i[122]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input260 (.A(sports_i[127]),
    .X(net260));
 sky130_fd_sc_hd__buf_1 input261 (.A(sports_i[128]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 input262 (.A(sports_i[129]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 input263 (.A(sports_i[12]),
    .X(net263));
 sky130_fd_sc_hd__buf_1 input264 (.A(sports_i[130]),
    .X(net264));
 sky130_fd_sc_hd__buf_1 input265 (.A(sports_i[131]),
    .X(net265));
 sky130_fd_sc_hd__buf_1 input266 (.A(sports_i[132]),
    .X(net266));
 sky130_fd_sc_hd__buf_1 input267 (.A(sports_i[133]),
    .X(net267));
 sky130_fd_sc_hd__buf_2 input268 (.A(sports_i[134]),
    .X(net268));
 sky130_fd_sc_hd__buf_1 input269 (.A(sports_i[135]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(mports_i[123]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input270 (.A(sports_i[13]),
    .X(net270));
 sky130_fd_sc_hd__buf_1 input271 (.A(sports_i[14]),
    .X(net271));
 sky130_fd_sc_hd__buf_1 input272 (.A(sports_i[15]),
    .X(net272));
 sky130_fd_sc_hd__buf_1 input273 (.A(sports_i[16]),
    .X(net273));
 sky130_fd_sc_hd__buf_1 input274 (.A(sports_i[17]),
    .X(net274));
 sky130_fd_sc_hd__buf_1 input275 (.A(sports_i[18]),
    .X(net275));
 sky130_fd_sc_hd__buf_1 input276 (.A(sports_i[19]),
    .X(net276));
 sky130_fd_sc_hd__buf_1 input277 (.A(sports_i[1]),
    .X(net277));
 sky130_fd_sc_hd__buf_1 input278 (.A(sports_i[20]),
    .X(net278));
 sky130_fd_sc_hd__buf_1 input279 (.A(sports_i[21]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(mports_i[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input280 (.A(sports_i[22]),
    .X(net280));
 sky130_fd_sc_hd__buf_1 input281 (.A(sports_i[23]),
    .X(net281));
 sky130_fd_sc_hd__buf_1 input282 (.A(sports_i[24]),
    .X(net282));
 sky130_fd_sc_hd__buf_1 input283 (.A(sports_i[25]),
    .X(net283));
 sky130_fd_sc_hd__buf_1 input284 (.A(sports_i[26]),
    .X(net284));
 sky130_fd_sc_hd__buf_1 input285 (.A(sports_i[27]),
    .X(net285));
 sky130_fd_sc_hd__buf_1 input286 (.A(sports_i[28]),
    .X(net286));
 sky130_fd_sc_hd__buf_1 input287 (.A(sports_i[29]),
    .X(net287));
 sky130_fd_sc_hd__buf_1 input288 (.A(sports_i[2]),
    .X(net288));
 sky130_fd_sc_hd__buf_1 input289 (.A(sports_i[30]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(mports_i[125]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input290 (.A(sports_i[31]),
    .X(net290));
 sky130_fd_sc_hd__buf_2 input291 (.A(sports_i[32]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 input292 (.A(sports_i[33]),
    .X(net292));
 sky130_fd_sc_hd__buf_1 input293 (.A(sports_i[34]),
    .X(net293));
 sky130_fd_sc_hd__buf_1 input294 (.A(sports_i[35]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 input295 (.A(sports_i[36]),
    .X(net295));
 sky130_fd_sc_hd__buf_1 input296 (.A(sports_i[37]),
    .X(net296));
 sky130_fd_sc_hd__buf_1 input297 (.A(sports_i[38]),
    .X(net297));
 sky130_fd_sc_hd__buf_1 input298 (.A(sports_i[39]),
    .X(net298));
 sky130_fd_sc_hd__buf_1 input299 (.A(sports_i[3]),
    .X(net299));
 sky130_fd_sc_hd__buf_1 input3 (.A(mports_i[101]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(mports_i[126]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input300 (.A(sports_i[40]),
    .X(net300));
 sky130_fd_sc_hd__buf_1 input301 (.A(sports_i[41]),
    .X(net301));
 sky130_fd_sc_hd__buf_1 input302 (.A(sports_i[42]),
    .X(net302));
 sky130_fd_sc_hd__buf_1 input303 (.A(sports_i[43]),
    .X(net303));
 sky130_fd_sc_hd__buf_1 input304 (.A(sports_i[44]),
    .X(net304));
 sky130_fd_sc_hd__buf_1 input305 (.A(sports_i[45]),
    .X(net305));
 sky130_fd_sc_hd__buf_1 input306 (.A(sports_i[46]),
    .X(net306));
 sky130_fd_sc_hd__buf_1 input307 (.A(sports_i[47]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 input308 (.A(sports_i[48]),
    .X(net308));
 sky130_fd_sc_hd__buf_1 input309 (.A(sports_i[49]),
    .X(net309));
 sky130_fd_sc_hd__buf_1 input31 (.A(mports_i[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input310 (.A(sports_i[4]),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 input311 (.A(sports_i[50]),
    .X(net311));
 sky130_fd_sc_hd__buf_1 input312 (.A(sports_i[51]),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 input313 (.A(sports_i[52]),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 input314 (.A(sports_i[53]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 input315 (.A(sports_i[54]),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 input316 (.A(sports_i[55]),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 input317 (.A(sports_i[56]),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 input318 (.A(sports_i[57]),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 input319 (.A(sports_i[58]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(mports_i[128]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input320 (.A(sports_i[59]),
    .X(net320));
 sky130_fd_sc_hd__buf_1 input321 (.A(sports_i[5]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 input322 (.A(sports_i[60]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 input323 (.A(sports_i[61]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 input324 (.A(sports_i[62]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 input325 (.A(sports_i[63]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 input326 (.A(sports_i[64]),
    .X(net326));
 sky130_fd_sc_hd__buf_1 input327 (.A(sports_i[65]),
    .X(net327));
 sky130_fd_sc_hd__buf_2 input328 (.A(sports_i[66]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 input329 (.A(sports_i[67]),
    .X(net329));
 sky130_fd_sc_hd__buf_1 input33 (.A(mports_i[129]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input330 (.A(sports_i[68]),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 input331 (.A(sports_i[69]),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 input332 (.A(sports_i[6]),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_1 input333 (.A(sports_i[70]),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 input334 (.A(sports_i[71]),
    .X(net334));
 sky130_fd_sc_hd__buf_1 input335 (.A(sports_i[72]),
    .X(net335));
 sky130_fd_sc_hd__buf_1 input336 (.A(sports_i[73]),
    .X(net336));
 sky130_fd_sc_hd__buf_1 input337 (.A(sports_i[74]),
    .X(net337));
 sky130_fd_sc_hd__buf_1 input338 (.A(sports_i[75]),
    .X(net338));
 sky130_fd_sc_hd__buf_1 input339 (.A(sports_i[76]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(mports_i[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input340 (.A(sports_i[77]),
    .X(net340));
 sky130_fd_sc_hd__buf_1 input341 (.A(sports_i[78]),
    .X(net341));
 sky130_fd_sc_hd__buf_1 input342 (.A(sports_i[79]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 input343 (.A(sports_i[7]),
    .X(net343));
 sky130_fd_sc_hd__buf_1 input344 (.A(sports_i[80]),
    .X(net344));
 sky130_fd_sc_hd__buf_1 input345 (.A(sports_i[81]),
    .X(net345));
 sky130_fd_sc_hd__buf_1 input346 (.A(sports_i[82]),
    .X(net346));
 sky130_fd_sc_hd__buf_1 input347 (.A(sports_i[83]),
    .X(net347));
 sky130_fd_sc_hd__buf_1 input348 (.A(sports_i[84]),
    .X(net348));
 sky130_fd_sc_hd__buf_1 input349 (.A(sports_i[85]),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(mports_i[130]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input350 (.A(sports_i[86]),
    .X(net350));
 sky130_fd_sc_hd__buf_1 input351 (.A(sports_i[87]),
    .X(net351));
 sky130_fd_sc_hd__buf_1 input352 (.A(sports_i[88]),
    .X(net352));
 sky130_fd_sc_hd__buf_1 input353 (.A(sports_i[89]),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 input354 (.A(sports_i[8]),
    .X(net354));
 sky130_fd_sc_hd__buf_1 input355 (.A(sports_i[90]),
    .X(net355));
 sky130_fd_sc_hd__buf_1 input356 (.A(sports_i[91]),
    .X(net356));
 sky130_fd_sc_hd__buf_1 input357 (.A(sports_i[92]),
    .X(net357));
 sky130_fd_sc_hd__buf_1 input358 (.A(sports_i[93]),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 input359 (.A(sports_i[94]),
    .X(net359));
 sky130_fd_sc_hd__buf_1 input36 (.A(mports_i[131]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input360 (.A(sports_i[95]),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 input361 (.A(sports_i[96]),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 input362 (.A(sports_i[97]),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 input363 (.A(sports_i[98]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 input364 (.A(sports_i[99]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 input365 (.A(sports_i[9]),
    .X(net365));
 sky130_fd_sc_hd__buf_1 input37 (.A(mports_i[132]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(mports_i[133]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(mports_i[134]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(mports_i[102]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(mports_i[135]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(mports_i[136]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(mports_i[137]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(mports_i[138]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(mports_i[139]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(mports_i[13]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(mports_i[140]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(mports_i[141]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(mports_i[142]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(mports_i[143]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(mports_i[103]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(mports_i[144]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(mports_i[145]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(mports_i[146]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(mports_i[147]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(mports_i[148]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(mports_i[149]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(mports_i[14]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(mports_i[150]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(mports_i[151]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(mports_i[152]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input6 (.A(mports_i[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input60 (.A(mports_i[153]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(mports_i[154]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(mports_i[155]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(mports_i[156]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(mports_i[157]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(mports_i[158]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(mports_i[159]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(mports_i[15]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(mports_i[160]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(mports_i[161]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(mports_i[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input70 (.A(mports_i[162]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(mports_i[163]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(mports_i[164]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(mports_i[165]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(mports_i[166]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(mports_i[167]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(mports_i[168]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(mports_i[169]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(mports_i[16]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(mports_i[170]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(mports_i[106]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input80 (.A(mports_i[171]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(mports_i[172]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(mports_i[173]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(mports_i[174]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(mports_i[175]),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 input85 (.A(mports_i[176]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(mports_i[177]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(mports_i[178]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(mports_i[179]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(mports_i[17]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(mports_i[107]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input90 (.A(mports_i[180]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(mports_i[181]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(mports_i[182]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(mports_i[183]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(mports_i[184]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(mports_i[185]),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 input96 (.A(mports_i[186]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(mports_i[187]),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 input98 (.A(mports_i[188]),
    .X(net98));
 sky130_fd_sc_hd__dlymetal6s2s_1 input99 (.A(mports_i[189]),
    .X(net99));
 sky130_fd_sc_hd__buf_12 output366 (.A(net366),
    .X(mports_o[0]));
 sky130_fd_sc_hd__buf_12 output367 (.A(net367),
    .X(mports_o[100]));
 sky130_fd_sc_hd__buf_12 output368 (.A(net368),
    .X(mports_o[101]));
 sky130_fd_sc_hd__buf_12 output369 (.A(net369),
    .X(mports_o[102]));
 sky130_fd_sc_hd__buf_12 output370 (.A(net370),
    .X(mports_o[103]));
 sky130_fd_sc_hd__buf_12 output371 (.A(net371),
    .X(mports_o[104]));
 sky130_fd_sc_hd__buf_12 output372 (.A(net372),
    .X(mports_o[105]));
 sky130_fd_sc_hd__buf_12 output373 (.A(net373),
    .X(mports_o[106]));
 sky130_fd_sc_hd__buf_12 output374 (.A(net374),
    .X(mports_o[107]));
 sky130_fd_sc_hd__buf_12 output375 (.A(net375),
    .X(mports_o[108]));
 sky130_fd_sc_hd__buf_12 output376 (.A(net376),
    .X(mports_o[109]));
 sky130_fd_sc_hd__buf_12 output377 (.A(net377),
    .X(mports_o[10]));
 sky130_fd_sc_hd__buf_12 output378 (.A(net378),
    .X(mports_o[110]));
 sky130_fd_sc_hd__buf_12 output379 (.A(net379),
    .X(mports_o[111]));
 sky130_fd_sc_hd__buf_12 output380 (.A(net380),
    .X(mports_o[112]));
 sky130_fd_sc_hd__buf_12 output381 (.A(net381),
    .X(mports_o[113]));
 sky130_fd_sc_hd__buf_12 output382 (.A(net382),
    .X(mports_o[114]));
 sky130_fd_sc_hd__buf_12 output383 (.A(net383),
    .X(mports_o[115]));
 sky130_fd_sc_hd__buf_12 output384 (.A(net384),
    .X(mports_o[116]));
 sky130_fd_sc_hd__buf_12 output385 (.A(net385),
    .X(mports_o[117]));
 sky130_fd_sc_hd__buf_12 output386 (.A(net386),
    .X(mports_o[118]));
 sky130_fd_sc_hd__buf_12 output387 (.A(net387),
    .X(mports_o[119]));
 sky130_fd_sc_hd__buf_12 output388 (.A(net388),
    .X(mports_o[11]));
 sky130_fd_sc_hd__buf_12 output389 (.A(net389),
    .X(mports_o[120]));
 sky130_fd_sc_hd__buf_12 output390 (.A(net390),
    .X(mports_o[121]));
 sky130_fd_sc_hd__buf_12 output391 (.A(net391),
    .X(mports_o[122]));
 sky130_fd_sc_hd__buf_12 output392 (.A(net392),
    .X(mports_o[123]));
 sky130_fd_sc_hd__buf_12 output393 (.A(net393),
    .X(mports_o[124]));
 sky130_fd_sc_hd__buf_12 output394 (.A(net394),
    .X(mports_o[125]));
 sky130_fd_sc_hd__buf_12 output395 (.A(net395),
    .X(mports_o[126]));
 sky130_fd_sc_hd__buf_12 output396 (.A(net396),
    .X(mports_o[127]));
 sky130_fd_sc_hd__buf_12 output397 (.A(net397),
    .X(mports_o[128]));
 sky130_fd_sc_hd__buf_12 output398 (.A(net398),
    .X(mports_o[129]));
 sky130_fd_sc_hd__buf_12 output399 (.A(net399),
    .X(mports_o[12]));
 sky130_fd_sc_hd__buf_12 output400 (.A(net400),
    .X(mports_o[130]));
 sky130_fd_sc_hd__buf_12 output401 (.A(net401),
    .X(mports_o[131]));
 sky130_fd_sc_hd__buf_12 output402 (.A(net402),
    .X(mports_o[132]));
 sky130_fd_sc_hd__buf_12 output403 (.A(net403),
    .X(mports_o[133]));
 sky130_fd_sc_hd__buf_12 output404 (.A(net404),
    .X(mports_o[134]));
 sky130_fd_sc_hd__buf_12 output405 (.A(net405),
    .X(mports_o[135]));
 sky130_fd_sc_hd__buf_12 output406 (.A(net406),
    .X(mports_o[13]));
 sky130_fd_sc_hd__buf_12 output407 (.A(net407),
    .X(mports_o[14]));
 sky130_fd_sc_hd__buf_12 output408 (.A(net408),
    .X(mports_o[15]));
 sky130_fd_sc_hd__buf_12 output409 (.A(net409),
    .X(mports_o[16]));
 sky130_fd_sc_hd__buf_12 output410 (.A(net410),
    .X(mports_o[17]));
 sky130_fd_sc_hd__buf_12 output411 (.A(net411),
    .X(mports_o[18]));
 sky130_fd_sc_hd__buf_12 output412 (.A(net412),
    .X(mports_o[19]));
 sky130_fd_sc_hd__buf_12 output413 (.A(net413),
    .X(mports_o[1]));
 sky130_fd_sc_hd__buf_12 output414 (.A(net414),
    .X(mports_o[20]));
 sky130_fd_sc_hd__buf_12 output415 (.A(net415),
    .X(mports_o[21]));
 sky130_fd_sc_hd__buf_12 output416 (.A(net416),
    .X(mports_o[22]));
 sky130_fd_sc_hd__buf_12 output417 (.A(net417),
    .X(mports_o[23]));
 sky130_fd_sc_hd__buf_12 output418 (.A(net418),
    .X(mports_o[24]));
 sky130_fd_sc_hd__buf_12 output419 (.A(net419),
    .X(mports_o[25]));
 sky130_fd_sc_hd__buf_12 output420 (.A(net420),
    .X(mports_o[26]));
 sky130_fd_sc_hd__buf_12 output421 (.A(net421),
    .X(mports_o[27]));
 sky130_fd_sc_hd__buf_12 output422 (.A(net422),
    .X(mports_o[28]));
 sky130_fd_sc_hd__buf_12 output423 (.A(net423),
    .X(mports_o[29]));
 sky130_fd_sc_hd__buf_12 output424 (.A(net424),
    .X(mports_o[2]));
 sky130_fd_sc_hd__buf_12 output425 (.A(net425),
    .X(mports_o[30]));
 sky130_fd_sc_hd__buf_12 output426 (.A(net426),
    .X(mports_o[31]));
 sky130_fd_sc_hd__buf_12 output427 (.A(net427),
    .X(mports_o[32]));
 sky130_fd_sc_hd__buf_12 output428 (.A(net428),
    .X(mports_o[33]));
 sky130_fd_sc_hd__buf_12 output429 (.A(net429),
    .X(mports_o[34]));
 sky130_fd_sc_hd__buf_12 output430 (.A(net430),
    .X(mports_o[35]));
 sky130_fd_sc_hd__buf_12 output431 (.A(net431),
    .X(mports_o[36]));
 sky130_fd_sc_hd__buf_12 output432 (.A(net432),
    .X(mports_o[37]));
 sky130_fd_sc_hd__buf_12 output433 (.A(net433),
    .X(mports_o[38]));
 sky130_fd_sc_hd__buf_12 output434 (.A(net434),
    .X(mports_o[39]));
 sky130_fd_sc_hd__buf_12 output435 (.A(net435),
    .X(mports_o[3]));
 sky130_fd_sc_hd__buf_12 output436 (.A(net436),
    .X(mports_o[40]));
 sky130_fd_sc_hd__buf_12 output437 (.A(net437),
    .X(mports_o[41]));
 sky130_fd_sc_hd__buf_12 output438 (.A(net438),
    .X(mports_o[42]));
 sky130_fd_sc_hd__buf_12 output439 (.A(net439),
    .X(mports_o[43]));
 sky130_fd_sc_hd__buf_12 output440 (.A(net440),
    .X(mports_o[44]));
 sky130_fd_sc_hd__buf_12 output441 (.A(net441),
    .X(mports_o[45]));
 sky130_fd_sc_hd__buf_12 output442 (.A(net442),
    .X(mports_o[46]));
 sky130_fd_sc_hd__buf_12 output443 (.A(net443),
    .X(mports_o[47]));
 sky130_fd_sc_hd__buf_12 output444 (.A(net444),
    .X(mports_o[48]));
 sky130_fd_sc_hd__buf_12 output445 (.A(net445),
    .X(mports_o[49]));
 sky130_fd_sc_hd__buf_12 output446 (.A(net446),
    .X(mports_o[4]));
 sky130_fd_sc_hd__buf_12 output447 (.A(net447),
    .X(mports_o[50]));
 sky130_fd_sc_hd__buf_12 output448 (.A(net448),
    .X(mports_o[51]));
 sky130_fd_sc_hd__buf_12 output449 (.A(net449),
    .X(mports_o[52]));
 sky130_fd_sc_hd__buf_12 output450 (.A(net450),
    .X(mports_o[53]));
 sky130_fd_sc_hd__buf_12 output451 (.A(net451),
    .X(mports_o[54]));
 sky130_fd_sc_hd__buf_12 output452 (.A(net452),
    .X(mports_o[55]));
 sky130_fd_sc_hd__buf_12 output453 (.A(net453),
    .X(mports_o[56]));
 sky130_fd_sc_hd__buf_12 output454 (.A(net454),
    .X(mports_o[57]));
 sky130_fd_sc_hd__buf_12 output455 (.A(net455),
    .X(mports_o[58]));
 sky130_fd_sc_hd__buf_12 output456 (.A(net456),
    .X(mports_o[59]));
 sky130_fd_sc_hd__buf_12 output457 (.A(net457),
    .X(mports_o[5]));
 sky130_fd_sc_hd__buf_12 output458 (.A(net458),
    .X(mports_o[60]));
 sky130_fd_sc_hd__buf_12 output459 (.A(net459),
    .X(mports_o[61]));
 sky130_fd_sc_hd__buf_12 output460 (.A(net460),
    .X(mports_o[62]));
 sky130_fd_sc_hd__buf_12 output461 (.A(net461),
    .X(mports_o[63]));
 sky130_fd_sc_hd__buf_12 output462 (.A(net462),
    .X(mports_o[64]));
 sky130_fd_sc_hd__buf_12 output463 (.A(net463),
    .X(mports_o[65]));
 sky130_fd_sc_hd__buf_12 output464 (.A(net464),
    .X(mports_o[66]));
 sky130_fd_sc_hd__buf_12 output465 (.A(net465),
    .X(mports_o[67]));
 sky130_fd_sc_hd__buf_12 output466 (.A(net466),
    .X(mports_o[68]));
 sky130_fd_sc_hd__buf_12 output467 (.A(net467),
    .X(mports_o[69]));
 sky130_fd_sc_hd__buf_12 output468 (.A(net468),
    .X(mports_o[6]));
 sky130_fd_sc_hd__buf_12 output469 (.A(net469),
    .X(mports_o[70]));
 sky130_fd_sc_hd__buf_12 output470 (.A(net470),
    .X(mports_o[71]));
 sky130_fd_sc_hd__buf_12 output471 (.A(net471),
    .X(mports_o[72]));
 sky130_fd_sc_hd__buf_12 output472 (.A(net472),
    .X(mports_o[73]));
 sky130_fd_sc_hd__buf_12 output473 (.A(net473),
    .X(mports_o[74]));
 sky130_fd_sc_hd__buf_12 output474 (.A(net474),
    .X(mports_o[75]));
 sky130_fd_sc_hd__buf_12 output475 (.A(net475),
    .X(mports_o[76]));
 sky130_fd_sc_hd__buf_12 output476 (.A(net476),
    .X(mports_o[77]));
 sky130_fd_sc_hd__buf_12 output477 (.A(net477),
    .X(mports_o[78]));
 sky130_fd_sc_hd__buf_12 output478 (.A(net478),
    .X(mports_o[79]));
 sky130_fd_sc_hd__buf_12 output479 (.A(net479),
    .X(mports_o[7]));
 sky130_fd_sc_hd__buf_12 output480 (.A(net480),
    .X(mports_o[80]));
 sky130_fd_sc_hd__buf_12 output481 (.A(net481),
    .X(mports_o[81]));
 sky130_fd_sc_hd__buf_12 output482 (.A(net482),
    .X(mports_o[82]));
 sky130_fd_sc_hd__buf_12 output483 (.A(net483),
    .X(mports_o[83]));
 sky130_fd_sc_hd__buf_12 output484 (.A(net484),
    .X(mports_o[84]));
 sky130_fd_sc_hd__buf_12 output485 (.A(net485),
    .X(mports_o[85]));
 sky130_fd_sc_hd__buf_12 output486 (.A(net486),
    .X(mports_o[86]));
 sky130_fd_sc_hd__buf_12 output487 (.A(net487),
    .X(mports_o[87]));
 sky130_fd_sc_hd__buf_12 output488 (.A(net488),
    .X(mports_o[88]));
 sky130_fd_sc_hd__buf_12 output489 (.A(net489),
    .X(mports_o[89]));
 sky130_fd_sc_hd__buf_12 output490 (.A(net490),
    .X(mports_o[8]));
 sky130_fd_sc_hd__buf_12 output491 (.A(net491),
    .X(mports_o[90]));
 sky130_fd_sc_hd__buf_12 output492 (.A(net492),
    .X(mports_o[91]));
 sky130_fd_sc_hd__buf_12 output493 (.A(net493),
    .X(mports_o[92]));
 sky130_fd_sc_hd__buf_12 output494 (.A(net494),
    .X(mports_o[93]));
 sky130_fd_sc_hd__buf_12 output495 (.A(net495),
    .X(mports_o[94]));
 sky130_fd_sc_hd__buf_12 output496 (.A(net496),
    .X(mports_o[95]));
 sky130_fd_sc_hd__buf_12 output497 (.A(net497),
    .X(mports_o[96]));
 sky130_fd_sc_hd__buf_12 output498 (.A(net498),
    .X(mports_o[97]));
 sky130_fd_sc_hd__buf_12 output499 (.A(net499),
    .X(mports_o[98]));
 sky130_fd_sc_hd__buf_12 output500 (.A(net500),
    .X(mports_o[99]));
 sky130_fd_sc_hd__buf_12 output501 (.A(net501),
    .X(mports_o[9]));
 sky130_fd_sc_hd__buf_12 output502 (.A(net502),
    .X(sports_o[0]));
 sky130_fd_sc_hd__buf_12 output503 (.A(net503),
    .X(sports_o[100]));
 sky130_fd_sc_hd__buf_12 output504 (.A(net504),
    .X(sports_o[101]));
 sky130_fd_sc_hd__buf_12 output505 (.A(net505),
    .X(sports_o[102]));
 sky130_fd_sc_hd__buf_12 output506 (.A(net506),
    .X(sports_o[103]));
 sky130_fd_sc_hd__buf_12 output507 (.A(net507),
    .X(sports_o[104]));
 sky130_fd_sc_hd__buf_12 output508 (.A(net508),
    .X(sports_o[105]));
 sky130_fd_sc_hd__buf_12 output509 (.A(net509),
    .X(sports_o[106]));
 sky130_fd_sc_hd__buf_12 output510 (.A(net510),
    .X(sports_o[107]));
 sky130_fd_sc_hd__buf_12 output511 (.A(net511),
    .X(sports_o[108]));
 sky130_fd_sc_hd__buf_12 output512 (.A(net512),
    .X(sports_o[109]));
 sky130_fd_sc_hd__buf_12 output513 (.A(net513),
    .X(sports_o[10]));
 sky130_fd_sc_hd__buf_12 output514 (.A(net514),
    .X(sports_o[110]));
 sky130_fd_sc_hd__buf_12 output515 (.A(net515),
    .X(sports_o[111]));
 sky130_fd_sc_hd__buf_12 output516 (.A(net516),
    .X(sports_o[112]));
 sky130_fd_sc_hd__buf_12 output517 (.A(net517),
    .X(sports_o[113]));
 sky130_fd_sc_hd__buf_12 output518 (.A(net518),
    .X(sports_o[114]));
 sky130_fd_sc_hd__buf_12 output519 (.A(net519),
    .X(sports_o[115]));
 sky130_fd_sc_hd__buf_12 output520 (.A(net520),
    .X(sports_o[116]));
 sky130_fd_sc_hd__buf_12 output521 (.A(net521),
    .X(sports_o[117]));
 sky130_fd_sc_hd__buf_12 output522 (.A(net522),
    .X(sports_o[118]));
 sky130_fd_sc_hd__buf_12 output523 (.A(net523),
    .X(sports_o[119]));
 sky130_fd_sc_hd__buf_12 output524 (.A(net524),
    .X(sports_o[11]));
 sky130_fd_sc_hd__buf_12 output525 (.A(net525),
    .X(sports_o[120]));
 sky130_fd_sc_hd__buf_12 output526 (.A(net526),
    .X(sports_o[121]));
 sky130_fd_sc_hd__buf_12 output527 (.A(net527),
    .X(sports_o[122]));
 sky130_fd_sc_hd__buf_12 output528 (.A(net528),
    .X(sports_o[123]));
 sky130_fd_sc_hd__buf_12 output529 (.A(net529),
    .X(sports_o[124]));
 sky130_fd_sc_hd__buf_12 output530 (.A(net530),
    .X(sports_o[125]));
 sky130_fd_sc_hd__buf_12 output531 (.A(net531),
    .X(sports_o[126]));
 sky130_fd_sc_hd__buf_12 output532 (.A(net532),
    .X(sports_o[127]));
 sky130_fd_sc_hd__buf_12 output533 (.A(net533),
    .X(sports_o[128]));
 sky130_fd_sc_hd__buf_12 output534 (.A(net534),
    .X(sports_o[129]));
 sky130_fd_sc_hd__buf_12 output535 (.A(net535),
    .X(sports_o[12]));
 sky130_fd_sc_hd__buf_12 output536 (.A(net536),
    .X(sports_o[130]));
 sky130_fd_sc_hd__buf_12 output537 (.A(net537),
    .X(sports_o[131]));
 sky130_fd_sc_hd__buf_12 output538 (.A(net538),
    .X(sports_o[132]));
 sky130_fd_sc_hd__buf_12 output539 (.A(net539),
    .X(sports_o[133]));
 sky130_fd_sc_hd__buf_12 output540 (.A(net540),
    .X(sports_o[134]));
 sky130_fd_sc_hd__buf_12 output541 (.A(net541),
    .X(sports_o[135]));
 sky130_fd_sc_hd__buf_12 output542 (.A(net542),
    .X(sports_o[136]));
 sky130_fd_sc_hd__buf_12 output543 (.A(net543),
    .X(sports_o[137]));
 sky130_fd_sc_hd__buf_12 output544 (.A(net544),
    .X(sports_o[138]));
 sky130_fd_sc_hd__buf_12 output545 (.A(net545),
    .X(sports_o[139]));
 sky130_fd_sc_hd__buf_12 output546 (.A(net546),
    .X(sports_o[13]));
 sky130_fd_sc_hd__buf_12 output547 (.A(net547),
    .X(sports_o[140]));
 sky130_fd_sc_hd__buf_12 output548 (.A(net548),
    .X(sports_o[141]));
 sky130_fd_sc_hd__buf_12 output549 (.A(net549),
    .X(sports_o[142]));
 sky130_fd_sc_hd__buf_12 output550 (.A(net550),
    .X(sports_o[143]));
 sky130_fd_sc_hd__buf_12 output551 (.A(net551),
    .X(sports_o[144]));
 sky130_fd_sc_hd__buf_12 output552 (.A(net552),
    .X(sports_o[145]));
 sky130_fd_sc_hd__buf_12 output553 (.A(net553),
    .X(sports_o[146]));
 sky130_fd_sc_hd__buf_12 output554 (.A(net554),
    .X(sports_o[147]));
 sky130_fd_sc_hd__buf_12 output555 (.A(net555),
    .X(sports_o[148]));
 sky130_fd_sc_hd__buf_12 output556 (.A(net556),
    .X(sports_o[149]));
 sky130_fd_sc_hd__buf_12 output557 (.A(net557),
    .X(sports_o[14]));
 sky130_fd_sc_hd__buf_12 output558 (.A(net558),
    .X(sports_o[150]));
 sky130_fd_sc_hd__buf_12 output559 (.A(net559),
    .X(sports_o[151]));
 sky130_fd_sc_hd__buf_12 output560 (.A(net560),
    .X(sports_o[152]));
 sky130_fd_sc_hd__buf_12 output561 (.A(net561),
    .X(sports_o[153]));
 sky130_fd_sc_hd__buf_12 output562 (.A(net562),
    .X(sports_o[154]));
 sky130_fd_sc_hd__buf_12 output563 (.A(net563),
    .X(sports_o[155]));
 sky130_fd_sc_hd__buf_12 output564 (.A(net564),
    .X(sports_o[156]));
 sky130_fd_sc_hd__buf_12 output565 (.A(net565),
    .X(sports_o[157]));
 sky130_fd_sc_hd__buf_12 output566 (.A(net566),
    .X(sports_o[158]));
 sky130_fd_sc_hd__buf_12 output567 (.A(net567),
    .X(sports_o[159]));
 sky130_fd_sc_hd__buf_12 output568 (.A(net568),
    .X(sports_o[15]));
 sky130_fd_sc_hd__buf_12 output569 (.A(net569),
    .X(sports_o[160]));
 sky130_fd_sc_hd__buf_12 output570 (.A(net570),
    .X(sports_o[161]));
 sky130_fd_sc_hd__buf_12 output571 (.A(net571),
    .X(sports_o[162]));
 sky130_fd_sc_hd__buf_12 output572 (.A(net572),
    .X(sports_o[163]));
 sky130_fd_sc_hd__buf_12 output573 (.A(net573),
    .X(sports_o[164]));
 sky130_fd_sc_hd__buf_12 output574 (.A(net574),
    .X(sports_o[165]));
 sky130_fd_sc_hd__buf_12 output575 (.A(net575),
    .X(sports_o[166]));
 sky130_fd_sc_hd__buf_12 output576 (.A(net576),
    .X(sports_o[167]));
 sky130_fd_sc_hd__buf_12 output577 (.A(net577),
    .X(sports_o[168]));
 sky130_fd_sc_hd__buf_12 output578 (.A(net578),
    .X(sports_o[169]));
 sky130_fd_sc_hd__buf_12 output579 (.A(net579),
    .X(sports_o[16]));
 sky130_fd_sc_hd__buf_12 output580 (.A(net580),
    .X(sports_o[170]));
 sky130_fd_sc_hd__buf_12 output581 (.A(net581),
    .X(sports_o[171]));
 sky130_fd_sc_hd__buf_12 output582 (.A(net582),
    .X(sports_o[172]));
 sky130_fd_sc_hd__buf_12 output583 (.A(net583),
    .X(sports_o[173]));
 sky130_fd_sc_hd__buf_12 output584 (.A(net584),
    .X(sports_o[174]));
 sky130_fd_sc_hd__buf_12 output585 (.A(net585),
    .X(sports_o[175]));
 sky130_fd_sc_hd__buf_12 output586 (.A(net586),
    .X(sports_o[176]));
 sky130_fd_sc_hd__buf_12 output587 (.A(net587),
    .X(sports_o[177]));
 sky130_fd_sc_hd__buf_12 output588 (.A(net588),
    .X(sports_o[178]));
 sky130_fd_sc_hd__buf_12 output589 (.A(net589),
    .X(sports_o[179]));
 sky130_fd_sc_hd__buf_12 output590 (.A(net590),
    .X(sports_o[17]));
 sky130_fd_sc_hd__buf_12 output591 (.A(net591),
    .X(sports_o[180]));
 sky130_fd_sc_hd__buf_12 output592 (.A(net592),
    .X(sports_o[181]));
 sky130_fd_sc_hd__buf_12 output593 (.A(net593),
    .X(sports_o[182]));
 sky130_fd_sc_hd__buf_12 output594 (.A(net594),
    .X(sports_o[183]));
 sky130_fd_sc_hd__buf_12 output595 (.A(net595),
    .X(sports_o[184]));
 sky130_fd_sc_hd__buf_12 output596 (.A(net596),
    .X(sports_o[185]));
 sky130_fd_sc_hd__buf_12 output597 (.A(net597),
    .X(sports_o[186]));
 sky130_fd_sc_hd__buf_12 output598 (.A(net598),
    .X(sports_o[187]));
 sky130_fd_sc_hd__buf_12 output599 (.A(net599),
    .X(sports_o[188]));
 sky130_fd_sc_hd__buf_12 output600 (.A(net600),
    .X(sports_o[189]));
 sky130_fd_sc_hd__buf_12 output601 (.A(net601),
    .X(sports_o[18]));
 sky130_fd_sc_hd__buf_12 output602 (.A(net602),
    .X(sports_o[190]));
 sky130_fd_sc_hd__buf_12 output603 (.A(net603),
    .X(sports_o[191]));
 sky130_fd_sc_hd__buf_12 output604 (.A(net604),
    .X(sports_o[192]));
 sky130_fd_sc_hd__buf_12 output605 (.A(net605),
    .X(sports_o[193]));
 sky130_fd_sc_hd__buf_12 output606 (.A(net606),
    .X(sports_o[194]));
 sky130_fd_sc_hd__buf_12 output607 (.A(net607),
    .X(sports_o[195]));
 sky130_fd_sc_hd__buf_12 output608 (.A(net608),
    .X(sports_o[196]));
 sky130_fd_sc_hd__buf_12 output609 (.A(net609),
    .X(sports_o[197]));
 sky130_fd_sc_hd__buf_12 output610 (.A(net610),
    .X(sports_o[198]));
 sky130_fd_sc_hd__buf_12 output611 (.A(net611),
    .X(sports_o[199]));
 sky130_fd_sc_hd__buf_12 output612 (.A(net612),
    .X(sports_o[19]));
 sky130_fd_sc_hd__buf_12 output613 (.A(net613),
    .X(sports_o[1]));
 sky130_fd_sc_hd__buf_12 output614 (.A(net614),
    .X(sports_o[200]));
 sky130_fd_sc_hd__buf_12 output615 (.A(net615),
    .X(sports_o[201]));
 sky130_fd_sc_hd__buf_12 output616 (.A(net616),
    .X(sports_o[202]));
 sky130_fd_sc_hd__buf_12 output617 (.A(net617),
    .X(sports_o[203]));
 sky130_fd_sc_hd__buf_12 output618 (.A(net618),
    .X(sports_o[204]));
 sky130_fd_sc_hd__buf_12 output619 (.A(net619),
    .X(sports_o[205]));
 sky130_fd_sc_hd__buf_12 output620 (.A(net620),
    .X(sports_o[206]));
 sky130_fd_sc_hd__buf_12 output621 (.A(net621),
    .X(sports_o[207]));
 sky130_fd_sc_hd__buf_12 output622 (.A(net622),
    .X(sports_o[208]));
 sky130_fd_sc_hd__buf_12 output623 (.A(net623),
    .X(sports_o[209]));
 sky130_fd_sc_hd__buf_12 output624 (.A(net624),
    .X(sports_o[20]));
 sky130_fd_sc_hd__buf_12 output625 (.A(net625),
    .X(sports_o[210]));
 sky130_fd_sc_hd__buf_12 output626 (.A(net626),
    .X(sports_o[211]));
 sky130_fd_sc_hd__buf_12 output627 (.A(net627),
    .X(sports_o[212]));
 sky130_fd_sc_hd__buf_12 output628 (.A(net628),
    .X(sports_o[213]));
 sky130_fd_sc_hd__buf_12 output629 (.A(net629),
    .X(sports_o[214]));
 sky130_fd_sc_hd__buf_12 output630 (.A(net630),
    .X(sports_o[215]));
 sky130_fd_sc_hd__buf_12 output631 (.A(net631),
    .X(sports_o[216]));
 sky130_fd_sc_hd__buf_12 output632 (.A(net632),
    .X(sports_o[217]));
 sky130_fd_sc_hd__buf_12 output633 (.A(net633),
    .X(sports_o[218]));
 sky130_fd_sc_hd__buf_12 output634 (.A(net634),
    .X(sports_o[219]));
 sky130_fd_sc_hd__buf_12 output635 (.A(net635),
    .X(sports_o[21]));
 sky130_fd_sc_hd__buf_12 output636 (.A(net636),
    .X(sports_o[220]));
 sky130_fd_sc_hd__buf_12 output637 (.A(net637),
    .X(sports_o[221]));
 sky130_fd_sc_hd__buf_12 output638 (.A(net638),
    .X(sports_o[222]));
 sky130_fd_sc_hd__buf_12 output639 (.A(net639),
    .X(sports_o[223]));
 sky130_fd_sc_hd__buf_12 output640 (.A(net640),
    .X(sports_o[224]));
 sky130_fd_sc_hd__buf_12 output641 (.A(net641),
    .X(sports_o[225]));
 sky130_fd_sc_hd__buf_12 output642 (.A(net642),
    .X(sports_o[226]));
 sky130_fd_sc_hd__buf_12 output643 (.A(net643),
    .X(sports_o[227]));
 sky130_fd_sc_hd__buf_12 output644 (.A(net644),
    .X(sports_o[22]));
 sky130_fd_sc_hd__buf_12 output645 (.A(net645),
    .X(sports_o[23]));
 sky130_fd_sc_hd__buf_12 output646 (.A(net646),
    .X(sports_o[24]));
 sky130_fd_sc_hd__buf_12 output647 (.A(net647),
    .X(sports_o[25]));
 sky130_fd_sc_hd__buf_12 output648 (.A(net648),
    .X(sports_o[26]));
 sky130_fd_sc_hd__buf_12 output649 (.A(net649),
    .X(sports_o[27]));
 sky130_fd_sc_hd__buf_12 output650 (.A(net650),
    .X(sports_o[28]));
 sky130_fd_sc_hd__buf_12 output651 (.A(net651),
    .X(sports_o[29]));
 sky130_fd_sc_hd__buf_12 output652 (.A(net652),
    .X(sports_o[2]));
 sky130_fd_sc_hd__buf_12 output653 (.A(net653),
    .X(sports_o[30]));
 sky130_fd_sc_hd__buf_12 output654 (.A(net654),
    .X(sports_o[31]));
 sky130_fd_sc_hd__buf_12 output655 (.A(net655),
    .X(sports_o[32]));
 sky130_fd_sc_hd__buf_12 output656 (.A(net656),
    .X(sports_o[33]));
 sky130_fd_sc_hd__buf_12 output657 (.A(net657),
    .X(sports_o[34]));
 sky130_fd_sc_hd__buf_12 output658 (.A(net658),
    .X(sports_o[35]));
 sky130_fd_sc_hd__buf_12 output659 (.A(net659),
    .X(sports_o[36]));
 sky130_fd_sc_hd__buf_12 output660 (.A(net660),
    .X(sports_o[37]));
 sky130_fd_sc_hd__buf_12 output661 (.A(net661),
    .X(sports_o[38]));
 sky130_fd_sc_hd__buf_12 output662 (.A(net662),
    .X(sports_o[39]));
 sky130_fd_sc_hd__buf_12 output663 (.A(net663),
    .X(sports_o[3]));
 sky130_fd_sc_hd__buf_12 output664 (.A(net664),
    .X(sports_o[40]));
 sky130_fd_sc_hd__buf_12 output665 (.A(net665),
    .X(sports_o[41]));
 sky130_fd_sc_hd__buf_12 output666 (.A(net666),
    .X(sports_o[42]));
 sky130_fd_sc_hd__buf_12 output667 (.A(net667),
    .X(sports_o[43]));
 sky130_fd_sc_hd__buf_12 output668 (.A(net668),
    .X(sports_o[44]));
 sky130_fd_sc_hd__buf_12 output669 (.A(net669),
    .X(sports_o[45]));
 sky130_fd_sc_hd__buf_12 output670 (.A(net670),
    .X(sports_o[46]));
 sky130_fd_sc_hd__buf_12 output671 (.A(net671),
    .X(sports_o[47]));
 sky130_fd_sc_hd__buf_12 output672 (.A(net672),
    .X(sports_o[48]));
 sky130_fd_sc_hd__buf_12 output673 (.A(net673),
    .X(sports_o[49]));
 sky130_fd_sc_hd__buf_12 output674 (.A(net674),
    .X(sports_o[4]));
 sky130_fd_sc_hd__buf_12 output675 (.A(net675),
    .X(sports_o[50]));
 sky130_fd_sc_hd__buf_12 output676 (.A(net676),
    .X(sports_o[51]));
 sky130_fd_sc_hd__buf_12 output677 (.A(net677),
    .X(sports_o[52]));
 sky130_fd_sc_hd__buf_12 output678 (.A(net678),
    .X(sports_o[53]));
 sky130_fd_sc_hd__buf_12 output679 (.A(net679),
    .X(sports_o[54]));
 sky130_fd_sc_hd__buf_12 output680 (.A(net680),
    .X(sports_o[55]));
 sky130_fd_sc_hd__buf_12 output681 (.A(net681),
    .X(sports_o[56]));
 sky130_fd_sc_hd__buf_12 output682 (.A(net682),
    .X(sports_o[57]));
 sky130_fd_sc_hd__buf_12 output683 (.A(net683),
    .X(sports_o[58]));
 sky130_fd_sc_hd__buf_12 output684 (.A(net684),
    .X(sports_o[59]));
 sky130_fd_sc_hd__buf_12 output685 (.A(net685),
    .X(sports_o[5]));
 sky130_fd_sc_hd__buf_12 output686 (.A(net686),
    .X(sports_o[60]));
 sky130_fd_sc_hd__buf_12 output687 (.A(net687),
    .X(sports_o[61]));
 sky130_fd_sc_hd__buf_12 output688 (.A(net688),
    .X(sports_o[62]));
 sky130_fd_sc_hd__buf_12 output689 (.A(net689),
    .X(sports_o[63]));
 sky130_fd_sc_hd__buf_12 output690 (.A(net690),
    .X(sports_o[64]));
 sky130_fd_sc_hd__buf_12 output691 (.A(net691),
    .X(sports_o[65]));
 sky130_fd_sc_hd__buf_12 output692 (.A(net692),
    .X(sports_o[66]));
 sky130_fd_sc_hd__buf_12 output693 (.A(net693),
    .X(sports_o[67]));
 sky130_fd_sc_hd__buf_12 output694 (.A(net694),
    .X(sports_o[68]));
 sky130_fd_sc_hd__buf_12 output695 (.A(net695),
    .X(sports_o[69]));
 sky130_fd_sc_hd__buf_12 output696 (.A(net696),
    .X(sports_o[6]));
 sky130_fd_sc_hd__buf_12 output697 (.A(net697),
    .X(sports_o[70]));
 sky130_fd_sc_hd__buf_12 output698 (.A(net698),
    .X(sports_o[71]));
 sky130_fd_sc_hd__buf_12 output699 (.A(net699),
    .X(sports_o[72]));
 sky130_fd_sc_hd__buf_12 output700 (.A(net700),
    .X(sports_o[73]));
 sky130_fd_sc_hd__buf_12 output701 (.A(net701),
    .X(sports_o[74]));
 sky130_fd_sc_hd__buf_12 output702 (.A(net702),
    .X(sports_o[75]));
 sky130_fd_sc_hd__buf_12 output703 (.A(net703),
    .X(sports_o[76]));
 sky130_fd_sc_hd__buf_12 output704 (.A(net704),
    .X(sports_o[77]));
 sky130_fd_sc_hd__buf_12 output705 (.A(net705),
    .X(sports_o[78]));
 sky130_fd_sc_hd__buf_12 output706 (.A(net706),
    .X(sports_o[79]));
 sky130_fd_sc_hd__buf_12 output707 (.A(net707),
    .X(sports_o[7]));
 sky130_fd_sc_hd__buf_12 output708 (.A(net708),
    .X(sports_o[80]));
 sky130_fd_sc_hd__buf_12 output709 (.A(net709),
    .X(sports_o[81]));
 sky130_fd_sc_hd__buf_12 output710 (.A(net710),
    .X(sports_o[82]));
 sky130_fd_sc_hd__buf_12 output711 (.A(net711),
    .X(sports_o[83]));
 sky130_fd_sc_hd__buf_12 output712 (.A(net712),
    .X(sports_o[84]));
 sky130_fd_sc_hd__buf_12 output713 (.A(net713),
    .X(sports_o[85]));
 sky130_fd_sc_hd__buf_12 output714 (.A(net714),
    .X(sports_o[86]));
 sky130_fd_sc_hd__buf_12 output715 (.A(net715),
    .X(sports_o[87]));
 sky130_fd_sc_hd__buf_12 output716 (.A(net716),
    .X(sports_o[88]));
 sky130_fd_sc_hd__buf_12 output717 (.A(net717),
    .X(sports_o[89]));
 sky130_fd_sc_hd__buf_12 output718 (.A(net718),
    .X(sports_o[8]));
 sky130_fd_sc_hd__buf_12 output719 (.A(net719),
    .X(sports_o[90]));
 sky130_fd_sc_hd__buf_12 output720 (.A(net720),
    .X(sports_o[91]));
 sky130_fd_sc_hd__buf_12 output721 (.A(net721),
    .X(sports_o[92]));
 sky130_fd_sc_hd__buf_12 output722 (.A(net722),
    .X(sports_o[93]));
 sky130_fd_sc_hd__buf_12 output723 (.A(net723),
    .X(sports_o[94]));
 sky130_fd_sc_hd__buf_12 output724 (.A(net724),
    .X(sports_o[95]));
 sky130_fd_sc_hd__buf_12 output725 (.A(net725),
    .X(sports_o[96]));
 sky130_fd_sc_hd__buf_12 output726 (.A(net726),
    .X(sports_o[97]));
 sky130_fd_sc_hd__buf_12 output727 (.A(net727),
    .X(sports_o[98]));
 sky130_fd_sc_hd__buf_12 output728 (.A(net728),
    .X(sports_o[99]));
 sky130_fd_sc_hd__buf_12 output729 (.A(net729),
    .X(sports_o[9]));
 sky130_fd_sc_hd__clkbuf_4 wire730 (.A(_1001_),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_4 wire731 (.A(_0691_),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_4 wire732 (.A(_0682_),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_4 wire733 (.A(_0680_),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_4 wire734 (.A(_1019_),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_4 wire735 (.A(_1015_),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_4 wire736 (.A(_1006_),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_4 wire737 (.A(_1004_),
    .X(net737));
endmodule

