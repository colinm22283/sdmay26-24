magic
tech sky130A
magscale 1 2
timestamp 1761157739
<< obsli1 >>
rect 1104 2159 88872 87601
<< obsm1 >>
rect 14 960 89962 89956
<< metal2 >>
rect 2778 89200 2834 90000
rect 3146 89200 3202 90000
rect 3514 89200 3570 90000
rect 3882 89200 3938 90000
rect 4250 89200 4306 90000
rect 4618 89200 4674 90000
rect 4986 89200 5042 90000
rect 5354 89200 5410 90000
rect 5722 89200 5778 90000
rect 6090 89200 6146 90000
rect 6458 89200 6514 90000
rect 6826 89200 6882 90000
rect 7194 89200 7250 90000
rect 7562 89200 7618 90000
rect 7930 89200 7986 90000
rect 8298 89200 8354 90000
rect 8666 89200 8722 90000
rect 9034 89200 9090 90000
rect 9402 89200 9458 90000
rect 9770 89200 9826 90000
rect 10138 89200 10194 90000
rect 10506 89200 10562 90000
rect 10874 89200 10930 90000
rect 11242 89200 11298 90000
rect 11610 89200 11666 90000
rect 11978 89200 12034 90000
rect 12346 89200 12402 90000
rect 12714 89200 12770 90000
rect 13082 89200 13138 90000
rect 13450 89200 13506 90000
rect 13818 89200 13874 90000
rect 14186 89200 14242 90000
rect 14554 89200 14610 90000
rect 14922 89200 14978 90000
rect 15290 89200 15346 90000
rect 15658 89200 15714 90000
rect 16026 89200 16082 90000
rect 16394 89200 16450 90000
rect 16762 89200 16818 90000
rect 17130 89200 17186 90000
rect 17498 89200 17554 90000
rect 17866 89200 17922 90000
rect 18234 89200 18290 90000
rect 18602 89200 18658 90000
rect 18970 89200 19026 90000
rect 19338 89200 19394 90000
rect 19706 89200 19762 90000
rect 20074 89200 20130 90000
rect 20442 89200 20498 90000
rect 20810 89200 20866 90000
rect 21178 89200 21234 90000
rect 21546 89200 21602 90000
rect 21914 89200 21970 90000
rect 22282 89200 22338 90000
rect 22650 89200 22706 90000
rect 23018 89200 23074 90000
rect 23386 89200 23442 90000
rect 23754 89200 23810 90000
rect 24122 89200 24178 90000
rect 24490 89200 24546 90000
rect 24858 89200 24914 90000
rect 25226 89200 25282 90000
rect 25594 89200 25650 90000
rect 25962 89200 26018 90000
rect 26330 89200 26386 90000
rect 26698 89200 26754 90000
rect 27066 89200 27122 90000
rect 27434 89200 27490 90000
rect 27802 89200 27858 90000
rect 28170 89200 28226 90000
rect 28538 89200 28594 90000
rect 28906 89200 28962 90000
rect 29274 89200 29330 90000
rect 29642 89200 29698 90000
rect 30010 89200 30066 90000
rect 30378 89200 30434 90000
rect 30746 89200 30802 90000
rect 31114 89200 31170 90000
rect 31482 89200 31538 90000
rect 31850 89200 31906 90000
rect 32218 89200 32274 90000
rect 32586 89200 32642 90000
rect 32954 89200 33010 90000
rect 33322 89200 33378 90000
rect 33690 89200 33746 90000
rect 34058 89200 34114 90000
rect 34426 89200 34482 90000
rect 34794 89200 34850 90000
rect 35162 89200 35218 90000
rect 35530 89200 35586 90000
rect 35898 89200 35954 90000
rect 36266 89200 36322 90000
rect 36634 89200 36690 90000
rect 37002 89200 37058 90000
rect 37370 89200 37426 90000
rect 37738 89200 37794 90000
rect 38106 89200 38162 90000
rect 38474 89200 38530 90000
rect 38842 89200 38898 90000
rect 39210 89200 39266 90000
rect 39578 89200 39634 90000
rect 39946 89200 40002 90000
rect 40314 89200 40370 90000
rect 40682 89200 40738 90000
rect 41050 89200 41106 90000
rect 41418 89200 41474 90000
rect 41786 89200 41842 90000
rect 42154 89200 42210 90000
rect 42522 89200 42578 90000
rect 42890 89200 42946 90000
rect 43258 89200 43314 90000
rect 43626 89200 43682 90000
rect 43994 89200 44050 90000
rect 44362 89200 44418 90000
rect 44730 89200 44786 90000
rect 45098 89200 45154 90000
rect 45466 89200 45522 90000
rect 45834 89200 45890 90000
rect 46202 89200 46258 90000
rect 46570 89200 46626 90000
rect 46938 89200 46994 90000
rect 47306 89200 47362 90000
rect 47674 89200 47730 90000
rect 48042 89200 48098 90000
rect 48410 89200 48466 90000
rect 48778 89200 48834 90000
rect 49146 89200 49202 90000
rect 49514 89200 49570 90000
rect 49882 89200 49938 90000
rect 50250 89200 50306 90000
rect 50618 89200 50674 90000
rect 50986 89200 51042 90000
rect 51354 89200 51410 90000
rect 51722 89200 51778 90000
rect 52090 89200 52146 90000
rect 52458 89200 52514 90000
rect 52826 89200 52882 90000
rect 53194 89200 53250 90000
rect 53562 89200 53618 90000
rect 53930 89200 53986 90000
rect 54298 89200 54354 90000
rect 54666 89200 54722 90000
rect 55034 89200 55090 90000
rect 55402 89200 55458 90000
rect 55770 89200 55826 90000
rect 56138 89200 56194 90000
rect 56506 89200 56562 90000
rect 56874 89200 56930 90000
rect 57242 89200 57298 90000
rect 57610 89200 57666 90000
rect 57978 89200 58034 90000
rect 58346 89200 58402 90000
rect 58714 89200 58770 90000
rect 59082 89200 59138 90000
rect 59450 89200 59506 90000
rect 59818 89200 59874 90000
rect 60186 89200 60242 90000
rect 60554 89200 60610 90000
rect 60922 89200 60978 90000
rect 61290 89200 61346 90000
rect 61658 89200 61714 90000
rect 62026 89200 62082 90000
rect 62394 89200 62450 90000
rect 62762 89200 62818 90000
rect 63130 89200 63186 90000
rect 63498 89200 63554 90000
rect 63866 89200 63922 90000
rect 64234 89200 64290 90000
rect 64602 89200 64658 90000
rect 64970 89200 65026 90000
rect 65338 89200 65394 90000
rect 65706 89200 65762 90000
rect 66074 89200 66130 90000
rect 66442 89200 66498 90000
rect 66810 89200 66866 90000
rect 67178 89200 67234 90000
rect 67546 89200 67602 90000
rect 67914 89200 67970 90000
rect 68282 89200 68338 90000
rect 68650 89200 68706 90000
rect 69018 89200 69074 90000
rect 69386 89200 69442 90000
rect 69754 89200 69810 90000
rect 70122 89200 70178 90000
rect 70490 89200 70546 90000
rect 70858 89200 70914 90000
rect 71226 89200 71282 90000
rect 71594 89200 71650 90000
rect 71962 89200 72018 90000
rect 72330 89200 72386 90000
rect 72698 89200 72754 90000
rect 73066 89200 73122 90000
rect 73434 89200 73490 90000
rect 73802 89200 73858 90000
rect 74170 89200 74226 90000
rect 74538 89200 74594 90000
rect 74906 89200 74962 90000
rect 75274 89200 75330 90000
rect 75642 89200 75698 90000
rect 76010 89200 76066 90000
rect 76378 89200 76434 90000
rect 76746 89200 76802 90000
rect 77114 89200 77170 90000
rect 77482 89200 77538 90000
rect 77850 89200 77906 90000
rect 78218 89200 78274 90000
rect 78586 89200 78642 90000
rect 78954 89200 79010 90000
rect 79322 89200 79378 90000
rect 79690 89200 79746 90000
rect 80058 89200 80114 90000
rect 80426 89200 80482 90000
rect 80794 89200 80850 90000
rect 81162 89200 81218 90000
rect 81530 89200 81586 90000
rect 81898 89200 81954 90000
rect 82266 89200 82322 90000
rect 82634 89200 82690 90000
rect 83002 89200 83058 90000
rect 83370 89200 83426 90000
rect 83738 89200 83794 90000
rect 84106 89200 84162 90000
rect 84474 89200 84530 90000
rect 84842 89200 84898 90000
rect 85210 89200 85266 90000
rect 85578 89200 85634 90000
rect 85946 89200 86002 90000
rect 86314 89200 86370 90000
rect 86682 89200 86738 90000
rect 87050 89200 87106 90000
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9218 0 9274 800
rect 9862 0 9918 800
rect 10506 0 10562 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 13082 0 13138 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16302 0 16358 800
rect 16946 0 17002 800
rect 17590 0 17646 800
rect 18234 0 18290 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 24030 0 24086 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 25962 0 26018 800
rect 26606 0 26662 800
rect 27250 0 27306 800
rect 27894 0 27950 800
rect 28538 0 28594 800
rect 29182 0 29238 800
rect 29826 0 29882 800
rect 30470 0 30526 800
rect 31114 0 31170 800
rect 31758 0 31814 800
rect 32402 0 32458 800
rect 33046 0 33102 800
rect 33690 0 33746 800
rect 34334 0 34390 800
rect 34978 0 35034 800
rect 35622 0 35678 800
rect 36266 0 36322 800
rect 36910 0 36966 800
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38842 0 38898 800
rect 39486 0 39542 800
rect 40130 0 40186 800
rect 40774 0 40830 800
rect 41418 0 41474 800
rect 42062 0 42118 800
rect 42706 0 42762 800
rect 43350 0 43406 800
rect 43994 0 44050 800
rect 44638 0 44694 800
rect 45282 0 45338 800
rect 45926 0 45982 800
rect 46570 0 46626 800
rect 47214 0 47270 800
rect 47858 0 47914 800
rect 48502 0 48558 800
rect 49146 0 49202 800
rect 49790 0 49846 800
rect 50434 0 50490 800
rect 51078 0 51134 800
rect 51722 0 51778 800
rect 52366 0 52422 800
rect 53010 0 53066 800
rect 53654 0 53710 800
rect 54298 0 54354 800
rect 54942 0 54998 800
rect 55586 0 55642 800
rect 56230 0 56286 800
rect 56874 0 56930 800
rect 57518 0 57574 800
rect 58162 0 58218 800
rect 58806 0 58862 800
rect 59450 0 59506 800
rect 60094 0 60150 800
rect 60738 0 60794 800
rect 61382 0 61438 800
rect 62026 0 62082 800
rect 62670 0 62726 800
rect 63314 0 63370 800
rect 63958 0 64014 800
rect 64602 0 64658 800
rect 65246 0 65302 800
rect 65890 0 65946 800
rect 66534 0 66590 800
rect 67178 0 67234 800
rect 67822 0 67878 800
rect 68466 0 68522 800
rect 69110 0 69166 800
rect 69754 0 69810 800
rect 70398 0 70454 800
rect 71042 0 71098 800
rect 71686 0 71742 800
rect 72330 0 72386 800
rect 72974 0 73030 800
rect 73618 0 73674 800
rect 74262 0 74318 800
rect 74906 0 74962 800
rect 75550 0 75606 800
rect 76194 0 76250 800
rect 76838 0 76894 800
rect 77482 0 77538 800
rect 78126 0 78182 800
rect 78770 0 78826 800
rect 79414 0 79470 800
rect 80058 0 80114 800
rect 80702 0 80758 800
rect 81346 0 81402 800
rect 81990 0 82046 800
rect 82634 0 82690 800
rect 83278 0 83334 800
rect 83922 0 83978 800
rect 84566 0 84622 800
rect 85210 0 85266 800
rect 85854 0 85910 800
rect 86498 0 86554 800
rect 87142 0 87198 800
rect 87786 0 87842 800
rect 88430 0 88486 800
<< obsm2 >>
rect 20 89144 2722 89962
rect 2890 89144 3090 89962
rect 3258 89144 3458 89962
rect 3626 89144 3826 89962
rect 3994 89144 4194 89962
rect 4362 89144 4562 89962
rect 4730 89144 4930 89962
rect 5098 89144 5298 89962
rect 5466 89144 5666 89962
rect 5834 89144 6034 89962
rect 6202 89144 6402 89962
rect 6570 89144 6770 89962
rect 6938 89144 7138 89962
rect 7306 89144 7506 89962
rect 7674 89144 7874 89962
rect 8042 89144 8242 89962
rect 8410 89144 8610 89962
rect 8778 89144 8978 89962
rect 9146 89144 9346 89962
rect 9514 89144 9714 89962
rect 9882 89144 10082 89962
rect 10250 89144 10450 89962
rect 10618 89144 10818 89962
rect 10986 89144 11186 89962
rect 11354 89144 11554 89962
rect 11722 89144 11922 89962
rect 12090 89144 12290 89962
rect 12458 89144 12658 89962
rect 12826 89144 13026 89962
rect 13194 89144 13394 89962
rect 13562 89144 13762 89962
rect 13930 89144 14130 89962
rect 14298 89144 14498 89962
rect 14666 89144 14866 89962
rect 15034 89144 15234 89962
rect 15402 89144 15602 89962
rect 15770 89144 15970 89962
rect 16138 89144 16338 89962
rect 16506 89144 16706 89962
rect 16874 89144 17074 89962
rect 17242 89144 17442 89962
rect 17610 89144 17810 89962
rect 17978 89144 18178 89962
rect 18346 89144 18546 89962
rect 18714 89144 18914 89962
rect 19082 89144 19282 89962
rect 19450 89144 19650 89962
rect 19818 89144 20018 89962
rect 20186 89144 20386 89962
rect 20554 89144 20754 89962
rect 20922 89144 21122 89962
rect 21290 89144 21490 89962
rect 21658 89144 21858 89962
rect 22026 89144 22226 89962
rect 22394 89144 22594 89962
rect 22762 89144 22962 89962
rect 23130 89144 23330 89962
rect 23498 89144 23698 89962
rect 23866 89144 24066 89962
rect 24234 89144 24434 89962
rect 24602 89144 24802 89962
rect 24970 89144 25170 89962
rect 25338 89144 25538 89962
rect 25706 89144 25906 89962
rect 26074 89144 26274 89962
rect 26442 89144 26642 89962
rect 26810 89144 27010 89962
rect 27178 89144 27378 89962
rect 27546 89144 27746 89962
rect 27914 89144 28114 89962
rect 28282 89144 28482 89962
rect 28650 89144 28850 89962
rect 29018 89144 29218 89962
rect 29386 89144 29586 89962
rect 29754 89144 29954 89962
rect 30122 89144 30322 89962
rect 30490 89144 30690 89962
rect 30858 89144 31058 89962
rect 31226 89144 31426 89962
rect 31594 89144 31794 89962
rect 31962 89144 32162 89962
rect 32330 89144 32530 89962
rect 32698 89144 32898 89962
rect 33066 89144 33266 89962
rect 33434 89144 33634 89962
rect 33802 89144 34002 89962
rect 34170 89144 34370 89962
rect 34538 89144 34738 89962
rect 34906 89144 35106 89962
rect 35274 89144 35474 89962
rect 35642 89144 35842 89962
rect 36010 89144 36210 89962
rect 36378 89144 36578 89962
rect 36746 89144 36946 89962
rect 37114 89144 37314 89962
rect 37482 89144 37682 89962
rect 37850 89144 38050 89962
rect 38218 89144 38418 89962
rect 38586 89144 38786 89962
rect 38954 89144 39154 89962
rect 39322 89144 39522 89962
rect 39690 89144 39890 89962
rect 40058 89144 40258 89962
rect 40426 89144 40626 89962
rect 40794 89144 40994 89962
rect 41162 89144 41362 89962
rect 41530 89144 41730 89962
rect 41898 89144 42098 89962
rect 42266 89144 42466 89962
rect 42634 89144 42834 89962
rect 43002 89144 43202 89962
rect 43370 89144 43570 89962
rect 43738 89144 43938 89962
rect 44106 89144 44306 89962
rect 44474 89144 44674 89962
rect 44842 89144 45042 89962
rect 45210 89144 45410 89962
rect 45578 89144 45778 89962
rect 45946 89144 46146 89962
rect 46314 89144 46514 89962
rect 46682 89144 46882 89962
rect 47050 89144 47250 89962
rect 47418 89144 47618 89962
rect 47786 89144 47986 89962
rect 48154 89144 48354 89962
rect 48522 89144 48722 89962
rect 48890 89144 49090 89962
rect 49258 89144 49458 89962
rect 49626 89144 49826 89962
rect 49994 89144 50194 89962
rect 50362 89144 50562 89962
rect 50730 89144 50930 89962
rect 51098 89144 51298 89962
rect 51466 89144 51666 89962
rect 51834 89144 52034 89962
rect 52202 89144 52402 89962
rect 52570 89144 52770 89962
rect 52938 89144 53138 89962
rect 53306 89144 53506 89962
rect 53674 89144 53874 89962
rect 54042 89144 54242 89962
rect 54410 89144 54610 89962
rect 54778 89144 54978 89962
rect 55146 89144 55346 89962
rect 55514 89144 55714 89962
rect 55882 89144 56082 89962
rect 56250 89144 56450 89962
rect 56618 89144 56818 89962
rect 56986 89144 57186 89962
rect 57354 89144 57554 89962
rect 57722 89144 57922 89962
rect 58090 89144 58290 89962
rect 58458 89144 58658 89962
rect 58826 89144 59026 89962
rect 59194 89144 59394 89962
rect 59562 89144 59762 89962
rect 59930 89144 60130 89962
rect 60298 89144 60498 89962
rect 60666 89144 60866 89962
rect 61034 89144 61234 89962
rect 61402 89144 61602 89962
rect 61770 89144 61970 89962
rect 62138 89144 62338 89962
rect 62506 89144 62706 89962
rect 62874 89144 63074 89962
rect 63242 89144 63442 89962
rect 63610 89144 63810 89962
rect 63978 89144 64178 89962
rect 64346 89144 64546 89962
rect 64714 89144 64914 89962
rect 65082 89144 65282 89962
rect 65450 89144 65650 89962
rect 65818 89144 66018 89962
rect 66186 89144 66386 89962
rect 66554 89144 66754 89962
rect 66922 89144 67122 89962
rect 67290 89144 67490 89962
rect 67658 89144 67858 89962
rect 68026 89144 68226 89962
rect 68394 89144 68594 89962
rect 68762 89144 68962 89962
rect 69130 89144 69330 89962
rect 69498 89144 69698 89962
rect 69866 89144 70066 89962
rect 70234 89144 70434 89962
rect 70602 89144 70802 89962
rect 70970 89144 71170 89962
rect 71338 89144 71538 89962
rect 71706 89144 71906 89962
rect 72074 89144 72274 89962
rect 72442 89144 72642 89962
rect 72810 89144 73010 89962
rect 73178 89144 73378 89962
rect 73546 89144 73746 89962
rect 73914 89144 74114 89962
rect 74282 89144 74482 89962
rect 74650 89144 74850 89962
rect 75018 89144 75218 89962
rect 75386 89144 75586 89962
rect 75754 89144 75954 89962
rect 76122 89144 76322 89962
rect 76490 89144 76690 89962
rect 76858 89144 77058 89962
rect 77226 89144 77426 89962
rect 77594 89144 77794 89962
rect 77962 89144 78162 89962
rect 78330 89144 78530 89962
rect 78698 89144 78898 89962
rect 79066 89144 79266 89962
rect 79434 89144 79634 89962
rect 79802 89144 80002 89962
rect 80170 89144 80370 89962
rect 80538 89144 80738 89962
rect 80906 89144 81106 89962
rect 81274 89144 81474 89962
rect 81642 89144 81842 89962
rect 82010 89144 82210 89962
rect 82378 89144 82578 89962
rect 82746 89144 82946 89962
rect 83114 89144 83314 89962
rect 83482 89144 83682 89962
rect 83850 89144 84050 89962
rect 84218 89144 84418 89962
rect 84586 89144 84786 89962
rect 84954 89144 85154 89962
rect 85322 89144 85522 89962
rect 85690 89144 85890 89962
rect 86058 89144 86258 89962
rect 86426 89144 86626 89962
rect 86794 89144 86994 89962
rect 87162 89144 89956 89962
rect 20 856 89956 89144
rect 20 734 1434 856
rect 1602 734 2078 856
rect 2246 734 2722 856
rect 2890 734 3366 856
rect 3534 734 4010 856
rect 4178 734 4654 856
rect 4822 734 5298 856
rect 5466 734 5942 856
rect 6110 734 6586 856
rect 6754 734 7230 856
rect 7398 734 7874 856
rect 8042 734 8518 856
rect 8686 734 9162 856
rect 9330 734 9806 856
rect 9974 734 10450 856
rect 10618 734 11094 856
rect 11262 734 11738 856
rect 11906 734 12382 856
rect 12550 734 13026 856
rect 13194 734 13670 856
rect 13838 734 14314 856
rect 14482 734 14958 856
rect 15126 734 15602 856
rect 15770 734 16246 856
rect 16414 734 16890 856
rect 17058 734 17534 856
rect 17702 734 18178 856
rect 18346 734 18822 856
rect 18990 734 19466 856
rect 19634 734 20110 856
rect 20278 734 20754 856
rect 20922 734 21398 856
rect 21566 734 22042 856
rect 22210 734 22686 856
rect 22854 734 23330 856
rect 23498 734 23974 856
rect 24142 734 24618 856
rect 24786 734 25262 856
rect 25430 734 25906 856
rect 26074 734 26550 856
rect 26718 734 27194 856
rect 27362 734 27838 856
rect 28006 734 28482 856
rect 28650 734 29126 856
rect 29294 734 29770 856
rect 29938 734 30414 856
rect 30582 734 31058 856
rect 31226 734 31702 856
rect 31870 734 32346 856
rect 32514 734 32990 856
rect 33158 734 33634 856
rect 33802 734 34278 856
rect 34446 734 34922 856
rect 35090 734 35566 856
rect 35734 734 36210 856
rect 36378 734 36854 856
rect 37022 734 37498 856
rect 37666 734 38142 856
rect 38310 734 38786 856
rect 38954 734 39430 856
rect 39598 734 40074 856
rect 40242 734 40718 856
rect 40886 734 41362 856
rect 41530 734 42006 856
rect 42174 734 42650 856
rect 42818 734 43294 856
rect 43462 734 43938 856
rect 44106 734 44582 856
rect 44750 734 45226 856
rect 45394 734 45870 856
rect 46038 734 46514 856
rect 46682 734 47158 856
rect 47326 734 47802 856
rect 47970 734 48446 856
rect 48614 734 49090 856
rect 49258 734 49734 856
rect 49902 734 50378 856
rect 50546 734 51022 856
rect 51190 734 51666 856
rect 51834 734 52310 856
rect 52478 734 52954 856
rect 53122 734 53598 856
rect 53766 734 54242 856
rect 54410 734 54886 856
rect 55054 734 55530 856
rect 55698 734 56174 856
rect 56342 734 56818 856
rect 56986 734 57462 856
rect 57630 734 58106 856
rect 58274 734 58750 856
rect 58918 734 59394 856
rect 59562 734 60038 856
rect 60206 734 60682 856
rect 60850 734 61326 856
rect 61494 734 61970 856
rect 62138 734 62614 856
rect 62782 734 63258 856
rect 63426 734 63902 856
rect 64070 734 64546 856
rect 64714 734 65190 856
rect 65358 734 65834 856
rect 66002 734 66478 856
rect 66646 734 67122 856
rect 67290 734 67766 856
rect 67934 734 68410 856
rect 68578 734 69054 856
rect 69222 734 69698 856
rect 69866 734 70342 856
rect 70510 734 70986 856
rect 71154 734 71630 856
rect 71798 734 72274 856
rect 72442 734 72918 856
rect 73086 734 73562 856
rect 73730 734 74206 856
rect 74374 734 74850 856
rect 75018 734 75494 856
rect 75662 734 76138 856
rect 76306 734 76782 856
rect 76950 734 77426 856
rect 77594 734 78070 856
rect 78238 734 78714 856
rect 78882 734 79358 856
rect 79526 734 80002 856
rect 80170 734 80646 856
rect 80814 734 81290 856
rect 81458 734 81934 856
rect 82102 734 82578 856
rect 82746 734 83222 856
rect 83390 734 83866 856
rect 84034 734 84510 856
rect 84678 734 85154 856
rect 85322 734 85798 856
rect 85966 734 86442 856
rect 86610 734 87086 856
rect 87254 734 87730 856
rect 87898 734 88374 856
rect 88542 734 89956 856
<< metal3 >>
rect 89200 81608 90000 81728
rect 89200 81064 90000 81184
rect 89200 80520 90000 80640
rect 89200 79976 90000 80096
rect 89200 79432 90000 79552
rect 89200 78888 90000 79008
rect 89200 78344 90000 78464
rect 89200 77800 90000 77920
rect 89200 77256 90000 77376
rect 89200 76712 90000 76832
rect 89200 76168 90000 76288
rect 0 75624 800 75744
rect 89200 75624 90000 75744
rect 0 75352 800 75472
rect 0 75080 800 75200
rect 89200 75080 90000 75200
rect 0 74808 800 74928
rect 0 74536 800 74656
rect 89200 74536 90000 74656
rect 0 74264 800 74384
rect 0 73992 800 74112
rect 89200 73992 90000 74112
rect 0 73720 800 73840
rect 0 73448 800 73568
rect 89200 73448 90000 73568
rect 0 73176 800 73296
rect 0 72904 800 73024
rect 89200 72904 90000 73024
rect 0 72632 800 72752
rect 0 72360 800 72480
rect 89200 72360 90000 72480
rect 0 72088 800 72208
rect 0 71816 800 71936
rect 89200 71816 90000 71936
rect 0 71544 800 71664
rect 0 71272 800 71392
rect 89200 71272 90000 71392
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 89200 70728 90000 70848
rect 0 70456 800 70576
rect 0 70184 800 70304
rect 89200 70184 90000 70304
rect 0 69912 800 70032
rect 0 69640 800 69760
rect 89200 69640 90000 69760
rect 0 69368 800 69488
rect 0 69096 800 69216
rect 89200 69096 90000 69216
rect 0 68824 800 68944
rect 0 68552 800 68672
rect 89200 68552 90000 68672
rect 0 68280 800 68400
rect 0 68008 800 68128
rect 89200 68008 90000 68128
rect 0 67736 800 67856
rect 0 67464 800 67584
rect 89200 67464 90000 67584
rect 0 67192 800 67312
rect 0 66920 800 67040
rect 89200 66920 90000 67040
rect 0 66648 800 66768
rect 0 66376 800 66496
rect 89200 66376 90000 66496
rect 0 66104 800 66224
rect 0 65832 800 65952
rect 89200 65832 90000 65952
rect 0 65560 800 65680
rect 0 65288 800 65408
rect 89200 65288 90000 65408
rect 0 65016 800 65136
rect 0 64744 800 64864
rect 89200 64744 90000 64864
rect 0 64472 800 64592
rect 0 64200 800 64320
rect 89200 64200 90000 64320
rect 0 63928 800 64048
rect 0 63656 800 63776
rect 89200 63656 90000 63776
rect 0 63384 800 63504
rect 0 63112 800 63232
rect 89200 63112 90000 63232
rect 0 62840 800 62960
rect 0 62568 800 62688
rect 89200 62568 90000 62688
rect 0 62296 800 62416
rect 0 62024 800 62144
rect 89200 62024 90000 62144
rect 0 61752 800 61872
rect 0 61480 800 61600
rect 89200 61480 90000 61600
rect 0 61208 800 61328
rect 0 60936 800 61056
rect 89200 60936 90000 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 89200 60392 90000 60512
rect 0 60120 800 60240
rect 0 59848 800 59968
rect 89200 59848 90000 59968
rect 0 59576 800 59696
rect 0 59304 800 59424
rect 89200 59304 90000 59424
rect 0 59032 800 59152
rect 0 58760 800 58880
rect 89200 58760 90000 58880
rect 0 58488 800 58608
rect 0 58216 800 58336
rect 89200 58216 90000 58336
rect 0 57944 800 58064
rect 0 57672 800 57792
rect 89200 57672 90000 57792
rect 0 57400 800 57520
rect 0 57128 800 57248
rect 89200 57128 90000 57248
rect 0 56856 800 56976
rect 0 56584 800 56704
rect 89200 56584 90000 56704
rect 0 56312 800 56432
rect 0 56040 800 56160
rect 89200 56040 90000 56160
rect 0 55768 800 55888
rect 0 55496 800 55616
rect 89200 55496 90000 55616
rect 0 55224 800 55344
rect 0 54952 800 55072
rect 89200 54952 90000 55072
rect 0 54680 800 54800
rect 0 54408 800 54528
rect 89200 54408 90000 54528
rect 0 54136 800 54256
rect 0 53864 800 53984
rect 89200 53864 90000 53984
rect 0 53592 800 53712
rect 0 53320 800 53440
rect 89200 53320 90000 53440
rect 0 53048 800 53168
rect 0 52776 800 52896
rect 89200 52776 90000 52896
rect 0 52504 800 52624
rect 0 52232 800 52352
rect 89200 52232 90000 52352
rect 0 51960 800 52080
rect 0 51688 800 51808
rect 89200 51688 90000 51808
rect 0 51416 800 51536
rect 0 51144 800 51264
rect 89200 51144 90000 51264
rect 0 50872 800 50992
rect 0 50600 800 50720
rect 89200 50600 90000 50720
rect 0 50328 800 50448
rect 0 50056 800 50176
rect 89200 50056 90000 50176
rect 0 49784 800 49904
rect 0 49512 800 49632
rect 89200 49512 90000 49632
rect 0 49240 800 49360
rect 0 48968 800 49088
rect 89200 48968 90000 49088
rect 0 48696 800 48816
rect 0 48424 800 48544
rect 89200 48424 90000 48544
rect 0 48152 800 48272
rect 0 47880 800 48000
rect 89200 47880 90000 48000
rect 0 47608 800 47728
rect 0 47336 800 47456
rect 89200 47336 90000 47456
rect 0 47064 800 47184
rect 0 46792 800 46912
rect 89200 46792 90000 46912
rect 0 46520 800 46640
rect 0 46248 800 46368
rect 89200 46248 90000 46368
rect 0 45976 800 46096
rect 0 45704 800 45824
rect 89200 45704 90000 45824
rect 0 45432 800 45552
rect 0 45160 800 45280
rect 89200 45160 90000 45280
rect 0 44888 800 45008
rect 0 44616 800 44736
rect 89200 44616 90000 44736
rect 0 44344 800 44464
rect 0 44072 800 44192
rect 89200 44072 90000 44192
rect 0 43800 800 43920
rect 0 43528 800 43648
rect 89200 43528 90000 43648
rect 0 43256 800 43376
rect 0 42984 800 43104
rect 89200 42984 90000 43104
rect 0 42712 800 42832
rect 0 42440 800 42560
rect 89200 42440 90000 42560
rect 0 42168 800 42288
rect 0 41896 800 42016
rect 89200 41896 90000 42016
rect 0 41624 800 41744
rect 0 41352 800 41472
rect 89200 41352 90000 41472
rect 0 41080 800 41200
rect 0 40808 800 40928
rect 89200 40808 90000 40928
rect 0 40536 800 40656
rect 0 40264 800 40384
rect 89200 40264 90000 40384
rect 0 39992 800 40112
rect 0 39720 800 39840
rect 89200 39720 90000 39840
rect 0 39448 800 39568
rect 0 39176 800 39296
rect 89200 39176 90000 39296
rect 0 38904 800 39024
rect 0 38632 800 38752
rect 89200 38632 90000 38752
rect 0 38360 800 38480
rect 0 38088 800 38208
rect 89200 38088 90000 38208
rect 0 37816 800 37936
rect 0 37544 800 37664
rect 89200 37544 90000 37664
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 89200 37000 90000 37120
rect 0 36728 800 36848
rect 0 36456 800 36576
rect 89200 36456 90000 36576
rect 0 36184 800 36304
rect 0 35912 800 36032
rect 89200 35912 90000 36032
rect 0 35640 800 35760
rect 0 35368 800 35488
rect 89200 35368 90000 35488
rect 0 35096 800 35216
rect 0 34824 800 34944
rect 89200 34824 90000 34944
rect 0 34552 800 34672
rect 0 34280 800 34400
rect 89200 34280 90000 34400
rect 0 34008 800 34128
rect 0 33736 800 33856
rect 89200 33736 90000 33856
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 89200 33192 90000 33312
rect 0 32920 800 33040
rect 0 32648 800 32768
rect 89200 32648 90000 32768
rect 0 32376 800 32496
rect 0 32104 800 32224
rect 89200 32104 90000 32224
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 89200 31560 90000 31680
rect 0 31288 800 31408
rect 0 31016 800 31136
rect 89200 31016 90000 31136
rect 0 30744 800 30864
rect 0 30472 800 30592
rect 89200 30472 90000 30592
rect 0 30200 800 30320
rect 0 29928 800 30048
rect 89200 29928 90000 30048
rect 0 29656 800 29776
rect 0 29384 800 29504
rect 89200 29384 90000 29504
rect 0 29112 800 29232
rect 0 28840 800 28960
rect 89200 28840 90000 28960
rect 0 28568 800 28688
rect 0 28296 800 28416
rect 89200 28296 90000 28416
rect 0 28024 800 28144
rect 0 27752 800 27872
rect 89200 27752 90000 27872
rect 0 27480 800 27600
rect 0 27208 800 27328
rect 89200 27208 90000 27328
rect 0 26936 800 27056
rect 0 26664 800 26784
rect 89200 26664 90000 26784
rect 0 26392 800 26512
rect 0 26120 800 26240
rect 89200 26120 90000 26240
rect 0 25848 800 25968
rect 0 25576 800 25696
rect 89200 25576 90000 25696
rect 0 25304 800 25424
rect 0 25032 800 25152
rect 89200 25032 90000 25152
rect 0 24760 800 24880
rect 0 24488 800 24608
rect 89200 24488 90000 24608
rect 0 24216 800 24336
rect 0 23944 800 24064
rect 89200 23944 90000 24064
rect 0 23672 800 23792
rect 0 23400 800 23520
rect 89200 23400 90000 23520
rect 0 23128 800 23248
rect 0 22856 800 22976
rect 89200 22856 90000 22976
rect 0 22584 800 22704
rect 0 22312 800 22432
rect 89200 22312 90000 22432
rect 0 22040 800 22160
rect 0 21768 800 21888
rect 89200 21768 90000 21888
rect 0 21496 800 21616
rect 0 21224 800 21344
rect 89200 21224 90000 21344
rect 0 20952 800 21072
rect 0 20680 800 20800
rect 89200 20680 90000 20800
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 89200 20136 90000 20256
rect 0 19864 800 19984
rect 0 19592 800 19712
rect 89200 19592 90000 19712
rect 0 19320 800 19440
rect 0 19048 800 19168
rect 89200 19048 90000 19168
rect 0 18776 800 18896
rect 0 18504 800 18624
rect 89200 18504 90000 18624
rect 0 18232 800 18352
rect 0 17960 800 18080
rect 89200 17960 90000 18080
rect 0 17688 800 17808
rect 0 17416 800 17536
rect 89200 17416 90000 17536
rect 0 17144 800 17264
rect 0 16872 800 16992
rect 89200 16872 90000 16992
rect 0 16600 800 16720
rect 0 16328 800 16448
rect 89200 16328 90000 16448
rect 0 16056 800 16176
rect 0 15784 800 15904
rect 89200 15784 90000 15904
rect 0 15512 800 15632
rect 0 15240 800 15360
rect 89200 15240 90000 15360
rect 0 14968 800 15088
rect 0 14696 800 14816
rect 89200 14696 90000 14816
rect 0 14424 800 14544
rect 0 14152 800 14272
rect 89200 14152 90000 14272
rect 0 13880 800 14000
rect 89200 13608 90000 13728
rect 89200 13064 90000 13184
rect 89200 12520 90000 12640
rect 89200 11976 90000 12096
rect 89200 11432 90000 11552
rect 89200 10888 90000 11008
rect 89200 10344 90000 10464
rect 89200 9800 90000 9920
rect 89200 9256 90000 9376
rect 89200 8712 90000 8832
rect 89200 8168 90000 8288
<< obsm3 >>
rect 800 81808 89227 89861
rect 800 81528 89120 81808
rect 800 81264 89227 81528
rect 800 80984 89120 81264
rect 800 80720 89227 80984
rect 800 80440 89120 80720
rect 800 80176 89227 80440
rect 800 79896 89120 80176
rect 800 79632 89227 79896
rect 800 79352 89120 79632
rect 800 79088 89227 79352
rect 800 78808 89120 79088
rect 800 78544 89227 78808
rect 800 78264 89120 78544
rect 800 78000 89227 78264
rect 800 77720 89120 78000
rect 800 77456 89227 77720
rect 800 77176 89120 77456
rect 800 76912 89227 77176
rect 800 76632 89120 76912
rect 800 76368 89227 76632
rect 800 76088 89120 76368
rect 800 75824 89227 76088
rect 880 75544 89120 75824
rect 880 75280 89227 75544
rect 880 75000 89120 75280
rect 880 74736 89227 75000
rect 880 74456 89120 74736
rect 880 74192 89227 74456
rect 880 73912 89120 74192
rect 880 73648 89227 73912
rect 880 73368 89120 73648
rect 880 73104 89227 73368
rect 880 72824 89120 73104
rect 880 72560 89227 72824
rect 880 72280 89120 72560
rect 880 72016 89227 72280
rect 880 71736 89120 72016
rect 880 71472 89227 71736
rect 880 71192 89120 71472
rect 880 70928 89227 71192
rect 880 70648 89120 70928
rect 880 70384 89227 70648
rect 880 70104 89120 70384
rect 880 69840 89227 70104
rect 880 69560 89120 69840
rect 880 69296 89227 69560
rect 880 69016 89120 69296
rect 880 68752 89227 69016
rect 880 68472 89120 68752
rect 880 68208 89227 68472
rect 880 67928 89120 68208
rect 880 67664 89227 67928
rect 880 67384 89120 67664
rect 880 67120 89227 67384
rect 880 66840 89120 67120
rect 880 66576 89227 66840
rect 880 66296 89120 66576
rect 880 66032 89227 66296
rect 880 65752 89120 66032
rect 880 65488 89227 65752
rect 880 65208 89120 65488
rect 880 64944 89227 65208
rect 880 64664 89120 64944
rect 880 64400 89227 64664
rect 880 64120 89120 64400
rect 880 63856 89227 64120
rect 880 63576 89120 63856
rect 880 63312 89227 63576
rect 880 63032 89120 63312
rect 880 62768 89227 63032
rect 880 62488 89120 62768
rect 880 62224 89227 62488
rect 880 61944 89120 62224
rect 880 61680 89227 61944
rect 880 61400 89120 61680
rect 880 61136 89227 61400
rect 880 60856 89120 61136
rect 880 60592 89227 60856
rect 880 60312 89120 60592
rect 880 60048 89227 60312
rect 880 59768 89120 60048
rect 880 59504 89227 59768
rect 880 59224 89120 59504
rect 880 58960 89227 59224
rect 880 58680 89120 58960
rect 880 58416 89227 58680
rect 880 58136 89120 58416
rect 880 57872 89227 58136
rect 880 57592 89120 57872
rect 880 57328 89227 57592
rect 880 57048 89120 57328
rect 880 56784 89227 57048
rect 880 56504 89120 56784
rect 880 56240 89227 56504
rect 880 55960 89120 56240
rect 880 55696 89227 55960
rect 880 55416 89120 55696
rect 880 55152 89227 55416
rect 880 54872 89120 55152
rect 880 54608 89227 54872
rect 880 54328 89120 54608
rect 880 54064 89227 54328
rect 880 53784 89120 54064
rect 880 53520 89227 53784
rect 880 53240 89120 53520
rect 880 52976 89227 53240
rect 880 52696 89120 52976
rect 880 52432 89227 52696
rect 880 52152 89120 52432
rect 880 51888 89227 52152
rect 880 51608 89120 51888
rect 880 51344 89227 51608
rect 880 51064 89120 51344
rect 880 50800 89227 51064
rect 880 50520 89120 50800
rect 880 50256 89227 50520
rect 880 49976 89120 50256
rect 880 49712 89227 49976
rect 880 49432 89120 49712
rect 880 49168 89227 49432
rect 880 48888 89120 49168
rect 880 48624 89227 48888
rect 880 48344 89120 48624
rect 880 48080 89227 48344
rect 880 47800 89120 48080
rect 880 47536 89227 47800
rect 880 47256 89120 47536
rect 880 46992 89227 47256
rect 880 46712 89120 46992
rect 880 46448 89227 46712
rect 880 46168 89120 46448
rect 880 45904 89227 46168
rect 880 45624 89120 45904
rect 880 45360 89227 45624
rect 880 45080 89120 45360
rect 880 44816 89227 45080
rect 880 44536 89120 44816
rect 880 44272 89227 44536
rect 880 43992 89120 44272
rect 880 43728 89227 43992
rect 880 43448 89120 43728
rect 880 43184 89227 43448
rect 880 42904 89120 43184
rect 880 42640 89227 42904
rect 880 42360 89120 42640
rect 880 42096 89227 42360
rect 880 41816 89120 42096
rect 880 41552 89227 41816
rect 880 41272 89120 41552
rect 880 41008 89227 41272
rect 880 40728 89120 41008
rect 880 40464 89227 40728
rect 880 40184 89120 40464
rect 880 39920 89227 40184
rect 880 39640 89120 39920
rect 880 39376 89227 39640
rect 880 39096 89120 39376
rect 880 38832 89227 39096
rect 880 38552 89120 38832
rect 880 38288 89227 38552
rect 880 38008 89120 38288
rect 880 37744 89227 38008
rect 880 37464 89120 37744
rect 880 37200 89227 37464
rect 880 36920 89120 37200
rect 880 36656 89227 36920
rect 880 36376 89120 36656
rect 880 36112 89227 36376
rect 880 35832 89120 36112
rect 880 35568 89227 35832
rect 880 35288 89120 35568
rect 880 35024 89227 35288
rect 880 34744 89120 35024
rect 880 34480 89227 34744
rect 880 34200 89120 34480
rect 880 33936 89227 34200
rect 880 33656 89120 33936
rect 880 33392 89227 33656
rect 880 33112 89120 33392
rect 880 32848 89227 33112
rect 880 32568 89120 32848
rect 880 32304 89227 32568
rect 880 32024 89120 32304
rect 880 31760 89227 32024
rect 880 31480 89120 31760
rect 880 31216 89227 31480
rect 880 30936 89120 31216
rect 880 30672 89227 30936
rect 880 30392 89120 30672
rect 880 30128 89227 30392
rect 880 29848 89120 30128
rect 880 29584 89227 29848
rect 880 29304 89120 29584
rect 880 29040 89227 29304
rect 880 28760 89120 29040
rect 880 28496 89227 28760
rect 880 28216 89120 28496
rect 880 27952 89227 28216
rect 880 27672 89120 27952
rect 880 27408 89227 27672
rect 880 27128 89120 27408
rect 880 26864 89227 27128
rect 880 26584 89120 26864
rect 880 26320 89227 26584
rect 880 26040 89120 26320
rect 880 25776 89227 26040
rect 880 25496 89120 25776
rect 880 25232 89227 25496
rect 880 24952 89120 25232
rect 880 24688 89227 24952
rect 880 24408 89120 24688
rect 880 24144 89227 24408
rect 880 23864 89120 24144
rect 880 23600 89227 23864
rect 880 23320 89120 23600
rect 880 23056 89227 23320
rect 880 22776 89120 23056
rect 880 22512 89227 22776
rect 880 22232 89120 22512
rect 880 21968 89227 22232
rect 880 21688 89120 21968
rect 880 21424 89227 21688
rect 880 21144 89120 21424
rect 880 20880 89227 21144
rect 880 20600 89120 20880
rect 880 20336 89227 20600
rect 880 20056 89120 20336
rect 880 19792 89227 20056
rect 880 19512 89120 19792
rect 880 19248 89227 19512
rect 880 18968 89120 19248
rect 880 18704 89227 18968
rect 880 18424 89120 18704
rect 880 18160 89227 18424
rect 880 17880 89120 18160
rect 880 17616 89227 17880
rect 880 17336 89120 17616
rect 880 17072 89227 17336
rect 880 16792 89120 17072
rect 880 16528 89227 16792
rect 880 16248 89120 16528
rect 880 15984 89227 16248
rect 880 15704 89120 15984
rect 880 15440 89227 15704
rect 880 15160 89120 15440
rect 880 14896 89227 15160
rect 880 14616 89120 14896
rect 880 14352 89227 14616
rect 880 14072 89120 14352
rect 880 13808 89227 14072
rect 880 13800 89120 13808
rect 800 13528 89120 13800
rect 800 13264 89227 13528
rect 800 12984 89120 13264
rect 800 12720 89227 12984
rect 800 12440 89120 12720
rect 800 12176 89227 12440
rect 800 11896 89120 12176
rect 800 11632 89227 11896
rect 800 11352 89120 11632
rect 800 11088 89227 11352
rect 800 10808 89120 11088
rect 800 10544 89227 10808
rect 800 10264 89120 10544
rect 800 10000 89227 10264
rect 800 9720 89120 10000
rect 800 9456 89227 9720
rect 800 9176 89120 9456
rect 800 8912 89227 9176
rect 800 8632 89120 8912
rect 800 8368 89227 8632
rect 800 8088 89120 8368
rect 800 1123 89227 8088
<< metal4 >>
rect 4208 2128 4528 87632
rect 19568 2128 19888 87632
rect 34928 2128 35248 87632
rect 50288 2128 50608 87632
rect 65648 2128 65968 87632
rect 81008 2128 81328 87632
<< obsm4 >>
rect 430 87712 88813 89861
rect 430 2048 4128 87712
rect 4608 2048 19488 87712
rect 19968 2048 34848 87712
rect 35328 2048 50208 87712
rect 50688 2048 65568 87712
rect 66048 2048 80928 87712
rect 81408 2048 88813 87712
rect 430 1123 88813 2048
<< labels >>
rlabel metal2 s 2778 89200 2834 90000 6 clk_i
port 1 nsew signal input
rlabel metal2 s 3514 89200 3570 90000 6 mports_i[0]
port 2 nsew signal input
rlabel metal2 s 40314 89200 40370 90000 6 mports_i[100]
port 3 nsew signal input
rlabel metal2 s 40682 89200 40738 90000 6 mports_i[101]
port 4 nsew signal input
rlabel metal2 s 41050 89200 41106 90000 6 mports_i[102]
port 5 nsew signal input
rlabel metal2 s 41418 89200 41474 90000 6 mports_i[103]
port 6 nsew signal input
rlabel metal2 s 41786 89200 41842 90000 6 mports_i[104]
port 7 nsew signal input
rlabel metal2 s 42154 89200 42210 90000 6 mports_i[105]
port 8 nsew signal input
rlabel metal2 s 42522 89200 42578 90000 6 mports_i[106]
port 9 nsew signal input
rlabel metal2 s 42890 89200 42946 90000 6 mports_i[107]
port 10 nsew signal input
rlabel metal2 s 43258 89200 43314 90000 6 mports_i[108]
port 11 nsew signal input
rlabel metal2 s 43626 89200 43682 90000 6 mports_i[109]
port 12 nsew signal input
rlabel metal2 s 7194 89200 7250 90000 6 mports_i[10]
port 13 nsew signal input
rlabel metal2 s 43994 89200 44050 90000 6 mports_i[110]
port 14 nsew signal input
rlabel metal2 s 44362 89200 44418 90000 6 mports_i[111]
port 15 nsew signal input
rlabel metal2 s 44730 89200 44786 90000 6 mports_i[112]
port 16 nsew signal input
rlabel metal2 s 45098 89200 45154 90000 6 mports_i[113]
port 17 nsew signal input
rlabel metal2 s 45466 89200 45522 90000 6 mports_i[114]
port 18 nsew signal input
rlabel metal2 s 45834 89200 45890 90000 6 mports_i[115]
port 19 nsew signal input
rlabel metal2 s 46202 89200 46258 90000 6 mports_i[116]
port 20 nsew signal input
rlabel metal2 s 46570 89200 46626 90000 6 mports_i[117]
port 21 nsew signal input
rlabel metal2 s 46938 89200 46994 90000 6 mports_i[118]
port 22 nsew signal input
rlabel metal2 s 47306 89200 47362 90000 6 mports_i[119]
port 23 nsew signal input
rlabel metal2 s 7562 89200 7618 90000 6 mports_i[11]
port 24 nsew signal input
rlabel metal2 s 47674 89200 47730 90000 6 mports_i[120]
port 25 nsew signal input
rlabel metal2 s 48042 89200 48098 90000 6 mports_i[121]
port 26 nsew signal input
rlabel metal2 s 48410 89200 48466 90000 6 mports_i[122]
port 27 nsew signal input
rlabel metal2 s 48778 89200 48834 90000 6 mports_i[123]
port 28 nsew signal input
rlabel metal2 s 49146 89200 49202 90000 6 mports_i[124]
port 29 nsew signal input
rlabel metal2 s 49514 89200 49570 90000 6 mports_i[125]
port 30 nsew signal input
rlabel metal2 s 49882 89200 49938 90000 6 mports_i[126]
port 31 nsew signal input
rlabel metal2 s 50250 89200 50306 90000 6 mports_i[127]
port 32 nsew signal input
rlabel metal2 s 50618 89200 50674 90000 6 mports_i[128]
port 33 nsew signal input
rlabel metal2 s 50986 89200 51042 90000 6 mports_i[129]
port 34 nsew signal input
rlabel metal2 s 7930 89200 7986 90000 6 mports_i[12]
port 35 nsew signal input
rlabel metal2 s 51354 89200 51410 90000 6 mports_i[130]
port 36 nsew signal input
rlabel metal2 s 51722 89200 51778 90000 6 mports_i[131]
port 37 nsew signal input
rlabel metal2 s 52090 89200 52146 90000 6 mports_i[132]
port 38 nsew signal input
rlabel metal2 s 52458 89200 52514 90000 6 mports_i[133]
port 39 nsew signal input
rlabel metal2 s 52826 89200 52882 90000 6 mports_i[134]
port 40 nsew signal input
rlabel metal2 s 53194 89200 53250 90000 6 mports_i[135]
port 41 nsew signal input
rlabel metal2 s 53562 89200 53618 90000 6 mports_i[136]
port 42 nsew signal input
rlabel metal2 s 53930 89200 53986 90000 6 mports_i[137]
port 43 nsew signal input
rlabel metal2 s 54298 89200 54354 90000 6 mports_i[138]
port 44 nsew signal input
rlabel metal2 s 54666 89200 54722 90000 6 mports_i[139]
port 45 nsew signal input
rlabel metal2 s 8298 89200 8354 90000 6 mports_i[13]
port 46 nsew signal input
rlabel metal2 s 55034 89200 55090 90000 6 mports_i[140]
port 47 nsew signal input
rlabel metal2 s 55402 89200 55458 90000 6 mports_i[141]
port 48 nsew signal input
rlabel metal2 s 55770 89200 55826 90000 6 mports_i[142]
port 49 nsew signal input
rlabel metal2 s 56138 89200 56194 90000 6 mports_i[143]
port 50 nsew signal input
rlabel metal2 s 56506 89200 56562 90000 6 mports_i[144]
port 51 nsew signal input
rlabel metal2 s 56874 89200 56930 90000 6 mports_i[145]
port 52 nsew signal input
rlabel metal2 s 57242 89200 57298 90000 6 mports_i[146]
port 53 nsew signal input
rlabel metal2 s 57610 89200 57666 90000 6 mports_i[147]
port 54 nsew signal input
rlabel metal2 s 57978 89200 58034 90000 6 mports_i[148]
port 55 nsew signal input
rlabel metal2 s 58346 89200 58402 90000 6 mports_i[149]
port 56 nsew signal input
rlabel metal2 s 8666 89200 8722 90000 6 mports_i[14]
port 57 nsew signal input
rlabel metal2 s 58714 89200 58770 90000 6 mports_i[150]
port 58 nsew signal input
rlabel metal2 s 59082 89200 59138 90000 6 mports_i[151]
port 59 nsew signal input
rlabel metal2 s 59450 89200 59506 90000 6 mports_i[152]
port 60 nsew signal input
rlabel metal2 s 59818 89200 59874 90000 6 mports_i[153]
port 61 nsew signal input
rlabel metal2 s 60186 89200 60242 90000 6 mports_i[154]
port 62 nsew signal input
rlabel metal2 s 60554 89200 60610 90000 6 mports_i[155]
port 63 nsew signal input
rlabel metal2 s 60922 89200 60978 90000 6 mports_i[156]
port 64 nsew signal input
rlabel metal2 s 61290 89200 61346 90000 6 mports_i[157]
port 65 nsew signal input
rlabel metal2 s 61658 89200 61714 90000 6 mports_i[158]
port 66 nsew signal input
rlabel metal2 s 62026 89200 62082 90000 6 mports_i[159]
port 67 nsew signal input
rlabel metal2 s 9034 89200 9090 90000 6 mports_i[15]
port 68 nsew signal input
rlabel metal2 s 62394 89200 62450 90000 6 mports_i[160]
port 69 nsew signal input
rlabel metal2 s 62762 89200 62818 90000 6 mports_i[161]
port 70 nsew signal input
rlabel metal2 s 63130 89200 63186 90000 6 mports_i[162]
port 71 nsew signal input
rlabel metal2 s 63498 89200 63554 90000 6 mports_i[163]
port 72 nsew signal input
rlabel metal2 s 63866 89200 63922 90000 6 mports_i[164]
port 73 nsew signal input
rlabel metal2 s 64234 89200 64290 90000 6 mports_i[165]
port 74 nsew signal input
rlabel metal2 s 64602 89200 64658 90000 6 mports_i[166]
port 75 nsew signal input
rlabel metal2 s 64970 89200 65026 90000 6 mports_i[167]
port 76 nsew signal input
rlabel metal2 s 65338 89200 65394 90000 6 mports_i[168]
port 77 nsew signal input
rlabel metal2 s 65706 89200 65762 90000 6 mports_i[169]
port 78 nsew signal input
rlabel metal2 s 9402 89200 9458 90000 6 mports_i[16]
port 79 nsew signal input
rlabel metal2 s 66074 89200 66130 90000 6 mports_i[170]
port 80 nsew signal input
rlabel metal2 s 66442 89200 66498 90000 6 mports_i[171]
port 81 nsew signal input
rlabel metal2 s 66810 89200 66866 90000 6 mports_i[172]
port 82 nsew signal input
rlabel metal2 s 67178 89200 67234 90000 6 mports_i[173]
port 83 nsew signal input
rlabel metal2 s 67546 89200 67602 90000 6 mports_i[174]
port 84 nsew signal input
rlabel metal2 s 67914 89200 67970 90000 6 mports_i[175]
port 85 nsew signal input
rlabel metal2 s 68282 89200 68338 90000 6 mports_i[176]
port 86 nsew signal input
rlabel metal2 s 68650 89200 68706 90000 6 mports_i[177]
port 87 nsew signal input
rlabel metal2 s 69018 89200 69074 90000 6 mports_i[178]
port 88 nsew signal input
rlabel metal2 s 69386 89200 69442 90000 6 mports_i[179]
port 89 nsew signal input
rlabel metal2 s 9770 89200 9826 90000 6 mports_i[17]
port 90 nsew signal input
rlabel metal2 s 69754 89200 69810 90000 6 mports_i[180]
port 91 nsew signal input
rlabel metal2 s 70122 89200 70178 90000 6 mports_i[181]
port 92 nsew signal input
rlabel metal2 s 70490 89200 70546 90000 6 mports_i[182]
port 93 nsew signal input
rlabel metal2 s 70858 89200 70914 90000 6 mports_i[183]
port 94 nsew signal input
rlabel metal2 s 71226 89200 71282 90000 6 mports_i[184]
port 95 nsew signal input
rlabel metal2 s 71594 89200 71650 90000 6 mports_i[185]
port 96 nsew signal input
rlabel metal2 s 71962 89200 72018 90000 6 mports_i[186]
port 97 nsew signal input
rlabel metal2 s 72330 89200 72386 90000 6 mports_i[187]
port 98 nsew signal input
rlabel metal2 s 72698 89200 72754 90000 6 mports_i[188]
port 99 nsew signal input
rlabel metal2 s 73066 89200 73122 90000 6 mports_i[189]
port 100 nsew signal input
rlabel metal2 s 10138 89200 10194 90000 6 mports_i[18]
port 101 nsew signal input
rlabel metal2 s 73434 89200 73490 90000 6 mports_i[190]
port 102 nsew signal input
rlabel metal2 s 73802 89200 73858 90000 6 mports_i[191]
port 103 nsew signal input
rlabel metal2 s 74170 89200 74226 90000 6 mports_i[192]
port 104 nsew signal input
rlabel metal2 s 74538 89200 74594 90000 6 mports_i[193]
port 105 nsew signal input
rlabel metal2 s 74906 89200 74962 90000 6 mports_i[194]
port 106 nsew signal input
rlabel metal2 s 75274 89200 75330 90000 6 mports_i[195]
port 107 nsew signal input
rlabel metal2 s 75642 89200 75698 90000 6 mports_i[196]
port 108 nsew signal input
rlabel metal2 s 76010 89200 76066 90000 6 mports_i[197]
port 109 nsew signal input
rlabel metal2 s 76378 89200 76434 90000 6 mports_i[198]
port 110 nsew signal input
rlabel metal2 s 76746 89200 76802 90000 6 mports_i[199]
port 111 nsew signal input
rlabel metal2 s 10506 89200 10562 90000 6 mports_i[19]
port 112 nsew signal input
rlabel metal2 s 3882 89200 3938 90000 6 mports_i[1]
port 113 nsew signal input
rlabel metal2 s 77114 89200 77170 90000 6 mports_i[200]
port 114 nsew signal input
rlabel metal2 s 77482 89200 77538 90000 6 mports_i[201]
port 115 nsew signal input
rlabel metal2 s 77850 89200 77906 90000 6 mports_i[202]
port 116 nsew signal input
rlabel metal2 s 78218 89200 78274 90000 6 mports_i[203]
port 117 nsew signal input
rlabel metal2 s 78586 89200 78642 90000 6 mports_i[204]
port 118 nsew signal input
rlabel metal2 s 78954 89200 79010 90000 6 mports_i[205]
port 119 nsew signal input
rlabel metal2 s 79322 89200 79378 90000 6 mports_i[206]
port 120 nsew signal input
rlabel metal2 s 79690 89200 79746 90000 6 mports_i[207]
port 121 nsew signal input
rlabel metal2 s 80058 89200 80114 90000 6 mports_i[208]
port 122 nsew signal input
rlabel metal2 s 80426 89200 80482 90000 6 mports_i[209]
port 123 nsew signal input
rlabel metal2 s 10874 89200 10930 90000 6 mports_i[20]
port 124 nsew signal input
rlabel metal2 s 80794 89200 80850 90000 6 mports_i[210]
port 125 nsew signal input
rlabel metal2 s 81162 89200 81218 90000 6 mports_i[211]
port 126 nsew signal input
rlabel metal2 s 81530 89200 81586 90000 6 mports_i[212]
port 127 nsew signal input
rlabel metal2 s 81898 89200 81954 90000 6 mports_i[213]
port 128 nsew signal input
rlabel metal2 s 82266 89200 82322 90000 6 mports_i[214]
port 129 nsew signal input
rlabel metal2 s 82634 89200 82690 90000 6 mports_i[215]
port 130 nsew signal input
rlabel metal2 s 83002 89200 83058 90000 6 mports_i[216]
port 131 nsew signal input
rlabel metal2 s 83370 89200 83426 90000 6 mports_i[217]
port 132 nsew signal input
rlabel metal2 s 83738 89200 83794 90000 6 mports_i[218]
port 133 nsew signal input
rlabel metal2 s 84106 89200 84162 90000 6 mports_i[219]
port 134 nsew signal input
rlabel metal2 s 11242 89200 11298 90000 6 mports_i[21]
port 135 nsew signal input
rlabel metal2 s 84474 89200 84530 90000 6 mports_i[220]
port 136 nsew signal input
rlabel metal2 s 84842 89200 84898 90000 6 mports_i[221]
port 137 nsew signal input
rlabel metal2 s 85210 89200 85266 90000 6 mports_i[222]
port 138 nsew signal input
rlabel metal2 s 85578 89200 85634 90000 6 mports_i[223]
port 139 nsew signal input
rlabel metal2 s 85946 89200 86002 90000 6 mports_i[224]
port 140 nsew signal input
rlabel metal2 s 86314 89200 86370 90000 6 mports_i[225]
port 141 nsew signal input
rlabel metal2 s 86682 89200 86738 90000 6 mports_i[226]
port 142 nsew signal input
rlabel metal2 s 87050 89200 87106 90000 6 mports_i[227]
port 143 nsew signal input
rlabel metal2 s 11610 89200 11666 90000 6 mports_i[22]
port 144 nsew signal input
rlabel metal2 s 11978 89200 12034 90000 6 mports_i[23]
port 145 nsew signal input
rlabel metal2 s 12346 89200 12402 90000 6 mports_i[24]
port 146 nsew signal input
rlabel metal2 s 12714 89200 12770 90000 6 mports_i[25]
port 147 nsew signal input
rlabel metal2 s 13082 89200 13138 90000 6 mports_i[26]
port 148 nsew signal input
rlabel metal2 s 13450 89200 13506 90000 6 mports_i[27]
port 149 nsew signal input
rlabel metal2 s 13818 89200 13874 90000 6 mports_i[28]
port 150 nsew signal input
rlabel metal2 s 14186 89200 14242 90000 6 mports_i[29]
port 151 nsew signal input
rlabel metal2 s 4250 89200 4306 90000 6 mports_i[2]
port 152 nsew signal input
rlabel metal2 s 14554 89200 14610 90000 6 mports_i[30]
port 153 nsew signal input
rlabel metal2 s 14922 89200 14978 90000 6 mports_i[31]
port 154 nsew signal input
rlabel metal2 s 15290 89200 15346 90000 6 mports_i[32]
port 155 nsew signal input
rlabel metal2 s 15658 89200 15714 90000 6 mports_i[33]
port 156 nsew signal input
rlabel metal2 s 16026 89200 16082 90000 6 mports_i[34]
port 157 nsew signal input
rlabel metal2 s 16394 89200 16450 90000 6 mports_i[35]
port 158 nsew signal input
rlabel metal2 s 16762 89200 16818 90000 6 mports_i[36]
port 159 nsew signal input
rlabel metal2 s 17130 89200 17186 90000 6 mports_i[37]
port 160 nsew signal input
rlabel metal2 s 17498 89200 17554 90000 6 mports_i[38]
port 161 nsew signal input
rlabel metal2 s 17866 89200 17922 90000 6 mports_i[39]
port 162 nsew signal input
rlabel metal2 s 4618 89200 4674 90000 6 mports_i[3]
port 163 nsew signal input
rlabel metal2 s 18234 89200 18290 90000 6 mports_i[40]
port 164 nsew signal input
rlabel metal2 s 18602 89200 18658 90000 6 mports_i[41]
port 165 nsew signal input
rlabel metal2 s 18970 89200 19026 90000 6 mports_i[42]
port 166 nsew signal input
rlabel metal2 s 19338 89200 19394 90000 6 mports_i[43]
port 167 nsew signal input
rlabel metal2 s 19706 89200 19762 90000 6 mports_i[44]
port 168 nsew signal input
rlabel metal2 s 20074 89200 20130 90000 6 mports_i[45]
port 169 nsew signal input
rlabel metal2 s 20442 89200 20498 90000 6 mports_i[46]
port 170 nsew signal input
rlabel metal2 s 20810 89200 20866 90000 6 mports_i[47]
port 171 nsew signal input
rlabel metal2 s 21178 89200 21234 90000 6 mports_i[48]
port 172 nsew signal input
rlabel metal2 s 21546 89200 21602 90000 6 mports_i[49]
port 173 nsew signal input
rlabel metal2 s 4986 89200 5042 90000 6 mports_i[4]
port 174 nsew signal input
rlabel metal2 s 21914 89200 21970 90000 6 mports_i[50]
port 175 nsew signal input
rlabel metal2 s 22282 89200 22338 90000 6 mports_i[51]
port 176 nsew signal input
rlabel metal2 s 22650 89200 22706 90000 6 mports_i[52]
port 177 nsew signal input
rlabel metal2 s 23018 89200 23074 90000 6 mports_i[53]
port 178 nsew signal input
rlabel metal2 s 23386 89200 23442 90000 6 mports_i[54]
port 179 nsew signal input
rlabel metal2 s 23754 89200 23810 90000 6 mports_i[55]
port 180 nsew signal input
rlabel metal2 s 24122 89200 24178 90000 6 mports_i[56]
port 181 nsew signal input
rlabel metal2 s 24490 89200 24546 90000 6 mports_i[57]
port 182 nsew signal input
rlabel metal2 s 24858 89200 24914 90000 6 mports_i[58]
port 183 nsew signal input
rlabel metal2 s 25226 89200 25282 90000 6 mports_i[59]
port 184 nsew signal input
rlabel metal2 s 5354 89200 5410 90000 6 mports_i[5]
port 185 nsew signal input
rlabel metal2 s 25594 89200 25650 90000 6 mports_i[60]
port 186 nsew signal input
rlabel metal2 s 25962 89200 26018 90000 6 mports_i[61]
port 187 nsew signal input
rlabel metal2 s 26330 89200 26386 90000 6 mports_i[62]
port 188 nsew signal input
rlabel metal2 s 26698 89200 26754 90000 6 mports_i[63]
port 189 nsew signal input
rlabel metal2 s 27066 89200 27122 90000 6 mports_i[64]
port 190 nsew signal input
rlabel metal2 s 27434 89200 27490 90000 6 mports_i[65]
port 191 nsew signal input
rlabel metal2 s 27802 89200 27858 90000 6 mports_i[66]
port 192 nsew signal input
rlabel metal2 s 28170 89200 28226 90000 6 mports_i[67]
port 193 nsew signal input
rlabel metal2 s 28538 89200 28594 90000 6 mports_i[68]
port 194 nsew signal input
rlabel metal2 s 28906 89200 28962 90000 6 mports_i[69]
port 195 nsew signal input
rlabel metal2 s 5722 89200 5778 90000 6 mports_i[6]
port 196 nsew signal input
rlabel metal2 s 29274 89200 29330 90000 6 mports_i[70]
port 197 nsew signal input
rlabel metal2 s 29642 89200 29698 90000 6 mports_i[71]
port 198 nsew signal input
rlabel metal2 s 30010 89200 30066 90000 6 mports_i[72]
port 199 nsew signal input
rlabel metal2 s 30378 89200 30434 90000 6 mports_i[73]
port 200 nsew signal input
rlabel metal2 s 30746 89200 30802 90000 6 mports_i[74]
port 201 nsew signal input
rlabel metal2 s 31114 89200 31170 90000 6 mports_i[75]
port 202 nsew signal input
rlabel metal2 s 31482 89200 31538 90000 6 mports_i[76]
port 203 nsew signal input
rlabel metal2 s 31850 89200 31906 90000 6 mports_i[77]
port 204 nsew signal input
rlabel metal2 s 32218 89200 32274 90000 6 mports_i[78]
port 205 nsew signal input
rlabel metal2 s 32586 89200 32642 90000 6 mports_i[79]
port 206 nsew signal input
rlabel metal2 s 6090 89200 6146 90000 6 mports_i[7]
port 207 nsew signal input
rlabel metal2 s 32954 89200 33010 90000 6 mports_i[80]
port 208 nsew signal input
rlabel metal2 s 33322 89200 33378 90000 6 mports_i[81]
port 209 nsew signal input
rlabel metal2 s 33690 89200 33746 90000 6 mports_i[82]
port 210 nsew signal input
rlabel metal2 s 34058 89200 34114 90000 6 mports_i[83]
port 211 nsew signal input
rlabel metal2 s 34426 89200 34482 90000 6 mports_i[84]
port 212 nsew signal input
rlabel metal2 s 34794 89200 34850 90000 6 mports_i[85]
port 213 nsew signal input
rlabel metal2 s 35162 89200 35218 90000 6 mports_i[86]
port 214 nsew signal input
rlabel metal2 s 35530 89200 35586 90000 6 mports_i[87]
port 215 nsew signal input
rlabel metal2 s 35898 89200 35954 90000 6 mports_i[88]
port 216 nsew signal input
rlabel metal2 s 36266 89200 36322 90000 6 mports_i[89]
port 217 nsew signal input
rlabel metal2 s 6458 89200 6514 90000 6 mports_i[8]
port 218 nsew signal input
rlabel metal2 s 36634 89200 36690 90000 6 mports_i[90]
port 219 nsew signal input
rlabel metal2 s 37002 89200 37058 90000 6 mports_i[91]
port 220 nsew signal input
rlabel metal2 s 37370 89200 37426 90000 6 mports_i[92]
port 221 nsew signal input
rlabel metal2 s 37738 89200 37794 90000 6 mports_i[93]
port 222 nsew signal input
rlabel metal2 s 38106 89200 38162 90000 6 mports_i[94]
port 223 nsew signal input
rlabel metal2 s 38474 89200 38530 90000 6 mports_i[95]
port 224 nsew signal input
rlabel metal2 s 38842 89200 38898 90000 6 mports_i[96]
port 225 nsew signal input
rlabel metal2 s 39210 89200 39266 90000 6 mports_i[97]
port 226 nsew signal input
rlabel metal2 s 39578 89200 39634 90000 6 mports_i[98]
port 227 nsew signal input
rlabel metal2 s 39946 89200 40002 90000 6 mports_i[99]
port 228 nsew signal input
rlabel metal2 s 6826 89200 6882 90000 6 mports_i[9]
port 229 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 mports_o[0]
port 230 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 mports_o[100]
port 231 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 mports_o[101]
port 232 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 mports_o[102]
port 233 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 mports_o[103]
port 234 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 mports_o[104]
port 235 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 mports_o[105]
port 236 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 mports_o[106]
port 237 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 mports_o[107]
port 238 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 mports_o[108]
port 239 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 mports_o[109]
port 240 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 mports_o[10]
port 241 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 mports_o[110]
port 242 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 mports_o[111]
port 243 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 mports_o[112]
port 244 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 mports_o[113]
port 245 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 mports_o[114]
port 246 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 mports_o[115]
port 247 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 mports_o[116]
port 248 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 mports_o[117]
port 249 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 mports_o[118]
port 250 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 mports_o[119]
port 251 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 mports_o[11]
port 252 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 mports_o[120]
port 253 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 mports_o[121]
port 254 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 mports_o[122]
port 255 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 mports_o[123]
port 256 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 mports_o[124]
port 257 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 mports_o[125]
port 258 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 mports_o[126]
port 259 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 mports_o[127]
port 260 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 mports_o[128]
port 261 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 mports_o[129]
port 262 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 mports_o[12]
port 263 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 mports_o[130]
port 264 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 mports_o[131]
port 265 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 mports_o[132]
port 266 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 mports_o[133]
port 267 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 mports_o[134]
port 268 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 mports_o[135]
port 269 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 mports_o[13]
port 270 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 mports_o[14]
port 271 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 mports_o[15]
port 272 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 mports_o[16]
port 273 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 mports_o[17]
port 274 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 mports_o[18]
port 275 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 mports_o[19]
port 276 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 mports_o[1]
port 277 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 mports_o[20]
port 278 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 mports_o[21]
port 279 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 mports_o[22]
port 280 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 mports_o[23]
port 281 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 mports_o[24]
port 282 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 mports_o[25]
port 283 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 mports_o[26]
port 284 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 mports_o[27]
port 285 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 mports_o[28]
port 286 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 mports_o[29]
port 287 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 mports_o[2]
port 288 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 mports_o[30]
port 289 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 mports_o[31]
port 290 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 mports_o[32]
port 291 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 mports_o[33]
port 292 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 mports_o[34]
port 293 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 mports_o[35]
port 294 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 mports_o[36]
port 295 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 mports_o[37]
port 296 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 mports_o[38]
port 297 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 mports_o[39]
port 298 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 mports_o[3]
port 299 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 mports_o[40]
port 300 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 mports_o[41]
port 301 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 mports_o[42]
port 302 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 mports_o[43]
port 303 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 mports_o[44]
port 304 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 mports_o[45]
port 305 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 mports_o[46]
port 306 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 mports_o[47]
port 307 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 mports_o[48]
port 308 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 mports_o[49]
port 309 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 mports_o[4]
port 310 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 mports_o[50]
port 311 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 mports_o[51]
port 312 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 mports_o[52]
port 313 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 mports_o[53]
port 314 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 mports_o[54]
port 315 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 mports_o[55]
port 316 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 mports_o[56]
port 317 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 mports_o[57]
port 318 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 mports_o[58]
port 319 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 mports_o[59]
port 320 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 mports_o[5]
port 321 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 mports_o[60]
port 322 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 mports_o[61]
port 323 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 mports_o[62]
port 324 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 mports_o[63]
port 325 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 mports_o[64]
port 326 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 mports_o[65]
port 327 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 mports_o[66]
port 328 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 mports_o[67]
port 329 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 mports_o[68]
port 330 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 mports_o[69]
port 331 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 mports_o[6]
port 332 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 mports_o[70]
port 333 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 mports_o[71]
port 334 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 mports_o[72]
port 335 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 mports_o[73]
port 336 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 mports_o[74]
port 337 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 mports_o[75]
port 338 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 mports_o[76]
port 339 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 mports_o[77]
port 340 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 mports_o[78]
port 341 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 mports_o[79]
port 342 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 mports_o[7]
port 343 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 mports_o[80]
port 344 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 mports_o[81]
port 345 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 mports_o[82]
port 346 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 mports_o[83]
port 347 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 mports_o[84]
port 348 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 mports_o[85]
port 349 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 mports_o[86]
port 350 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 mports_o[87]
port 351 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 mports_o[88]
port 352 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 mports_o[89]
port 353 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 mports_o[8]
port 354 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 mports_o[90]
port 355 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 mports_o[91]
port 356 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 mports_o[92]
port 357 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 mports_o[93]
port 358 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 mports_o[94]
port 359 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 mports_o[95]
port 360 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 mports_o[96]
port 361 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 mports_o[97]
port 362 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 mports_o[98]
port 363 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 mports_o[99]
port 364 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 mports_o[9]
port 365 nsew signal output
rlabel metal2 s 3146 89200 3202 90000 6 nrst_i
port 366 nsew signal input
rlabel metal3 s 89200 8168 90000 8288 6 sports_i[0]
port 367 nsew signal input
rlabel metal3 s 89200 62568 90000 62688 6 sports_i[100]
port 368 nsew signal input
rlabel metal3 s 89200 63112 90000 63232 6 sports_i[101]
port 369 nsew signal input
rlabel metal3 s 89200 63656 90000 63776 6 sports_i[102]
port 370 nsew signal input
rlabel metal3 s 89200 64200 90000 64320 6 sports_i[103]
port 371 nsew signal input
rlabel metal3 s 89200 64744 90000 64864 6 sports_i[104]
port 372 nsew signal input
rlabel metal3 s 89200 65288 90000 65408 6 sports_i[105]
port 373 nsew signal input
rlabel metal3 s 89200 65832 90000 65952 6 sports_i[106]
port 374 nsew signal input
rlabel metal3 s 89200 66376 90000 66496 6 sports_i[107]
port 375 nsew signal input
rlabel metal3 s 89200 66920 90000 67040 6 sports_i[108]
port 376 nsew signal input
rlabel metal3 s 89200 67464 90000 67584 6 sports_i[109]
port 377 nsew signal input
rlabel metal3 s 89200 13608 90000 13728 6 sports_i[10]
port 378 nsew signal input
rlabel metal3 s 89200 68008 90000 68128 6 sports_i[110]
port 379 nsew signal input
rlabel metal3 s 89200 68552 90000 68672 6 sports_i[111]
port 380 nsew signal input
rlabel metal3 s 89200 69096 90000 69216 6 sports_i[112]
port 381 nsew signal input
rlabel metal3 s 89200 69640 90000 69760 6 sports_i[113]
port 382 nsew signal input
rlabel metal3 s 89200 70184 90000 70304 6 sports_i[114]
port 383 nsew signal input
rlabel metal3 s 89200 70728 90000 70848 6 sports_i[115]
port 384 nsew signal input
rlabel metal3 s 89200 71272 90000 71392 6 sports_i[116]
port 385 nsew signal input
rlabel metal3 s 89200 71816 90000 71936 6 sports_i[117]
port 386 nsew signal input
rlabel metal3 s 89200 72360 90000 72480 6 sports_i[118]
port 387 nsew signal input
rlabel metal3 s 89200 72904 90000 73024 6 sports_i[119]
port 388 nsew signal input
rlabel metal3 s 89200 14152 90000 14272 6 sports_i[11]
port 389 nsew signal input
rlabel metal3 s 89200 73448 90000 73568 6 sports_i[120]
port 390 nsew signal input
rlabel metal3 s 89200 73992 90000 74112 6 sports_i[121]
port 391 nsew signal input
rlabel metal3 s 89200 74536 90000 74656 6 sports_i[122]
port 392 nsew signal input
rlabel metal3 s 89200 75080 90000 75200 6 sports_i[123]
port 393 nsew signal input
rlabel metal3 s 89200 75624 90000 75744 6 sports_i[124]
port 394 nsew signal input
rlabel metal3 s 89200 76168 90000 76288 6 sports_i[125]
port 395 nsew signal input
rlabel metal3 s 89200 76712 90000 76832 6 sports_i[126]
port 396 nsew signal input
rlabel metal3 s 89200 77256 90000 77376 6 sports_i[127]
port 397 nsew signal input
rlabel metal3 s 89200 77800 90000 77920 6 sports_i[128]
port 398 nsew signal input
rlabel metal3 s 89200 78344 90000 78464 6 sports_i[129]
port 399 nsew signal input
rlabel metal3 s 89200 14696 90000 14816 6 sports_i[12]
port 400 nsew signal input
rlabel metal3 s 89200 78888 90000 79008 6 sports_i[130]
port 401 nsew signal input
rlabel metal3 s 89200 79432 90000 79552 6 sports_i[131]
port 402 nsew signal input
rlabel metal3 s 89200 79976 90000 80096 6 sports_i[132]
port 403 nsew signal input
rlabel metal3 s 89200 80520 90000 80640 6 sports_i[133]
port 404 nsew signal input
rlabel metal3 s 89200 81064 90000 81184 6 sports_i[134]
port 405 nsew signal input
rlabel metal3 s 89200 81608 90000 81728 6 sports_i[135]
port 406 nsew signal input
rlabel metal3 s 89200 15240 90000 15360 6 sports_i[13]
port 407 nsew signal input
rlabel metal3 s 89200 15784 90000 15904 6 sports_i[14]
port 408 nsew signal input
rlabel metal3 s 89200 16328 90000 16448 6 sports_i[15]
port 409 nsew signal input
rlabel metal3 s 89200 16872 90000 16992 6 sports_i[16]
port 410 nsew signal input
rlabel metal3 s 89200 17416 90000 17536 6 sports_i[17]
port 411 nsew signal input
rlabel metal3 s 89200 17960 90000 18080 6 sports_i[18]
port 412 nsew signal input
rlabel metal3 s 89200 18504 90000 18624 6 sports_i[19]
port 413 nsew signal input
rlabel metal3 s 89200 8712 90000 8832 6 sports_i[1]
port 414 nsew signal input
rlabel metal3 s 89200 19048 90000 19168 6 sports_i[20]
port 415 nsew signal input
rlabel metal3 s 89200 19592 90000 19712 6 sports_i[21]
port 416 nsew signal input
rlabel metal3 s 89200 20136 90000 20256 6 sports_i[22]
port 417 nsew signal input
rlabel metal3 s 89200 20680 90000 20800 6 sports_i[23]
port 418 nsew signal input
rlabel metal3 s 89200 21224 90000 21344 6 sports_i[24]
port 419 nsew signal input
rlabel metal3 s 89200 21768 90000 21888 6 sports_i[25]
port 420 nsew signal input
rlabel metal3 s 89200 22312 90000 22432 6 sports_i[26]
port 421 nsew signal input
rlabel metal3 s 89200 22856 90000 22976 6 sports_i[27]
port 422 nsew signal input
rlabel metal3 s 89200 23400 90000 23520 6 sports_i[28]
port 423 nsew signal input
rlabel metal3 s 89200 23944 90000 24064 6 sports_i[29]
port 424 nsew signal input
rlabel metal3 s 89200 9256 90000 9376 6 sports_i[2]
port 425 nsew signal input
rlabel metal3 s 89200 24488 90000 24608 6 sports_i[30]
port 426 nsew signal input
rlabel metal3 s 89200 25032 90000 25152 6 sports_i[31]
port 427 nsew signal input
rlabel metal3 s 89200 25576 90000 25696 6 sports_i[32]
port 428 nsew signal input
rlabel metal3 s 89200 26120 90000 26240 6 sports_i[33]
port 429 nsew signal input
rlabel metal3 s 89200 26664 90000 26784 6 sports_i[34]
port 430 nsew signal input
rlabel metal3 s 89200 27208 90000 27328 6 sports_i[35]
port 431 nsew signal input
rlabel metal3 s 89200 27752 90000 27872 6 sports_i[36]
port 432 nsew signal input
rlabel metal3 s 89200 28296 90000 28416 6 sports_i[37]
port 433 nsew signal input
rlabel metal3 s 89200 28840 90000 28960 6 sports_i[38]
port 434 nsew signal input
rlabel metal3 s 89200 29384 90000 29504 6 sports_i[39]
port 435 nsew signal input
rlabel metal3 s 89200 9800 90000 9920 6 sports_i[3]
port 436 nsew signal input
rlabel metal3 s 89200 29928 90000 30048 6 sports_i[40]
port 437 nsew signal input
rlabel metal3 s 89200 30472 90000 30592 6 sports_i[41]
port 438 nsew signal input
rlabel metal3 s 89200 31016 90000 31136 6 sports_i[42]
port 439 nsew signal input
rlabel metal3 s 89200 31560 90000 31680 6 sports_i[43]
port 440 nsew signal input
rlabel metal3 s 89200 32104 90000 32224 6 sports_i[44]
port 441 nsew signal input
rlabel metal3 s 89200 32648 90000 32768 6 sports_i[45]
port 442 nsew signal input
rlabel metal3 s 89200 33192 90000 33312 6 sports_i[46]
port 443 nsew signal input
rlabel metal3 s 89200 33736 90000 33856 6 sports_i[47]
port 444 nsew signal input
rlabel metal3 s 89200 34280 90000 34400 6 sports_i[48]
port 445 nsew signal input
rlabel metal3 s 89200 34824 90000 34944 6 sports_i[49]
port 446 nsew signal input
rlabel metal3 s 89200 10344 90000 10464 6 sports_i[4]
port 447 nsew signal input
rlabel metal3 s 89200 35368 90000 35488 6 sports_i[50]
port 448 nsew signal input
rlabel metal3 s 89200 35912 90000 36032 6 sports_i[51]
port 449 nsew signal input
rlabel metal3 s 89200 36456 90000 36576 6 sports_i[52]
port 450 nsew signal input
rlabel metal3 s 89200 37000 90000 37120 6 sports_i[53]
port 451 nsew signal input
rlabel metal3 s 89200 37544 90000 37664 6 sports_i[54]
port 452 nsew signal input
rlabel metal3 s 89200 38088 90000 38208 6 sports_i[55]
port 453 nsew signal input
rlabel metal3 s 89200 38632 90000 38752 6 sports_i[56]
port 454 nsew signal input
rlabel metal3 s 89200 39176 90000 39296 6 sports_i[57]
port 455 nsew signal input
rlabel metal3 s 89200 39720 90000 39840 6 sports_i[58]
port 456 nsew signal input
rlabel metal3 s 89200 40264 90000 40384 6 sports_i[59]
port 457 nsew signal input
rlabel metal3 s 89200 10888 90000 11008 6 sports_i[5]
port 458 nsew signal input
rlabel metal3 s 89200 40808 90000 40928 6 sports_i[60]
port 459 nsew signal input
rlabel metal3 s 89200 41352 90000 41472 6 sports_i[61]
port 460 nsew signal input
rlabel metal3 s 89200 41896 90000 42016 6 sports_i[62]
port 461 nsew signal input
rlabel metal3 s 89200 42440 90000 42560 6 sports_i[63]
port 462 nsew signal input
rlabel metal3 s 89200 42984 90000 43104 6 sports_i[64]
port 463 nsew signal input
rlabel metal3 s 89200 43528 90000 43648 6 sports_i[65]
port 464 nsew signal input
rlabel metal3 s 89200 44072 90000 44192 6 sports_i[66]
port 465 nsew signal input
rlabel metal3 s 89200 44616 90000 44736 6 sports_i[67]
port 466 nsew signal input
rlabel metal3 s 89200 45160 90000 45280 6 sports_i[68]
port 467 nsew signal input
rlabel metal3 s 89200 45704 90000 45824 6 sports_i[69]
port 468 nsew signal input
rlabel metal3 s 89200 11432 90000 11552 6 sports_i[6]
port 469 nsew signal input
rlabel metal3 s 89200 46248 90000 46368 6 sports_i[70]
port 470 nsew signal input
rlabel metal3 s 89200 46792 90000 46912 6 sports_i[71]
port 471 nsew signal input
rlabel metal3 s 89200 47336 90000 47456 6 sports_i[72]
port 472 nsew signal input
rlabel metal3 s 89200 47880 90000 48000 6 sports_i[73]
port 473 nsew signal input
rlabel metal3 s 89200 48424 90000 48544 6 sports_i[74]
port 474 nsew signal input
rlabel metal3 s 89200 48968 90000 49088 6 sports_i[75]
port 475 nsew signal input
rlabel metal3 s 89200 49512 90000 49632 6 sports_i[76]
port 476 nsew signal input
rlabel metal3 s 89200 50056 90000 50176 6 sports_i[77]
port 477 nsew signal input
rlabel metal3 s 89200 50600 90000 50720 6 sports_i[78]
port 478 nsew signal input
rlabel metal3 s 89200 51144 90000 51264 6 sports_i[79]
port 479 nsew signal input
rlabel metal3 s 89200 11976 90000 12096 6 sports_i[7]
port 480 nsew signal input
rlabel metal3 s 89200 51688 90000 51808 6 sports_i[80]
port 481 nsew signal input
rlabel metal3 s 89200 52232 90000 52352 6 sports_i[81]
port 482 nsew signal input
rlabel metal3 s 89200 52776 90000 52896 6 sports_i[82]
port 483 nsew signal input
rlabel metal3 s 89200 53320 90000 53440 6 sports_i[83]
port 484 nsew signal input
rlabel metal3 s 89200 53864 90000 53984 6 sports_i[84]
port 485 nsew signal input
rlabel metal3 s 89200 54408 90000 54528 6 sports_i[85]
port 486 nsew signal input
rlabel metal3 s 89200 54952 90000 55072 6 sports_i[86]
port 487 nsew signal input
rlabel metal3 s 89200 55496 90000 55616 6 sports_i[87]
port 488 nsew signal input
rlabel metal3 s 89200 56040 90000 56160 6 sports_i[88]
port 489 nsew signal input
rlabel metal3 s 89200 56584 90000 56704 6 sports_i[89]
port 490 nsew signal input
rlabel metal3 s 89200 12520 90000 12640 6 sports_i[8]
port 491 nsew signal input
rlabel metal3 s 89200 57128 90000 57248 6 sports_i[90]
port 492 nsew signal input
rlabel metal3 s 89200 57672 90000 57792 6 sports_i[91]
port 493 nsew signal input
rlabel metal3 s 89200 58216 90000 58336 6 sports_i[92]
port 494 nsew signal input
rlabel metal3 s 89200 58760 90000 58880 6 sports_i[93]
port 495 nsew signal input
rlabel metal3 s 89200 59304 90000 59424 6 sports_i[94]
port 496 nsew signal input
rlabel metal3 s 89200 59848 90000 59968 6 sports_i[95]
port 497 nsew signal input
rlabel metal3 s 89200 60392 90000 60512 6 sports_i[96]
port 498 nsew signal input
rlabel metal3 s 89200 60936 90000 61056 6 sports_i[97]
port 499 nsew signal input
rlabel metal3 s 89200 61480 90000 61600 6 sports_i[98]
port 500 nsew signal input
rlabel metal3 s 89200 62024 90000 62144 6 sports_i[99]
port 501 nsew signal input
rlabel metal3 s 89200 13064 90000 13184 6 sports_i[9]
port 502 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 sports_o[0]
port 503 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 sports_o[100]
port 504 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 sports_o[101]
port 505 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 sports_o[102]
port 506 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 sports_o[103]
port 507 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 sports_o[104]
port 508 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 sports_o[105]
port 509 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 sports_o[106]
port 510 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 sports_o[107]
port 511 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 sports_o[108]
port 512 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 sports_o[109]
port 513 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 sports_o[10]
port 514 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 sports_o[110]
port 515 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 sports_o[111]
port 516 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 sports_o[112]
port 517 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 sports_o[113]
port 518 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 sports_o[114]
port 519 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 sports_o[115]
port 520 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 sports_o[116]
port 521 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 sports_o[117]
port 522 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 sports_o[118]
port 523 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 sports_o[119]
port 524 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 sports_o[11]
port 525 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 sports_o[120]
port 526 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 sports_o[121]
port 527 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 sports_o[122]
port 528 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 sports_o[123]
port 529 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 sports_o[124]
port 530 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 sports_o[125]
port 531 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 sports_o[126]
port 532 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 sports_o[127]
port 533 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 sports_o[128]
port 534 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 sports_o[129]
port 535 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 sports_o[12]
port 536 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 sports_o[130]
port 537 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 sports_o[131]
port 538 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 sports_o[132]
port 539 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 sports_o[133]
port 540 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 sports_o[134]
port 541 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 sports_o[135]
port 542 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 sports_o[136]
port 543 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 sports_o[137]
port 544 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 sports_o[138]
port 545 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 sports_o[139]
port 546 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 sports_o[13]
port 547 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 sports_o[140]
port 548 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 sports_o[141]
port 549 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 sports_o[142]
port 550 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 sports_o[143]
port 551 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 sports_o[144]
port 552 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 sports_o[145]
port 553 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 sports_o[146]
port 554 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 sports_o[147]
port 555 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 sports_o[148]
port 556 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 sports_o[149]
port 557 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 sports_o[14]
port 558 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 sports_o[150]
port 559 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 sports_o[151]
port 560 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 sports_o[152]
port 561 nsew signal output
rlabel metal3 s 0 55496 800 55616 6 sports_o[153]
port 562 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 sports_o[154]
port 563 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 sports_o[155]
port 564 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 sports_o[156]
port 565 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 sports_o[157]
port 566 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 sports_o[158]
port 567 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 sports_o[159]
port 568 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 sports_o[15]
port 569 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 sports_o[160]
port 570 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 sports_o[161]
port 571 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 sports_o[162]
port 572 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 sports_o[163]
port 573 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 sports_o[164]
port 574 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 sports_o[165]
port 575 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 sports_o[166]
port 576 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 sports_o[167]
port 577 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 sports_o[168]
port 578 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 sports_o[169]
port 579 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 sports_o[16]
port 580 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 sports_o[170]
port 581 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 sports_o[171]
port 582 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 sports_o[172]
port 583 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 sports_o[173]
port 584 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 sports_o[174]
port 585 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 sports_o[175]
port 586 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 sports_o[176]
port 587 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 sports_o[177]
port 588 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 sports_o[178]
port 589 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 sports_o[179]
port 590 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 sports_o[17]
port 591 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 sports_o[180]
port 592 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 sports_o[181]
port 593 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 sports_o[182]
port 594 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 sports_o[183]
port 595 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 sports_o[184]
port 596 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 sports_o[185]
port 597 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 sports_o[186]
port 598 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 sports_o[187]
port 599 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 sports_o[188]
port 600 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 sports_o[189]
port 601 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 sports_o[18]
port 602 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 sports_o[190]
port 603 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 sports_o[191]
port 604 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 sports_o[192]
port 605 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 sports_o[193]
port 606 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 sports_o[194]
port 607 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 sports_o[195]
port 608 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 sports_o[196]
port 609 nsew signal output
rlabel metal3 s 0 67464 800 67584 6 sports_o[197]
port 610 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 sports_o[198]
port 611 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 sports_o[199]
port 612 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 sports_o[19]
port 613 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 sports_o[1]
port 614 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 sports_o[200]
port 615 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 sports_o[201]
port 616 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 sports_o[202]
port 617 nsew signal output
rlabel metal3 s 0 69096 800 69216 6 sports_o[203]
port 618 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 sports_o[204]
port 619 nsew signal output
rlabel metal3 s 0 69640 800 69760 6 sports_o[205]
port 620 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 sports_o[206]
port 621 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 sports_o[207]
port 622 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 sports_o[208]
port 623 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 sports_o[209]
port 624 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 sports_o[20]
port 625 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 sports_o[210]
port 626 nsew signal output
rlabel metal3 s 0 71272 800 71392 6 sports_o[211]
port 627 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 sports_o[212]
port 628 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 sports_o[213]
port 629 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 sports_o[214]
port 630 nsew signal output
rlabel metal3 s 0 72360 800 72480 6 sports_o[215]
port 631 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 sports_o[216]
port 632 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 sports_o[217]
port 633 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 sports_o[218]
port 634 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 sports_o[219]
port 635 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 sports_o[21]
port 636 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 sports_o[220]
port 637 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 sports_o[221]
port 638 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 sports_o[222]
port 639 nsew signal output
rlabel metal3 s 0 74536 800 74656 6 sports_o[223]
port 640 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 sports_o[224]
port 641 nsew signal output
rlabel metal3 s 0 75080 800 75200 6 sports_o[225]
port 642 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 sports_o[226]
port 643 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 sports_o[227]
port 644 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 sports_o[22]
port 645 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 sports_o[23]
port 646 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 sports_o[24]
port 647 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 sports_o[25]
port 648 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 sports_o[26]
port 649 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 sports_o[27]
port 650 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 sports_o[28]
port 651 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 sports_o[29]
port 652 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 sports_o[2]
port 653 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 sports_o[30]
port 654 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 sports_o[31]
port 655 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 sports_o[32]
port 656 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 sports_o[33]
port 657 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 sports_o[34]
port 658 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 sports_o[35]
port 659 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 sports_o[36]
port 660 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 sports_o[37]
port 661 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 sports_o[38]
port 662 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 sports_o[39]
port 663 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 sports_o[3]
port 664 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 sports_o[40]
port 665 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 sports_o[41]
port 666 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 sports_o[42]
port 667 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 sports_o[43]
port 668 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 sports_o[44]
port 669 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 sports_o[45]
port 670 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 sports_o[46]
port 671 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 sports_o[47]
port 672 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 sports_o[48]
port 673 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 sports_o[49]
port 674 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 sports_o[4]
port 675 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 sports_o[50]
port 676 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 sports_o[51]
port 677 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 sports_o[52]
port 678 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 sports_o[53]
port 679 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 sports_o[54]
port 680 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 sports_o[55]
port 681 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 sports_o[56]
port 682 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 sports_o[57]
port 683 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 sports_o[58]
port 684 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 sports_o[59]
port 685 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 sports_o[5]
port 686 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 sports_o[60]
port 687 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 sports_o[61]
port 688 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 sports_o[62]
port 689 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 sports_o[63]
port 690 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 sports_o[64]
port 691 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 sports_o[65]
port 692 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 sports_o[66]
port 693 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 sports_o[67]
port 694 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 sports_o[68]
port 695 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 sports_o[69]
port 696 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 sports_o[6]
port 697 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 sports_o[70]
port 698 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 sports_o[71]
port 699 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 sports_o[72]
port 700 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 sports_o[73]
port 701 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 sports_o[74]
port 702 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 sports_o[75]
port 703 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 sports_o[76]
port 704 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 sports_o[77]
port 705 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 sports_o[78]
port 706 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 sports_o[79]
port 707 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 sports_o[7]
port 708 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 sports_o[80]
port 709 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 sports_o[81]
port 710 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 sports_o[82]
port 711 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 sports_o[83]
port 712 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 sports_o[84]
port 713 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 sports_o[85]
port 714 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 sports_o[86]
port 715 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 sports_o[87]
port 716 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 sports_o[88]
port 717 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 sports_o[89]
port 718 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 sports_o[8]
port 719 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 sports_o[90]
port 720 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 sports_o[91]
port 721 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 sports_o[92]
port 722 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 sports_o[93]
port 723 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 sports_o[94]
port 724 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 sports_o[95]
port 725 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 sports_o[96]
port 726 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 sports_o[97]
port 727 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 sports_o[98]
port 728 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 sports_o[99]
port 729 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 sports_o[9]
port 730 nsew signal output
rlabel metal4 s 4208 2128 4528 87632 6 vccd1
port 731 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 87632 6 vccd1
port 731 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 87632 6 vccd1
port 731 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 87632 6 vssd1
port 732 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 87632 6 vssd1
port 732 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 87632 6 vssd1
port 732 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 24960800
string GDS_FILE /local/colinm22/sdmay26-24/openlane/busarb_2_2/runs/25_10_22_13_19/results/signoff/busarb_2_2.magic.gds
string GDS_START 876966
<< end >>

