VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac
  CLASS BLOCK ;
  FOREIGN mac ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 38.120 250.000 38.720 ;
    END
  END a_i[0]
  PIN a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 65.320 250.000 65.920 ;
    END
  END a_i[10]
  PIN a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 68.040 250.000 68.640 ;
    END
  END a_i[11]
  PIN a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 70.760 250.000 71.360 ;
    END
  END a_i[12]
  PIN a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 73.480 250.000 74.080 ;
    END
  END a_i[13]
  PIN a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 76.200 250.000 76.800 ;
    END
  END a_i[14]
  PIN a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 78.920 250.000 79.520 ;
    END
  END a_i[15]
  PIN a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 81.640 250.000 82.240 ;
    END
  END a_i[16]
  PIN a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 84.360 250.000 84.960 ;
    END
  END a_i[17]
  PIN a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 87.080 250.000 87.680 ;
    END
  END a_i[18]
  PIN a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 89.800 250.000 90.400 ;
    END
  END a_i[19]
  PIN a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 40.840 250.000 41.440 ;
    END
  END a_i[1]
  PIN a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 92.520 250.000 93.120 ;
    END
  END a_i[20]
  PIN a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 95.240 250.000 95.840 ;
    END
  END a_i[21]
  PIN a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 97.960 250.000 98.560 ;
    END
  END a_i[22]
  PIN a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 100.680 250.000 101.280 ;
    END
  END a_i[23]
  PIN a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 103.400 250.000 104.000 ;
    END
  END a_i[24]
  PIN a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 106.120 250.000 106.720 ;
    END
  END a_i[25]
  PIN a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 108.840 250.000 109.440 ;
    END
  END a_i[26]
  PIN a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 111.560 250.000 112.160 ;
    END
  END a_i[27]
  PIN a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 114.280 250.000 114.880 ;
    END
  END a_i[28]
  PIN a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 117.000 250.000 117.600 ;
    END
  END a_i[29]
  PIN a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 43.560 250.000 44.160 ;
    END
  END a_i[2]
  PIN a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 119.720 250.000 120.320 ;
    END
  END a_i[30]
  PIN a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 122.440 250.000 123.040 ;
    END
  END a_i[31]
  PIN a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 46.280 250.000 46.880 ;
    END
  END a_i[3]
  PIN a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 49.000 250.000 49.600 ;
    END
  END a_i[4]
  PIN a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 51.720 250.000 52.320 ;
    END
  END a_i[5]
  PIN a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 54.440 250.000 55.040 ;
    END
  END a_i[6]
  PIN a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 57.160 250.000 57.760 ;
    END
  END a_i[7]
  PIN a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 59.880 250.000 60.480 ;
    END
  END a_i[8]
  PIN a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 62.600 250.000 63.200 ;
    END
  END a_i[9]
  PIN b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 125.160 250.000 125.760 ;
    END
  END b_i[0]
  PIN b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 152.360 250.000 152.960 ;
    END
  END b_i[10]
  PIN b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 155.080 250.000 155.680 ;
    END
  END b_i[11]
  PIN b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 157.800 250.000 158.400 ;
    END
  END b_i[12]
  PIN b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 160.520 250.000 161.120 ;
    END
  END b_i[13]
  PIN b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 163.240 250.000 163.840 ;
    END
  END b_i[14]
  PIN b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 165.960 250.000 166.560 ;
    END
  END b_i[15]
  PIN b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 168.680 250.000 169.280 ;
    END
  END b_i[16]
  PIN b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 171.400 250.000 172.000 ;
    END
  END b_i[17]
  PIN b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 174.120 250.000 174.720 ;
    END
  END b_i[18]
  PIN b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 176.840 250.000 177.440 ;
    END
  END b_i[19]
  PIN b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 127.880 250.000 128.480 ;
    END
  END b_i[1]
  PIN b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 179.560 250.000 180.160 ;
    END
  END b_i[20]
  PIN b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 182.280 250.000 182.880 ;
    END
  END b_i[21]
  PIN b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 185.000 250.000 185.600 ;
    END
  END b_i[22]
  PIN b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 187.720 250.000 188.320 ;
    END
  END b_i[23]
  PIN b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 190.440 250.000 191.040 ;
    END
  END b_i[24]
  PIN b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 193.160 250.000 193.760 ;
    END
  END b_i[25]
  PIN b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 195.880 250.000 196.480 ;
    END
  END b_i[26]
  PIN b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 198.600 250.000 199.200 ;
    END
  END b_i[27]
  PIN b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 201.320 250.000 201.920 ;
    END
  END b_i[28]
  PIN b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 204.040 250.000 204.640 ;
    END
  END b_i[29]
  PIN b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 130.600 250.000 131.200 ;
    END
  END b_i[2]
  PIN b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 206.760 250.000 207.360 ;
    END
  END b_i[30]
  PIN b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 209.480 250.000 210.080 ;
    END
  END b_i[31]
  PIN b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 133.320 250.000 133.920 ;
    END
  END b_i[3]
  PIN b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 136.040 250.000 136.640 ;
    END
  END b_i[4]
  PIN b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 138.760 250.000 139.360 ;
    END
  END b_i[5]
  PIN b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 141.480 250.000 142.080 ;
    END
  END b_i[6]
  PIN b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 144.200 250.000 144.800 ;
    END
  END b_i[7]
  PIN b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 146.920 250.000 147.520 ;
    END
  END b_i[8]
  PIN b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 149.640 250.000 150.240 ;
    END
  END b_i[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END clk
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vssd1
  PIN y_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END y_o[0]
  PIN y_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END y_o[10]
  PIN y_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END y_o[11]
  PIN y_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END y_o[12]
  PIN y_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END y_o[13]
  PIN y_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END y_o[14]
  PIN y_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END y_o[15]
  PIN y_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END y_o[16]
  PIN y_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END y_o[17]
  PIN y_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END y_o[18]
  PIN y_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END y_o[19]
  PIN y_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END y_o[1]
  PIN y_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END y_o[20]
  PIN y_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END y_o[21]
  PIN y_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END y_o[22]
  PIN y_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END y_o[23]
  PIN y_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END y_o[24]
  PIN y_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END y_o[25]
  PIN y_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END y_o[26]
  PIN y_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END y_o[27]
  PIN y_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END y_o[28]
  PIN y_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END y_o[29]
  PIN y_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END y_o[2]
  PIN y_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END y_o[30]
  PIN y_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END y_o[31]
  PIN y_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END y_o[3]
  PIN y_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END y_o[4]
  PIN y_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END y_o[5]
  PIN y_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END y_o[6]
  PIN y_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END y_o[7]
  PIN y_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END y_o[8]
  PIN y_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END y_o[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 4.670 8.540 245.110 236.880 ;
      LAYER met2 ;
        RECT 4.690 4.280 245.090 236.825 ;
        RECT 4.690 4.000 61.910 4.280 ;
        RECT 62.750 4.000 186.570 4.280 ;
        RECT 187.410 4.000 245.090 4.280 ;
      LAYER met3 ;
        RECT 3.990 230.880 246.000 236.805 ;
        RECT 4.400 229.480 246.000 230.880 ;
        RECT 3.990 224.080 246.000 229.480 ;
        RECT 4.400 222.680 246.000 224.080 ;
        RECT 3.990 217.280 246.000 222.680 ;
        RECT 4.400 215.880 246.000 217.280 ;
        RECT 3.990 210.480 246.000 215.880 ;
        RECT 4.400 209.080 245.600 210.480 ;
        RECT 3.990 207.760 246.000 209.080 ;
        RECT 3.990 206.360 245.600 207.760 ;
        RECT 3.990 205.040 246.000 206.360 ;
        RECT 3.990 203.680 245.600 205.040 ;
        RECT 4.400 203.640 245.600 203.680 ;
        RECT 4.400 202.320 246.000 203.640 ;
        RECT 4.400 202.280 245.600 202.320 ;
        RECT 3.990 200.920 245.600 202.280 ;
        RECT 3.990 199.600 246.000 200.920 ;
        RECT 3.990 198.200 245.600 199.600 ;
        RECT 3.990 196.880 246.000 198.200 ;
        RECT 4.400 195.480 245.600 196.880 ;
        RECT 3.990 194.160 246.000 195.480 ;
        RECT 3.990 192.760 245.600 194.160 ;
        RECT 3.990 191.440 246.000 192.760 ;
        RECT 3.990 190.080 245.600 191.440 ;
        RECT 4.400 190.040 245.600 190.080 ;
        RECT 4.400 188.720 246.000 190.040 ;
        RECT 4.400 188.680 245.600 188.720 ;
        RECT 3.990 187.320 245.600 188.680 ;
        RECT 3.990 186.000 246.000 187.320 ;
        RECT 3.990 184.600 245.600 186.000 ;
        RECT 3.990 183.280 246.000 184.600 ;
        RECT 4.400 181.880 245.600 183.280 ;
        RECT 3.990 180.560 246.000 181.880 ;
        RECT 3.990 179.160 245.600 180.560 ;
        RECT 3.990 177.840 246.000 179.160 ;
        RECT 3.990 176.480 245.600 177.840 ;
        RECT 4.400 176.440 245.600 176.480 ;
        RECT 4.400 175.120 246.000 176.440 ;
        RECT 4.400 175.080 245.600 175.120 ;
        RECT 3.990 173.720 245.600 175.080 ;
        RECT 3.990 172.400 246.000 173.720 ;
        RECT 3.990 171.000 245.600 172.400 ;
        RECT 3.990 169.680 246.000 171.000 ;
        RECT 4.400 168.280 245.600 169.680 ;
        RECT 3.990 166.960 246.000 168.280 ;
        RECT 3.990 165.560 245.600 166.960 ;
        RECT 3.990 164.240 246.000 165.560 ;
        RECT 3.990 162.880 245.600 164.240 ;
        RECT 4.400 162.840 245.600 162.880 ;
        RECT 4.400 161.520 246.000 162.840 ;
        RECT 4.400 161.480 245.600 161.520 ;
        RECT 3.990 160.120 245.600 161.480 ;
        RECT 3.990 158.800 246.000 160.120 ;
        RECT 3.990 157.400 245.600 158.800 ;
        RECT 3.990 156.080 246.000 157.400 ;
        RECT 4.400 154.680 245.600 156.080 ;
        RECT 3.990 153.360 246.000 154.680 ;
        RECT 3.990 151.960 245.600 153.360 ;
        RECT 3.990 150.640 246.000 151.960 ;
        RECT 3.990 149.280 245.600 150.640 ;
        RECT 4.400 149.240 245.600 149.280 ;
        RECT 4.400 147.920 246.000 149.240 ;
        RECT 4.400 147.880 245.600 147.920 ;
        RECT 3.990 146.520 245.600 147.880 ;
        RECT 3.990 145.200 246.000 146.520 ;
        RECT 3.990 143.800 245.600 145.200 ;
        RECT 3.990 142.480 246.000 143.800 ;
        RECT 4.400 141.080 245.600 142.480 ;
        RECT 3.990 139.760 246.000 141.080 ;
        RECT 3.990 138.360 245.600 139.760 ;
        RECT 3.990 137.040 246.000 138.360 ;
        RECT 3.990 135.680 245.600 137.040 ;
        RECT 4.400 135.640 245.600 135.680 ;
        RECT 4.400 134.320 246.000 135.640 ;
        RECT 4.400 134.280 245.600 134.320 ;
        RECT 3.990 132.920 245.600 134.280 ;
        RECT 3.990 131.600 246.000 132.920 ;
        RECT 3.990 130.200 245.600 131.600 ;
        RECT 3.990 128.880 246.000 130.200 ;
        RECT 4.400 127.480 245.600 128.880 ;
        RECT 3.990 126.160 246.000 127.480 ;
        RECT 3.990 124.760 245.600 126.160 ;
        RECT 3.990 123.440 246.000 124.760 ;
        RECT 3.990 122.080 245.600 123.440 ;
        RECT 4.400 122.040 245.600 122.080 ;
        RECT 4.400 120.720 246.000 122.040 ;
        RECT 4.400 120.680 245.600 120.720 ;
        RECT 3.990 119.320 245.600 120.680 ;
        RECT 3.990 118.000 246.000 119.320 ;
        RECT 3.990 116.600 245.600 118.000 ;
        RECT 3.990 115.280 246.000 116.600 ;
        RECT 4.400 113.880 245.600 115.280 ;
        RECT 3.990 112.560 246.000 113.880 ;
        RECT 3.990 111.160 245.600 112.560 ;
        RECT 3.990 109.840 246.000 111.160 ;
        RECT 3.990 108.480 245.600 109.840 ;
        RECT 4.400 108.440 245.600 108.480 ;
        RECT 4.400 107.120 246.000 108.440 ;
        RECT 4.400 107.080 245.600 107.120 ;
        RECT 3.990 105.720 245.600 107.080 ;
        RECT 3.990 104.400 246.000 105.720 ;
        RECT 3.990 103.000 245.600 104.400 ;
        RECT 3.990 101.680 246.000 103.000 ;
        RECT 4.400 100.280 245.600 101.680 ;
        RECT 3.990 98.960 246.000 100.280 ;
        RECT 3.990 97.560 245.600 98.960 ;
        RECT 3.990 96.240 246.000 97.560 ;
        RECT 3.990 94.880 245.600 96.240 ;
        RECT 4.400 94.840 245.600 94.880 ;
        RECT 4.400 93.520 246.000 94.840 ;
        RECT 4.400 93.480 245.600 93.520 ;
        RECT 3.990 92.120 245.600 93.480 ;
        RECT 3.990 90.800 246.000 92.120 ;
        RECT 3.990 89.400 245.600 90.800 ;
        RECT 3.990 88.080 246.000 89.400 ;
        RECT 4.400 86.680 245.600 88.080 ;
        RECT 3.990 85.360 246.000 86.680 ;
        RECT 3.990 83.960 245.600 85.360 ;
        RECT 3.990 82.640 246.000 83.960 ;
        RECT 3.990 81.280 245.600 82.640 ;
        RECT 4.400 81.240 245.600 81.280 ;
        RECT 4.400 79.920 246.000 81.240 ;
        RECT 4.400 79.880 245.600 79.920 ;
        RECT 3.990 78.520 245.600 79.880 ;
        RECT 3.990 77.200 246.000 78.520 ;
        RECT 3.990 75.800 245.600 77.200 ;
        RECT 3.990 74.480 246.000 75.800 ;
        RECT 4.400 73.080 245.600 74.480 ;
        RECT 3.990 71.760 246.000 73.080 ;
        RECT 3.990 70.360 245.600 71.760 ;
        RECT 3.990 69.040 246.000 70.360 ;
        RECT 3.990 67.680 245.600 69.040 ;
        RECT 4.400 67.640 245.600 67.680 ;
        RECT 4.400 66.320 246.000 67.640 ;
        RECT 4.400 66.280 245.600 66.320 ;
        RECT 3.990 64.920 245.600 66.280 ;
        RECT 3.990 63.600 246.000 64.920 ;
        RECT 3.990 62.200 245.600 63.600 ;
        RECT 3.990 60.880 246.000 62.200 ;
        RECT 4.400 59.480 245.600 60.880 ;
        RECT 3.990 58.160 246.000 59.480 ;
        RECT 3.990 56.760 245.600 58.160 ;
        RECT 3.990 55.440 246.000 56.760 ;
        RECT 3.990 54.080 245.600 55.440 ;
        RECT 4.400 54.040 245.600 54.080 ;
        RECT 4.400 52.720 246.000 54.040 ;
        RECT 4.400 52.680 245.600 52.720 ;
        RECT 3.990 51.320 245.600 52.680 ;
        RECT 3.990 50.000 246.000 51.320 ;
        RECT 3.990 48.600 245.600 50.000 ;
        RECT 3.990 47.280 246.000 48.600 ;
        RECT 4.400 45.880 245.600 47.280 ;
        RECT 3.990 44.560 246.000 45.880 ;
        RECT 3.990 43.160 245.600 44.560 ;
        RECT 3.990 41.840 246.000 43.160 ;
        RECT 3.990 40.480 245.600 41.840 ;
        RECT 4.400 40.440 245.600 40.480 ;
        RECT 4.400 39.120 246.000 40.440 ;
        RECT 4.400 39.080 245.600 39.120 ;
        RECT 3.990 37.720 245.600 39.080 ;
        RECT 3.990 33.680 246.000 37.720 ;
        RECT 4.400 32.280 246.000 33.680 ;
        RECT 3.990 26.880 246.000 32.280 ;
        RECT 4.400 25.480 246.000 26.880 ;
        RECT 3.990 20.080 246.000 25.480 ;
        RECT 4.400 18.680 246.000 20.080 ;
        RECT 3.990 10.715 246.000 18.680 ;
      LAYER met4 ;
        RECT 19.615 19.215 20.640 228.305 ;
        RECT 23.040 19.215 97.440 228.305 ;
        RECT 99.840 19.215 174.240 228.305 ;
        RECT 176.640 19.215 240.745 228.305 ;
  END
END mac
END LIBRARY

