* NGSPICE file created from busarb_2_2.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt busarb_2_2 clk_i mports_i[0] mports_i[100] mports_i[101] mports_i[102] mports_i[103]
+ mports_i[104] mports_i[105] mports_i[106] mports_i[107] mports_i[108] mports_i[109]
+ mports_i[10] mports_i[110] mports_i[111] mports_i[112] mports_i[113] mports_i[114]
+ mports_i[115] mports_i[116] mports_i[117] mports_i[118] mports_i[119] mports_i[11]
+ mports_i[120] mports_i[121] mports_i[122] mports_i[123] mports_i[124] mports_i[125]
+ mports_i[126] mports_i[127] mports_i[128] mports_i[129] mports_i[12] mports_i[130]
+ mports_i[131] mports_i[132] mports_i[133] mports_i[134] mports_i[135] mports_i[136]
+ mports_i[137] mports_i[138] mports_i[139] mports_i[13] mports_i[140] mports_i[141]
+ mports_i[142] mports_i[143] mports_i[144] mports_i[145] mports_i[146] mports_i[147]
+ mports_i[148] mports_i[149] mports_i[14] mports_i[150] mports_i[151] mports_i[152]
+ mports_i[153] mports_i[154] mports_i[155] mports_i[156] mports_i[157] mports_i[158]
+ mports_i[159] mports_i[15] mports_i[160] mports_i[161] mports_i[162] mports_i[163]
+ mports_i[164] mports_i[165] mports_i[166] mports_i[167] mports_i[168] mports_i[169]
+ mports_i[16] mports_i[170] mports_i[171] mports_i[172] mports_i[173] mports_i[174]
+ mports_i[175] mports_i[176] mports_i[177] mports_i[178] mports_i[179] mports_i[17]
+ mports_i[180] mports_i[181] mports_i[182] mports_i[183] mports_i[184] mports_i[185]
+ mports_i[186] mports_i[187] mports_i[188] mports_i[189] mports_i[18] mports_i[190]
+ mports_i[191] mports_i[192] mports_i[193] mports_i[194] mports_i[195] mports_i[196]
+ mports_i[197] mports_i[198] mports_i[199] mports_i[19] mports_i[1] mports_i[200]
+ mports_i[201] mports_i[202] mports_i[203] mports_i[204] mports_i[205] mports_i[206]
+ mports_i[207] mports_i[208] mports_i[209] mports_i[20] mports_i[210] mports_i[211]
+ mports_i[212] mports_i[213] mports_i[214] mports_i[215] mports_i[216] mports_i[217]
+ mports_i[218] mports_i[219] mports_i[21] mports_i[220] mports_i[221] mports_i[222]
+ mports_i[223] mports_i[224] mports_i[225] mports_i[226] mports_i[227] mports_i[22]
+ mports_i[23] mports_i[24] mports_i[25] mports_i[26] mports_i[27] mports_i[28] mports_i[29]
+ mports_i[2] mports_i[30] mports_i[31] mports_i[32] mports_i[33] mports_i[34] mports_i[35]
+ mports_i[36] mports_i[37] mports_i[38] mports_i[39] mports_i[3] mports_i[40] mports_i[41]
+ mports_i[42] mports_i[43] mports_i[44] mports_i[45] mports_i[46] mports_i[47] mports_i[48]
+ mports_i[49] mports_i[4] mports_i[50] mports_i[51] mports_i[52] mports_i[53] mports_i[54]
+ mports_i[55] mports_i[56] mports_i[57] mports_i[58] mports_i[59] mports_i[5] mports_i[60]
+ mports_i[61] mports_i[62] mports_i[63] mports_i[64] mports_i[65] mports_i[66] mports_i[67]
+ mports_i[68] mports_i[69] mports_i[6] mports_i[70] mports_i[71] mports_i[72] mports_i[73]
+ mports_i[74] mports_i[75] mports_i[76] mports_i[77] mports_i[78] mports_i[79] mports_i[7]
+ mports_i[80] mports_i[81] mports_i[82] mports_i[83] mports_i[84] mports_i[85] mports_i[86]
+ mports_i[87] mports_i[88] mports_i[89] mports_i[8] mports_i[90] mports_i[91] mports_i[92]
+ mports_i[93] mports_i[94] mports_i[95] mports_i[96] mports_i[97] mports_i[98] mports_i[99]
+ mports_i[9] mports_o[0] mports_o[100] mports_o[101] mports_o[102] mports_o[103]
+ mports_o[104] mports_o[105] mports_o[106] mports_o[107] mports_o[108] mports_o[109]
+ mports_o[10] mports_o[110] mports_o[111] mports_o[112] mports_o[113] mports_o[114]
+ mports_o[115] mports_o[116] mports_o[117] mports_o[118] mports_o[119] mports_o[11]
+ mports_o[120] mports_o[121] mports_o[122] mports_o[123] mports_o[124] mports_o[125]
+ mports_o[126] mports_o[127] mports_o[128] mports_o[129] mports_o[12] mports_o[130]
+ mports_o[131] mports_o[132] mports_o[133] mports_o[134] mports_o[135] mports_o[13]
+ mports_o[14] mports_o[15] mports_o[16] mports_o[17] mports_o[18] mports_o[19] mports_o[1]
+ mports_o[20] mports_o[21] mports_o[22] mports_o[23] mports_o[24] mports_o[25] mports_o[26]
+ mports_o[27] mports_o[28] mports_o[29] mports_o[2] mports_o[30] mports_o[31] mports_o[32]
+ mports_o[33] mports_o[34] mports_o[35] mports_o[36] mports_o[37] mports_o[38] mports_o[39]
+ mports_o[3] mports_o[40] mports_o[41] mports_o[42] mports_o[43] mports_o[44] mports_o[45]
+ mports_o[46] mports_o[47] mports_o[48] mports_o[49] mports_o[4] mports_o[50] mports_o[51]
+ mports_o[52] mports_o[53] mports_o[54] mports_o[55] mports_o[56] mports_o[57] mports_o[58]
+ mports_o[59] mports_o[5] mports_o[60] mports_o[61] mports_o[62] mports_o[63] mports_o[64]
+ mports_o[65] mports_o[66] mports_o[67] mports_o[68] mports_o[69] mports_o[6] mports_o[70]
+ mports_o[71] mports_o[72] mports_o[73] mports_o[74] mports_o[75] mports_o[76] mports_o[77]
+ mports_o[78] mports_o[79] mports_o[7] mports_o[80] mports_o[81] mports_o[82] mports_o[83]
+ mports_o[84] mports_o[85] mports_o[86] mports_o[87] mports_o[88] mports_o[89] mports_o[8]
+ mports_o[90] mports_o[91] mports_o[92] mports_o[93] mports_o[94] mports_o[95] mports_o[96]
+ mports_o[97] mports_o[98] mports_o[99] mports_o[9] nrst_i sports_i[0] sports_i[100]
+ sports_i[101] sports_i[102] sports_i[103] sports_i[104] sports_i[105] sports_i[106]
+ sports_i[107] sports_i[108] sports_i[109] sports_i[10] sports_i[110] sports_i[111]
+ sports_i[112] sports_i[113] sports_i[114] sports_i[115] sports_i[116] sports_i[117]
+ sports_i[118] sports_i[119] sports_i[11] sports_i[120] sports_i[121] sports_i[122]
+ sports_i[123] sports_i[124] sports_i[125] sports_i[126] sports_i[127] sports_i[128]
+ sports_i[129] sports_i[12] sports_i[130] sports_i[131] sports_i[132] sports_i[133]
+ sports_i[134] sports_i[135] sports_i[13] sports_i[14] sports_i[15] sports_i[16]
+ sports_i[17] sports_i[18] sports_i[19] sports_i[1] sports_i[20] sports_i[21] sports_i[22]
+ sports_i[23] sports_i[24] sports_i[25] sports_i[26] sports_i[27] sports_i[28] sports_i[29]
+ sports_i[2] sports_i[30] sports_i[31] sports_i[32] sports_i[33] sports_i[34] sports_i[35]
+ sports_i[36] sports_i[37] sports_i[38] sports_i[39] sports_i[3] sports_i[40] sports_i[41]
+ sports_i[42] sports_i[43] sports_i[44] sports_i[45] sports_i[46] sports_i[47] sports_i[48]
+ sports_i[49] sports_i[4] sports_i[50] sports_i[51] sports_i[52] sports_i[53] sports_i[54]
+ sports_i[55] sports_i[56] sports_i[57] sports_i[58] sports_i[59] sports_i[5] sports_i[60]
+ sports_i[61] sports_i[62] sports_i[63] sports_i[64] sports_i[65] sports_i[66] sports_i[67]
+ sports_i[68] sports_i[69] sports_i[6] sports_i[70] sports_i[71] sports_i[72] sports_i[73]
+ sports_i[74] sports_i[75] sports_i[76] sports_i[77] sports_i[78] sports_i[79] sports_i[7]
+ sports_i[80] sports_i[81] sports_i[82] sports_i[83] sports_i[84] sports_i[85] sports_i[86]
+ sports_i[87] sports_i[88] sports_i[89] sports_i[8] sports_i[90] sports_i[91] sports_i[92]
+ sports_i[93] sports_i[94] sports_i[95] sports_i[96] sports_i[97] sports_i[98] sports_i[99]
+ sports_i[9] sports_o[0] sports_o[100] sports_o[101] sports_o[102] sports_o[103]
+ sports_o[104] sports_o[105] sports_o[106] sports_o[107] sports_o[108] sports_o[109]
+ sports_o[10] sports_o[110] sports_o[111] sports_o[112] sports_o[113] sports_o[114]
+ sports_o[115] sports_o[116] sports_o[117] sports_o[118] sports_o[119] sports_o[11]
+ sports_o[120] sports_o[121] sports_o[122] sports_o[123] sports_o[124] sports_o[125]
+ sports_o[126] sports_o[127] sports_o[128] sports_o[129] sports_o[12] sports_o[130]
+ sports_o[131] sports_o[132] sports_o[133] sports_o[134] sports_o[135] sports_o[136]
+ sports_o[137] sports_o[138] sports_o[139] sports_o[13] sports_o[140] sports_o[141]
+ sports_o[142] sports_o[143] sports_o[144] sports_o[145] sports_o[146] sports_o[147]
+ sports_o[148] sports_o[149] sports_o[14] sports_o[150] sports_o[151] sports_o[152]
+ sports_o[153] sports_o[154] sports_o[155] sports_o[156] sports_o[157] sports_o[158]
+ sports_o[159] sports_o[15] sports_o[160] sports_o[161] sports_o[162] sports_o[163]
+ sports_o[164] sports_o[165] sports_o[166] sports_o[167] sports_o[168] sports_o[169]
+ sports_o[16] sports_o[170] sports_o[171] sports_o[172] sports_o[173] sports_o[174]
+ sports_o[175] sports_o[176] sports_o[177] sports_o[178] sports_o[179] sports_o[17]
+ sports_o[180] sports_o[181] sports_o[182] sports_o[183] sports_o[184] sports_o[185]
+ sports_o[186] sports_o[187] sports_o[188] sports_o[189] sports_o[18] sports_o[190]
+ sports_o[191] sports_o[192] sports_o[193] sports_o[194] sports_o[195] sports_o[196]
+ sports_o[197] sports_o[198] sports_o[199] sports_o[19] sports_o[1] sports_o[200]
+ sports_o[201] sports_o[202] sports_o[203] sports_o[204] sports_o[205] sports_o[206]
+ sports_o[207] sports_o[208] sports_o[209] sports_o[20] sports_o[210] sports_o[211]
+ sports_o[212] sports_o[213] sports_o[214] sports_o[215] sports_o[216] sports_o[217]
+ sports_o[218] sports_o[219] sports_o[21] sports_o[220] sports_o[221] sports_o[222]
+ sports_o[223] sports_o[224] sports_o[225] sports_o[226] sports_o[227] sports_o[22]
+ sports_o[23] sports_o[24] sports_o[25] sports_o[26] sports_o[27] sports_o[28] sports_o[29]
+ sports_o[2] sports_o[30] sports_o[31] sports_o[32] sports_o[33] sports_o[34] sports_o[35]
+ sports_o[36] sports_o[37] sports_o[38] sports_o[39] sports_o[3] sports_o[40] sports_o[41]
+ sports_o[42] sports_o[43] sports_o[44] sports_o[45] sports_o[46] sports_o[47] sports_o[48]
+ sports_o[49] sports_o[4] sports_o[50] sports_o[51] sports_o[52] sports_o[53] sports_o[54]
+ sports_o[55] sports_o[56] sports_o[57] sports_o[58] sports_o[59] sports_o[5] sports_o[60]
+ sports_o[61] sports_o[62] sports_o[63] sports_o[64] sports_o[65] sports_o[66] sports_o[67]
+ sports_o[68] sports_o[69] sports_o[6] sports_o[70] sports_o[71] sports_o[72] sports_o[73]
+ sports_o[74] sports_o[75] sports_o[76] sports_o[77] sports_o[78] sports_o[79] sports_o[7]
+ sports_o[80] sports_o[81] sports_o[82] sports_o[83] sports_o[84] sports_o[85] sports_o[86]
+ sports_o[87] sports_o[88] sports_o[89] sports_o[8] sports_o[90] sports_o[91] sports_o[92]
+ sports_o[93] sports_o[94] sports_o[95] sports_o[96] sports_o[97] sports_o[98] sports_o[99]
+ sports_o[9] vccd1 vssd1
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7406__A1 _5248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8603__B1 _7832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7406__B2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4935__A _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7311__A _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7957__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7963_ _7963_/A vssd1 vssd1 vccd1 vccd1 _7963_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5968__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6914_ _7707_/B _6914_/B vssd1 vssd1 vccd1 vccd1 _6914_/X sky130_fd_sc_hd__or2_1
X_7894_ _8333_/A _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _7894_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__7709__A2 _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6845_ _6845_/A vssd1 vssd1 vccd1 vccd1 _7604_/B sky130_fd_sc_hd__inv_2
XFILLER_0_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8382__A2 _8381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8142__A _8142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6393__A1 _6400_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6776_ _6774_/X _6899_/B _7000_/S _6775_/X vssd1 vssd1 vccd1 vccd1 _6776_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6393__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8515_ _8515_/A _8516_/B vssd1 vssd1 vccd1 vccd1 _8515_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5727_ _5727_/A vssd1 vssd1 vccd1 vccd1 _5727_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_134_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8134__A2 _8133_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6145__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8446_ _8445_/Y _8416_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8446_/X sky130_fd_sc_hd__mux2_1
X_5658_ _5658_/A vssd1 vssd1 vccd1 vccd1 _7514_/A sky130_fd_sc_hd__inv_2
XANTENNA__6145__B2 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7893__A1 _7881_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4609_ _4608_/X _4511_/B _4511_/A _7510_/A vssd1 vssd1 vccd1 vccd1 _4610_/B sky130_fd_sc_hd__a31o_1
X_8377_ _8375_/Y _8376_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8378_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7893__B2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6597__A _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5589_ _5586_/X _5645_/A _6224_/S vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7328_ _4992_/X _7723_/B _7327_/X vssd1 vssd1 vccd1 vccd1 _7328_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7259_ _7258_/X _7725_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7260_/A sky130_fd_sc_hd__mux2_2
XANTENNA__5120__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8070__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6384__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8125__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6136__A1 _6136_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6136__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6687__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5895__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7115__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7636__A1 _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7939__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4960_ _4960_/A vssd1 vssd1 vccd1 vccd1 _6456_/A sky130_fd_sc_hd__inv_2
XFILLER_0_148_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4891_ _4891_/A vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__buf_8
XFILLER_0_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7021__C1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6630_ _6630_/A _6908_/B vssd1 vssd1 vccd1 vccd1 _6630_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5178__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6561_ _5219_/B _6913_/B _6557_/Y _6559_/Y _6560_/Y vssd1 vssd1 vccd1 vccd1 _6562_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8116__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8300_ _8455_/B _8300_/B vssd1 vssd1 vccd1 vccd1 _8755_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5274_/X _5543_/A1 _4896_/A input39/X vssd1 vssd1 vccd1 vccd1 _5512_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__6127__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6492_ _6958_/B _5109_/B _6450_/A vssd1 vssd1 vccd1 vccd1 _6492_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8231_ _6965_/A _8234_/A2 _8163_/A _8234_/B2 vssd1 vssd1 vccd1 vccd1 _8231_/X sky130_fd_sc_hd__a22o_1
X_5443_ _5440_/Y _4886_/A _5441_/Y _4891_/A _5442_/Y vssd1 vssd1 vccd1 vccd1 _6653_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput401 _8826_/X vssd1 vssd1 vccd1 vccd1 mports_o[131] sky130_fd_sc_hd__buf_12
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput412 _8057_/X vssd1 vssd1 vccd1 vccd1 mports_o[19] sky130_fd_sc_hd__buf_12
Xoutput423 _8213_/X vssd1 vssd1 vccd1 vccd1 mports_o[29] sky130_fd_sc_hd__buf_12
XANTENNA__7306__A _7306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput434 _8322_/X vssd1 vssd1 vccd1 vccd1 mports_o[39] sky130_fd_sc_hd__buf_12
X_8162_ _8162_/A vssd1 vssd1 vccd1 vccd1 _8174_/B sky130_fd_sc_hd__inv_2
XANTENNA__5350__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5374_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5374_/Y sky130_fd_sc_hd__inv_2
Xoutput445 _8411_/X vssd1 vssd1 vccd1 vccd1 mports_o[49] sky130_fd_sc_hd__buf_12
Xoutput456 _8528_/X vssd1 vssd1 vccd1 vccd1 mports_o[59] sky130_fd_sc_hd__buf_12
Xoutput467 _8596_/X vssd1 vssd1 vccd1 vccd1 mports_o[69] sky130_fd_sc_hd__buf_12
X_7113_ _7112_/X _5464_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7114_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7627__A1 _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput478 _8629_/X vssd1 vssd1 vccd1 vccd1 mports_o[79] sky130_fd_sc_hd__buf_12
X_4325_ _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__nand2_1
Xoutput489 _8664_/X vssd1 vssd1 vccd1 vccd1 mports_o[89] sky130_fd_sc_hd__buf_12
X_8093_ _8093_/A1 _7876_/X _8093_/B1 _7835_/A vssd1 vssd1 vccd1 vccd1 _8093_/Y sky130_fd_sc_hd__o22ai_1
X_7044_ _6488_/A _7088_/A _7043_/Y _7059_/A _7089_/A vssd1 vssd1 vccd1 vccd1 _7044_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6356__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6850__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8052__B2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4384__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6602__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7946_ _7777_/X _7945_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _7946_/X sky130_fd_sc_hd__o21ba_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7877_ _7877_/A1 _7876_/X _7877_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7877_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__8355__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6366__A1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6828_ _6828_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6828_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6366__B2 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7563__B1 _7559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6759_ _5737_/A _6912_/B _6755_/Y _6757_/Y _6758_/Y vssd1 vssd1 vccd1 vccd1 _6760_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8107__A2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7866__A1 _7877_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8429_ _8429_/A vssd1 vssd1 vccd1 vccd1 _8429_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7866__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4559__B hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7079__C1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7618__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8043__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5801__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7097__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__A1 _6357_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6357__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7554__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8510__A _8510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6109__A1 _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5868__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5332__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7609__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6965__A _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output728_A _6930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8282__A1 _7796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7085__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5090_ _5090_/A vssd1 vssd1 vccd1 vccd1 _8709_/B sky130_fd_sc_hd__buf_8
XFILLER_0_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6832__A2 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8034__A1 _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8391__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7800_ _4326_/B _6500_/A _7802_/A2 _7769_/X _7799_/X vssd1 vssd1 vccd1 vccd1 _7800_/X
+ sky130_fd_sc_hd__a221o_4
X_8780_ _8412_/A _8806_/B _8778_/X _8779_/X vssd1 vssd1 vccd1 vccd1 _8780_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5992_ _6079_/A _6046_/A vssd1 vssd1 vccd1 vccd1 _5992_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5399__A2 _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7731_ _6333_/Y _7349_/A _7266_/X _7753_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7731_/X
+ sky130_fd_sc_hd__a221o_1
X_4943_ _4943_/A vssd1 vssd1 vccd1 vccd1 _7372_/B sky130_fd_sc_hd__inv_6
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8404__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6348__A1 _6357_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7662_ _6112_/B _7696_/B _6915_/Y _7361_/X vssd1 vssd1 vccd1 vccd1 _7662_/X sky130_fd_sc_hd__a22o_1
X_4874_ _4874_/A vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__buf_8
XANTENNA__6348__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7545__B1 _7543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8742__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6613_ _6906_/A _6613_/B vssd1 vssd1 vccd1 vccd1 _6613_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7593_ _7532_/A _6809_/B _7348_/A vssd1 vssd1 vccd1 vccd1 _7593_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6544_ _6544_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6544_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5571__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6859__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6475_ _6475_/A vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__buf_6
XFILLER_0_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5859__B1 _5867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7036__A _7036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8214_ _7761_/A _8221_/A2 _5117_/A _4478_/B vssd1 vssd1 vccd1 vccd1 _8214_/X sky130_fd_sc_hd__a22o_1
X_5426_ _5426_/A vssd1 vssd1 vccd1 vccd1 _5426_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_140_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8145_ _8145_/A vssd1 vssd1 vccd1 vccd1 _8145_/Y sky130_fd_sc_hd__inv_2
X_5357_ input94/X _4935_/A input31/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5357_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8273__A1 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7076__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4308_ hold39/X _4719_/B vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__nor2_4
X_8076_ _8071_/Y _6079_/A _8072_/Y _6513_/A _8075_/Y vssd1 vssd1 vccd1 vccd1 _8483_/A
+ sky130_fd_sc_hd__a221oi_4
X_5288_ _5288_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _5288_/Y sky130_fd_sc_hd__nand2_1
X_7027_ _7027_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7027_/X sky130_fd_sc_hd__and2_1
XANTENNA__8025__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8978_ _8978_/CLK _8978_/D fanout732/X vssd1 vssd1 vccd1 vccd1 _8978_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__7784__B1 _7791_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4598__B1 _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7929_ _7922_/Y _7769_/X _7923_/Y _6500_/X _7928_/Y vssd1 vssd1 vccd1 vccd1 _7929_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8328__A2 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6339__A1 _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6115__A _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5562__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7839__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5314__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7067__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6275__B1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6814__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7775__B1 _7771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5250__A1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5250__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7527__B1 _7525_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8240__A _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4590_ _4590_/A _4590_/B vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5553__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6679__B _6679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6750__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6260_ _6253_/A _8516_/B input6/X _4913_/X _6259_/X vssd1 vssd1 vccd1 vccd1 _6261_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6502__A1 _6543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5211_ _5211_/A vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__inv_2
XANTENNA__6695__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6191_ _6170_/X _6402_/A _6179_/Y _6181_/Y _6190_/X vssd1 vssd1 vccd1 vccd1 _6191_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__7290__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5142_ _5139_/Y _8455_/B _5140_/Y _4891_/X _5141_/Y vssd1 vssd1 vccd1 vccd1 _6514_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6805__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5608__A3 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5073_ _5070_/Y _8455_/B _5071_/Y _4891_/X _5072_/Y vssd1 vssd1 vccd1 vccd1 _5075_/B
+ sky130_fd_sc_hd__o221a_2
X_8901_ _4800_/B _8706_/B _4662_/C _8574_/B vssd1 vssd1 vccd1 vccd1 _8901_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__8007__B2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8832_ _8230_/Y _8711_/A _8232_/X _8738_/A vssd1 vssd1 vccd1 vccd1 _8833_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5975_ _5972_/X _6837_/B _6711_/S vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__mux2_1
X_8763_ _8402_/X _8759_/Y _8762_/X _8725_/X vssd1 vssd1 vccd1 vccd1 _8763_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4662__B _7737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5241__A1 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5241__B2 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4926_ _4908_/X _4919_/X _6356_/S vssd1 vssd1 vccd1 vccd1 _4926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7714_ _6252_/X _7640_/B _7713_/X vssd1 vssd1 vccd1 vccd1 _7714_/X sky130_fd_sc_hd__o21a_1
XANTENNA__7518__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5792__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8694_ _8574_/B hold30/A _8263_/X _8693_/X _8590_/X vssd1 vssd1 vccd1 vccd1 _8694_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4857_ _8929_/B _4857_/B vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__nand2_1
X_7645_ _7646_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8191__B1 _8190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8730__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8150__A _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7576_ _5827_/A _7660_/B _7574_/X _7348_/A _7575_/Y vssd1 vssd1 vccd1 vccd1 _7576_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_145_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5544__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4788_ _4788_/A _4788_/B _4788_/C vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6527_ _6912_/B _5184_/X _7366_/B _6841_/A vssd1 vssd1 vccd1 vccd1 _6527_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_132_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6458_ _6724_/A vssd1 vssd1 vccd1 vccd1 _6473_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _6304_/A _7094_/A vssd1 vssd1 vccd1 vccd1 _5409_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6389_ _6402_/A _7750_/B vssd1 vssd1 vccd1 vccd1 _6389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8128_ _8123_/Y _6965_/A _8124_/Y _8163_/A _8127_/Y vssd1 vssd1 vccd1 vccd1 _8550_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7049__A2 _6499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8246__B2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5940__C _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8797__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8059_ _8059_/A vssd1 vssd1 vccd1 vccd1 _8059_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4807__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6009__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5480__A1 _5518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8549__A2 _8169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5480__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4991__B1 _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8182__B1 hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8721__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8237__A1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4747__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6248__B1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output426_A _8237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6799__A1 _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7748__B1 _7349_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4482__B _4566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5223__A1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5223__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5760_ _5760_/A _6593_/A vssd1 vssd1 vccd1 vccd1 _5760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4711_ _4711_/A hold35/X vssd1 vssd1 vccd1 vccd1 _4771_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5691_/A vssd1 vssd1 vccd1 vccd1 _7531_/A sky130_fd_sc_hd__inv_2
XANTENNA__7285__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7515__A3 _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7430_ _5317_/A _7681_/A _7673_/A _5353_/Y _7756_/A vssd1 vssd1 vccd1 vccd1 _7430_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4642_ hold30/A vssd1 vssd1 vccd1 vccd1 _4643_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6723__A1 _6719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7361_ _7476_/B vssd1 vssd1 vccd1 vccd1 _7361_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4573_ hold43/X vssd1 vssd1 vccd1 vccd1 _8336_/S sky130_fd_sc_hd__buf_4
XFILLER_0_71_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6202__B _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6312_ _6312_/A _6312_/B vssd1 vssd1 vccd1 vccd1 _6312_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7279__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7292_ _7753_/A _7059_/A _6397_/X _7088_/A _7089_/A vssd1 vssd1 vccd1 vccd1 _7292_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6243_ input68/X _8579_/C _6247_/A1 _8713_/C _6242_/X vssd1 vssd1 vccd1 vccd1 _6244_/A
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4938__A _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8228__A1 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6174_ _6174_/A1 _5192_/A input64/X _5193_/A vssd1 vssd1 vccd1 vccd1 _6174_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8228__B2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6239__B1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8779__A2 _8012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5125_ _5893_/B vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__clkbuf_8
X_5056_ _5056_/A vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__buf_6
XFILLER_0_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8815_ _8833_/B _8175_/Y _8725_/X vssd1 vssd1 vccd1 vccd1 _8815_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4392__B _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5214__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5214__B2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8746_ _8334_/A _8782_/A _8745_/X vssd1 vssd1 vccd1 vccd1 _8746_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5765__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5958_ _6059_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4909_ _4909_/A vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__buf_8
X_8677_ _8677_/A vssd1 vssd1 vccd1 vccd1 _8677_/X sky130_fd_sc_hd__buf_1
X_5889_ _5926_/B vssd1 vssd1 vccd1 vccd1 _5889_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7195__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8703__A2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7628_ _7378_/X _6059_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7628_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__6714__A1 _5659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7911__B1 _7918_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6714__B2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7559_ _6758_/B _7542_/A _7694_/A _5760_/Y vssd1 vssd1 vccd1 vccd1 _7559_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6190__A2 _7683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6112__B _6112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8219__A1 _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8219__B2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7690__A2 _6185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput301 sports_i[41] vssd1 vssd1 vccd1 vccd1 _7884_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__4567__B _7876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput312 sports_i[51] vssd1 vssd1 vccd1 vccd1 _8016_/A sky130_fd_sc_hd__clkbuf_1
Xinput323 sports_i[61] vssd1 vssd1 vccd1 vccd1 _8162_/A sky130_fd_sc_hd__clkbuf_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput334 sports_i[71] vssd1 vssd1 vccd1 vccd1 _7814_/B1 sky130_fd_sc_hd__clkbuf_4
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput345 sports_i[81] vssd1 vssd1 vccd1 vccd1 _7971_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7978__B1 _7985_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput356 sports_i[91] vssd1 vssd1 vccd1 vccd1 _8106_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7442__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6782__B _7171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6650__B1 _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5679__A _5679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__A _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5205__A1 _5208_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5205__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5756__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6953__A1 _6248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6303__A _6965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5508__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7902__B1 _7905_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _7155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7130__A1 _6697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6676__C _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7130__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8630__A1 _8358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7433__A2 _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8630__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6641__B1 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6930_ _6923_/X _6450_/X _6924_/X _6925_/Y _6929_/X vssd1 vssd1 vccd1 vccd1 _6930_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_107_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6861_ _6861_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6861_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7197__A1 _6002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7197__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8600_ _8309_/X _8581_/X _8313_/X _8583_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8600_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5812_ _5809_/Y _4886_/A _5810_/Y _4891_/A _5811_/Y vssd1 vssd1 vccd1 vccd1 _7171_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6792_ _7177_/A _6475_/X _5816_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6792_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5747__A2 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5743_ _5764_/A1 _4934_/A input48/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5743_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8531_ _8137_/X _8323_/X _8529_/X _8530_/Y vssd1 vssd1 vccd1 vccd1 _8531_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8412__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7309__A _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8462_ _8055_/Y _8567_/B _8497_/S _8461_/X vssd1 vssd1 vccd1 vccd1 _8462_/X sky130_fd_sc_hd__o211a_1
X_5674_ _6481_/B _5674_/B vssd1 vssd1 vccd1 vccd1 _5674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4625_ hold18/X _8759_/A vssd1 vssd1 vccd1 vccd1 _4626_/A sky130_fd_sc_hd__nor2_1
X_7413_ _7413_/A _7660_/B vssd1 vssd1 vccd1 vccd1 _7413_/X sky130_fd_sc_hd__and2_1
XFILLER_0_142_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8393_ _8441_/A _8349_/B _8555_/B vssd1 vssd1 vccd1 vccd1 _8393_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6172__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7344_ _5109_/B _7723_/B _7343_/X vssd1 vssd1 vccd1 vccd1 _7344_/Y sky130_fd_sc_hd__o21ai_1
X_4556_ _4595_/B _4612_/A _4612_/B vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__nand3_1
XANTENNA__6867__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6359__S _6359_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7275_ _7274_/X _7737_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7276_/A sky130_fd_sc_hd__mux2_1
X_4487_ hold36/A vssd1 vssd1 vccd1 vccd1 _8481_/S sky130_fd_sc_hd__clkinv_4
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5132__B1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6226_ _7705_/B vssd1 vssd1 vccd1 vccd1 _6948_/A sky130_fd_sc_hd__inv_2
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5683__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6880__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6157_ input2/X vssd1 vssd1 vccd1 vccd1 _6157_/Y sky130_fd_sc_hd__inv_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5108_/A _5108_/B vssd1 vssd1 vccd1 vccd1 _5108_/X sky130_fd_sc_hd__or2_1
XANTENNA__8621__A1 _8335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6088_ _6085_/X _6107_/A _6356_/S vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__mux2_2
X_5039_ input86/X _8271_/B input24/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__o22a_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5986__A2 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7188__A1 _5860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6107__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8385__B1 _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7188__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5199__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6935__A1 _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8729_ _7803_/Y _8820_/B _8829_/S vssd1 vssd1 vccd1 vccd1 _8729_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__8137__B1 _8142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8688__A1 _8203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8688__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6163__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5910__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4578__A _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7112__A1 _7470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5173__S _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7663__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8484__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput120 mports_i[207] vssd1 vssd1 vccd1 vccd1 _6007_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput131 mports_i[217] vssd1 vssd1 vccd1 vccd1 _6247_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5901__S _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput142 mports_i[227] vssd1 vssd1 vccd1 vccd1 _6400_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput153 mports_i[31] vssd1 vssd1 vccd1 vccd1 _5809_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8612__A1 _7867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput164 mports_i[41] vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__buf_2
Xinput175 mports_i[51] vssd1 vssd1 vccd1 vccd1 _6337_/B1 sky130_fd_sc_hd__clkbuf_2
Xinput186 mports_i[61] vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__clkbuf_2
Xinput197 mports_i[71] vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__buf_2
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5977__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6311__A1_N _6375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7179__A1 _6801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5856__B _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7129__A _7129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6968__A _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5872__A _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ _4504_/A _4611_/B _4504_/B vssd1 vssd1 vccd1 vccd1 _4456_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5390_ _5390_/A _6081_/S vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__nand2_1
Xoutput605 _5590_/X vssd1 vssd1 vccd1 vccd1 sports_o[193] sky130_fd_sc_hd__buf_12
XFILLER_0_151_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput616 _5851_/X vssd1 vssd1 vccd1 vccd1 sports_o[202] sky130_fd_sc_hd__buf_12
Xoutput627 _6146_/X vssd1 vssd1 vccd1 vccd1 sports_o[212] sky130_fd_sc_hd__buf_12
XFILLER_0_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput638 _6341_/X vssd1 vssd1 vccd1 vccd1 sports_o[222] sky130_fd_sc_hd__buf_12
X_4341_ _4341_/A _4341_/B vssd1 vssd1 vccd1 vccd1 _8239_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7103__A1 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput649 _7157_/X vssd1 vssd1 vccd1 vccd1 sports_o[27] sky130_fd_sc_hd__buf_12
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5114__B1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7060_ _7088_/A vssd1 vssd1 vccd1 vccd1 _7246_/B sky130_fd_sc_hd__buf_6
XFILLER_0_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6011_ _6089_/A1 _8709_/B input60/X _5091_/X vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__o22a_1
XANTENNA_hold26_A hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8603__A1 _7825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7406__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8603__B2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5417__A1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5417__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7311__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7962_ _7962_/A vssd1 vssd1 vccd1 vccd1 _7962_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5968__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6090__A1 _6020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6090__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6913_ _6913_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6913_/Y sky130_fd_sc_hd__nand2_1
X_7893_ _7881_/Y _7311_/A _7882_/Y _5230_/B _7892_/X vssd1 vssd1 vccd1 vccd1 _8333_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8423__A _8423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6844_ _6827_/A _5197_/X _8151_/B _6847_/A vssd1 vssd1 vccd1 vccd1 _6845_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6393__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8119__B1 _8119_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6775_ _6854_/A _5762_/B _5803_/A _6549_/A vssd1 vssd1 vccd1 vccd1 _6775_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8514_ _8117_/Y _8299_/X _8513_/Y _8304_/X _8496_/S vssd1 vssd1 vccd1 vccd1 _8514_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5726_ _6024_/A _6756_/B vssd1 vssd1 vccd1 vccd1 _5749_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8445_ _8445_/A vssd1 vssd1 vccd1 vccd1 _8445_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6145__A2 _6908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5657_ _5651_/X _5656_/Y _6926_/A vssd1 vssd1 vccd1 vccd1 _5657_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4608_ _6102_/B _4841_/B vssd1 vssd1 vccd1 vccd1 _4608_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5588_ _5575_/A _8491_/B _5576_/A _4933_/A _5587_/X vssd1 vssd1 vccd1 vccd1 _5645_/A
+ sky130_fd_sc_hd__o221a_4
X_8376_ _8376_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8376_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7893__A2 _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7327_ _7027_/A _7349_/A _6461_/A _7753_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7327_/X
+ sky130_fd_sc_hd__a221o_1
X_4539_ _8942_/A _4535_/Y _4586_/A vssd1 vssd1 vccd1 vccd1 _4863_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7258_ _6310_/X _7026_/X _7257_/X vssd1 vssd1 vccd1 vccd1 _7258_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5656__A1 _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6853__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6209_ _6209_/A _6870_/S vssd1 vssd1 vccd1 vccd1 _6209_/Y sky130_fd_sc_hd__nand2_1
X_7189_ _6827_/A _7023_/X _7188_/X vssd1 vssd1 vccd1 vccd1 _7189_/X sky130_fd_sc_hd__o21a_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8070__A2 _8491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5022__A _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8333__A _8333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6384__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6136__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7333__A1 _7328_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6788__A _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8530__B1 _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5895__A1 _5853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5895__B2 _5885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6844__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8597__B1 _8303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8061__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6028__A _6028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output506_A _6954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5867__A _5867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4890_ _4890_/A vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7572__A1 _5772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6560_ _6854_/A _6560_/B vssd1 vssd1 vccd1 vccd1 _6560_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5511_ _5511_/A vssd1 vssd1 vccd1 vccd1 _5511_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_109_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6491_ _6491_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6491_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6127__A2 _7660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8521__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5442_ _5274_/X input99/X _5275_/X input37/X vssd1 vssd1 vccd1 vccd1 _5442_/Y sky130_fd_sc_hd__a22oi_1
X_8230_ _8696_/B vssd1 vssd1 vccd1 vccd1 _8230_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput402 _8830_/X vssd1 vssd1 vccd1 vccd1 mports_o[132] sky130_fd_sc_hd__buf_12
XANTENNA__5886__A1 _5928_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5886__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput413 _7794_/X vssd1 vssd1 vccd1 vccd1 mports_o[1] sky130_fd_sc_hd__buf_12
XFILLER_0_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput424 _7805_/X vssd1 vssd1 vccd1 vccd1 mports_o[2] sky130_fd_sc_hd__buf_12
X_5373_ _6628_/B _5364_/Y _5372_/Y vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__o21ai_1
X_8161_ _8161_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _8161_/Y sky130_fd_sc_hd__nand2_1
Xoutput435 _7816_/X vssd1 vssd1 vccd1 vccd1 mports_o[3] sky130_fd_sc_hd__buf_12
XFILLER_0_22_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput446 _7839_/X vssd1 vssd1 vccd1 vccd1 mports_o[4] sky130_fd_sc_hd__buf_12
Xoutput457 _7863_/X vssd1 vssd1 vccd1 vccd1 mports_o[5] sky130_fd_sc_hd__buf_12
X_7112_ _7470_/A _7026_/X _7110_/X _7111_/X vssd1 vssd1 vccd1 vccd1 _7112_/X sky130_fd_sc_hd__o22a_2
X_4324_ _8160_/A _4591_/B _6231_/C vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__8824__A1 _8211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8285__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput468 _7880_/X vssd1 vssd1 vccd1 vccd1 mports_o[6] sky130_fd_sc_hd__buf_12
X_8092_ _8511_/A _7954_/X _8091_/Y _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8092_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput479 _7895_/X vssd1 vssd1 vccd1 vccd1 mports_o[7] sky130_fd_sc_hd__buf_12
XANTENNA__5638__A1 _5596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7043_ _8919_/A _7043_/B vssd1 vssd1 vccd1 vccd1 _7043_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4665__B _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8588__B1 _7771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8052__A2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7945_ _7935_/Y _7874_/X _7936_/Y _7875_/X _7944_/Y vssd1 vssd1 vccd1 vccd1 _7945_/Y
+ sky130_fd_sc_hd__a221oi_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7876_ _7876_/A vssd1 vssd1 vccd1 vccd1 _7876_/X sky130_fd_sc_hd__buf_8
XFILLER_0_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6827_ _6827_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6827_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6366__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7563__B2 _7562_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6758_ _6841_/A _6758_/B vssd1 vssd1 vccd1 vccd1 _6758_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5709_ _7532_/B vssd1 vssd1 vccd1 vccd1 _7148_/A sky130_fd_sc_hd__inv_2
XFILLER_0_150_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6689_ _5560_/Y _6666_/Y _6689_/S vssd1 vssd1 vccd1 vccd1 _7483_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8428_ _8427_/Y _8403_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8428_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7866__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8359_ _8359_/A _8455_/B vssd1 vssd1 vccd1 vccd1 _8359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5017__A _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7079__B1 _5280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8276__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7618__A2 _5923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5629__A1 _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6826__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8762__S _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8043__A2 _8042_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8958__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5801__A1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7003__B1 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6357__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7554__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5565__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8510__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7857__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5868__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output456_A _8528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7609__A2 _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6965__B _6965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6293__A1 _6326_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6293__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6045__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5991_ _5988_/Y _4886_/A _5989_/Y _4891_/A _5990_/Y vssd1 vssd1 vccd1 vccd1 _6046_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__7793__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6596__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7730_ _7728_/Y _7332_/A _7729_/Y vssd1 vssd1 vccd1 vccd1 _7730_/Y sky130_fd_sc_hd__a21oi_2
X_4942_ input1/X _4930_/X _4888_/A _4933_/X _4941_/X vssd1 vssd1 vccd1 vccd1 _4942_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7661_ _6912_/A _7680_/B _7659_/X _7640_/B _7660_/X vssd1 vssd1 vccd1 vccd1 _7661_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6348__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4873_ _5091_/A vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__buf_6
XFILLER_0_129_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8742__B1 _7871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7545__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6612_ _8924_/B _5362_/Y _6611_/Y vssd1 vssd1 vccd1 vccd1 _6613_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5556__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6753__C1 _6752_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7592_ _7592_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _7592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6543_ _6543_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6474_ _6474_/A vssd1 vssd1 vccd1 vccd1 _7032_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5859__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5859__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8213_ _7975_/X _8200_/X _8207_/X _8212_/Y vssd1 vssd1 vccd1 vccd1 _8213_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5425_ _7829_/A _6231_/C _5425_/C vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__or3_1
XANTENNA__6520__A2 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8144_ _8148_/A1 _6456_/B _8139_/Y _8141_/Y _8143_/Y vssd1 vssd1 vccd1 vccd1 _8145_/A
+ sky130_fd_sc_hd__o221ai_2
X_5356_ _6212_/A _5356_/B vssd1 vssd1 vccd1 vccd1 _5356_/X sky130_fd_sc_hd__or2_1
XANTENNA__6875__B _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6808__B1 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4307_ _4300_/Y _4305_/Y _4406_/A vssd1 vssd1 vccd1 vccd1 _4307_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8273__A2 _8235_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8075_ _8080_/A1 _5145_/A _8080_/B1 _5616_/A vssd1 vssd1 vccd1 vccd1 _8075_/Y sky130_fd_sc_hd__o22ai_2
X_5287_ _6284_/A _6578_/B _5762_/A _5264_/Y _5286_/X vssd1 vssd1 vccd1 vccd1 _5288_/A
+ sky130_fd_sc_hd__o221ai_4
X_7026_ _7138_/A vssd1 vssd1 vccd1 vccd1 _7026_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8025__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6891__A _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6036__A1 _6061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6036__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8977_ _8979_/CLK _8977_/D input229/X vssd1 vssd1 vccd1 vccd1 _8977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7784__A1 _7791_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7784__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4598__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7928_ _7931_/A1 _5780_/X _7931_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7928_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6115__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7859_ _8194_/A _7859_/B vssd1 vssd1 vccd1 vccd1 _7859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5547__B1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6830__S _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5446__S _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7227__A _7227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7839__A2 _7821_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6275__A1 _6309_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6275__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7472__B1 _5464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8492__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6027__A1 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6027__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7775__A1 _7765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7775__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5786__B1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5210__A _5359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5250__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7527__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6750__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7137__A _7137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6502__A2 _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5210_ _5359_/A vssd1 vssd1 vccd1 vccd1 _7013_/A sky130_fd_sc_hd__buf_12
X_6190_ _5741_/B _7683_/A _6189_/Y _5125_/X vssd1 vssd1 vccd1 vccd1 _6190_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6695__B _6695_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5141_ _4893_/A input87/X _4896_/A input25/X vssd1 vssd1 vccd1 vccd1 _5141_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_86_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8255__A2 _8222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5072_ _8713_/C input85/X _8579_/C input22/X vssd1 vssd1 vccd1 vccd1 _5072_/Y sky130_fd_sc_hd__a22oi_1
X_8900_ _8899_/Y _4800_/A _8880_/Y vssd1 vssd1 vccd1 vccd1 _8903_/A sky130_fd_sc_hd__a21o_1
XANTENNA__8007__A2 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6018__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8831_ _8833_/B _8235_/Y _8725_/X vssd1 vssd1 vccd1 vccd1 _8831_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8762_ _8760_/X _7945_/Y _8788_/S vssd1 vssd1 vccd1 vccd1 _8762_/X sky130_fd_sc_hd__mux2_1
X_5974_ _8140_/A _5870_/Y _5973_/Y vssd1 vssd1 vccd1 vccd1 _6837_/B sky130_fd_sc_hd__o21a_2
XANTENNA__4662__C _4662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5241__A2 _6567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7713_ _8755_/C _5299_/B _7246_/A _7712_/Y vssd1 vssd1 vccd1 vccd1 _7713_/X sky130_fd_sc_hd__a31o_1
X_4925_ _4925_/A vssd1 vssd1 vccd1 vccd1 _6356_/S sky130_fd_sc_hd__buf_8
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8693_ _8255_/X _8584_/B hold21/A _8698_/B _8692_/X vssd1 vssd1 vccd1 vccd1 _8693_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__7518__A1 _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7644_ _7378_/X _6058_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7646_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4856_ _8929_/A vssd1 vssd1 vccd1 vccd1 _4857_/B sky130_fd_sc_hd__inv_2
XANTENNA__8191__A1 _8187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8191__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8150__B _8150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7575_ _7575_/A _7575_/B vssd1 vssd1 vccd1 vccd1 _7575_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4787_ _4787_/A vssd1 vssd1 vccd1 vccd1 _4789_/A sky130_fd_sc_hd__inv_2
XANTENNA__6741__A2 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6526_ _6526_/A vssd1 vssd1 vccd1 vccd1 _7366_/B sky130_fd_sc_hd__inv_2
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6457_ _6470_/A _7829_/A vssd1 vssd1 vccd1 vccd1 _6457_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8962__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5408_ _6645_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5408_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5701__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6388_ _6388_/A1 _4930_/X input15/X _4933_/X _6387_/X vssd1 vssd1 vccd1 vccd1 _7750_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8127_ _8132_/A1 _5146_/A _8132_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _8127_/Y sky130_fd_sc_hd__o22ai_2
X_5339_ _5274_/A input96/X _5275_/A input33/X vssd1 vssd1 vccd1 vccd1 _5339_/Y sky130_fd_sc_hd__a22oi_2
XANTENNA__8246__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8651__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8058_ _8058_/A vssd1 vssd1 vccd1 vccd1 _8058_/Y sky130_fd_sc_hd__inv_2
X_7009_ _4876_/X _7004_/X _4899_/Y _7088_/A vssd1 vssd1 vccd1 vccd1 _7009_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6009__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5480__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4853__B _8976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5965__A _5965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4991__A1 _4978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4991__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8237__A2 _8226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8973__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6248__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7445__B1 _7372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7996__B2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8516__A _8516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output419_A _8135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7748__A1 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5223__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5875__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4710_ _4710_/A _8239_/A vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_155_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5690_ _5690_/A _6081_/S vssd1 vssd1 vccd1 vccd1 _5691_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4641_ hold31/A hold30/A vssd1 vssd1 vccd1 vccd1 _4934_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7920__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6723__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7360_ _7673_/A vssd1 vssd1 vccd1 vccd1 _7476_/B sky130_fd_sc_hd__inv_2
X_4572_ _7778_/B _5229_/A _4560_/Y _5230_/B _4571_/Y vssd1 vssd1 vccd1 vccd1 _4607_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_142_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6311_ _6375_/B _6312_/B _6261_/A _6310_/X vssd1 vssd1 vccd1 vccd1 _6311_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7291_ _7291_/A vssd1 vssd1 vccd1 vccd1 _7291_/X sky130_fd_sc_hd__buf_1
XANTENNA__5814__S _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6242_ _8444_/A _6248_/A1 _8257_/C input5/X vssd1 vssd1 vccd1 vccd1 _6242_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_122_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8228__A2 _8234_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6173_ _7696_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6173_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6239__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5124_ _7356_/B _8857_/B _5359_/B _7345_/B _5123_/Y vssd1 vssd1 vccd1 vccd1 _5124_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7987__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5055_/A vssd1 vssd1 vccd1 vccd1 _6304_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7739__A1 _6349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7739__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8814_ _8137_/X _8806_/B _8812_/X _8813_/Y vssd1 vssd1 vccd1 vccd1 _8814_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5214__A2 _5211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8745_ _7888_/Y _8738_/A _7890_/Y _8711_/A _8824_/S vssd1 vssd1 vccd1 vccd1 _8745_/X
+ sky130_fd_sc_hd__a221o_1
X_5957_ _5965_/A _4929_/A _5966_/A _4933_/A _5956_/X vssd1 vssd1 vccd1 vccd1 _6059_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4908_ _4876_/X _6234_/B _4899_/Y _5128_/A vssd1 vssd1 vccd1 vccd1 _4908_/X sky130_fd_sc_hd__a22o_1
X_8676_ _8675_/X _8523_/A _8690_/S vssd1 vssd1 vccd1 vccd1 _8677_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8164__A1 _8175_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5888_ _5885_/X _7316_/A _8194_/A _5899_/A vssd1 vssd1 vccd1 vccd1 _5926_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7627_ _7590_/A _7618_/Y _7619_/Y _7626_/X vssd1 vssd1 vccd1 vccd1 _7627_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__6175__B1 _6158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4839_ _4839_/A _4839_/B vssd1 vssd1 vccd1 vccd1 _4839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7911__A1 _7918_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6714__A2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7911__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5922__B1 _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7558_ _7558_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _7558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6509_ _5123_/B _6450_/X _6508_/X vssd1 vssd1 vccd1 vccd1 _6509_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7489_ _7542_/A _5500_/X _7326_/A vssd1 vssd1 vccd1 vccd1 _7489_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7505__A _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7224__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8219__A2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput302 sports_i[42] vssd1 vssd1 vccd1 vccd1 _7897_/A sky130_fd_sc_hd__buf_1
Xinput313 sports_i[52] vssd1 vssd1 vccd1 vccd1 _8031_/A sky130_fd_sc_hd__clkbuf_1
Xinput324 sports_i[62] vssd1 vssd1 vccd1 vccd1 _8196_/B1 sky130_fd_sc_hd__buf_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkbuf_4
Xinput335 sports_i[72] vssd1 vssd1 vccd1 vccd1 _7836_/A sky130_fd_sc_hd__buf_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7978__A1 _7985_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7978__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput346 sports_i[82] vssd1 vssd1 vccd1 vccd1 _7985_/B1 sky130_fd_sc_hd__buf_2
Xinput357 sports_i[92] vssd1 vssd1 vccd1 vccd1 _8119_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7240__A _7240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6650__A1 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__B _4909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5205__A2 _4927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4964__A1 _4963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8155__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7902__A1 _7905_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7902__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 _7155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7415__A _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7666__B1 _7372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4758__B _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7130__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5141__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__B2 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7969__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6465__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8630__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4774__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6641__A1 _7459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6641__B2 _6635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6860_ _6868_/A vssd1 vssd1 vccd1 vccd1 _6861_/A sky130_fd_sc_hd__inv_2
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7197__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5811_ _5274_/X _5825_/A1 _5275_/X input51/X vssd1 vssd1 vccd1 vccd1 _5811_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6791_ _6786_/X _6450_/X _6787_/Y _6788_/X _6790_/X vssd1 vssd1 vccd1 vccd1 _6791_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8530_ _8153_/X _8518_/B _8572_/S vssd1 vssd1 vccd1 vccd1 _8530_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4955__A1 _4956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5742_ _5125_/X _5720_/X _5739_/X _5740_/X _5741_/X vssd1 vssd1 vccd1 vccd1 _5742_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__4955__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8461_ _8457_/Y _8304_/A _8460_/Y _8299_/A _8496_/S vssd1 vssd1 vccd1 vccd1 _8461_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7309__B _7309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8697__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5673_ _5909_/B _7514_/A _5011_/Y _5660_/Y _5672_/Y vssd1 vssd1 vccd1 vccd1 _5673_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7412_ _5280_/A _7668_/B _5285_/X _7638_/B vssd1 vssd1 vccd1 vccd1 _7412_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4624_ _4593_/Y _4619_/Y _8926_/S vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_154_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8392_ _8392_/A vssd1 vssd1 vccd1 vccd1 _8441_/A sky130_fd_sc_hd__inv_2
XFILLER_0_114_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5380__A1 _5337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7343_ _6488_/A _7349_/A _7043_/Y _7753_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7343_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5380__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4555_ _4534_/B _4839_/B _4839_/A vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7325__A _7334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7274_ _4793_/A _7138_/X _7272_/X _7273_/X vssd1 vssd1 vccd1 vccd1 _7274_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4486_ _5077_/A vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__inv_6
X_6225_ _6225_/A vssd1 vssd1 vccd1 vccd1 _6225_/X sky130_fd_sc_hd__buf_1
XANTENNA__5132__B2 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6880__A1 _6867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6156_ _6156_/A vssd1 vssd1 vccd1 vccd1 _6156_/Y sky130_fd_sc_hd__inv_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6880__B2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5109_/B _5230_/B _7536_/B _6507_/B _5106_/Y vssd1 vssd1 vccd1 vccd1 _5108_/B
+ sky130_fd_sc_hd__a221o_1
X_6087_ _6020_/A _8271_/A _6021_/A _5191_/X _6086_/X vssd1 vssd1 vccd1 vccd1 _6107_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__7060__A _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5038_ _5070_/A _8335_/B _5071_/A _4913_/A _5037_/X vssd1 vssd1 vccd1 vccd1 _5109_/B
+ sky130_fd_sc_hd__o221a_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7188__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5199__A1 _5105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6396__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5199__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6989_ _6367_/B _6989_/B vssd1 vssd1 vccd1 vccd1 _6989_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_76_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6935__A2 _6212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8728_ _7798_/X _8803_/B _7800_/X _8711_/X _8820_/B vssd1 vssd1 vccd1 vccd1 _8728_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6404__A _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8137__A1 _8148_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8137__B2 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8659_ _8698_/B _8068_/Y _8590_/X vssd1 vssd1 vccd1 vccd1 _8659_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_91_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8976__D _8976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7112__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput110 mports_i[199] vssd1 vssd1 vccd1 vccd1 _5764_/A1 sky130_fd_sc_hd__buf_2
Xinput121 mports_i[208] vssd1 vssd1 vccd1 vccd1 _6031_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput132 mports_i[218] vssd1 vssd1 vccd1 vccd1 _6262_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput143 mports_i[22] vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__clkbuf_4
Xinput154 mports_i[32] vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8612__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput165 mports_i[42] vssd1 vssd1 vccd1 vccd1 _6141_/A1 sky130_fd_sc_hd__buf_2
Xinput176 mports_i[52] vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__clkbuf_1
Xinput187 mports_i[62] vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__clkbuf_2
Xinput198 mports_i[72] vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__buf_2
XFILLER_0_59_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7179__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6387__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6314__A _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8128__B2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6139__B1 _6158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7887__B1 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput606 _5650_/X vssd1 vssd1 vccd1 vccd1 sports_o[194] sky130_fd_sc_hd__buf_12
XFILLER_0_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput617 _5894_/X vssd1 vssd1 vccd1 vccd1 sports_o[203] sky130_fd_sc_hd__buf_12
Xoutput628 _6191_/X vssd1 vssd1 vccd1 vccd1 sports_o[213] sky130_fd_sc_hd__buf_12
XFILLER_0_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8836__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _4340_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4341_/B sky130_fd_sc_hd__nand2_1
Xoutput639 _6347_/X vssd1 vssd1 vccd1 vccd1 sports_o[223] sky130_fd_sc_hd__buf_12
XFILLER_0_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5114__A1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5114__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6311__B1 _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6010_ _5031_/X _5923_/A _6006_/Y _6009_/X vssd1 vssd1 vccd1 vccd1 _6010_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6862__A1 _5923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8064__B1 _8067_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8603__A2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5417__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6614__A1 _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7811__B1 _7814_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6614__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7961_ _7760_/X _8369_/A _7957_/X _7960_/X vssd1 vssd1 vccd1 vccd1 _7961_/X sky130_fd_sc_hd__a22o_2
XANTENNA__6090__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6912_ _6912_/A _6912_/B vssd1 vssd1 vccd1 vccd1 _6912_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7892_ _7874_/A _7883_/Y _4597_/A _7884_/Y vssd1 vssd1 vccd1 vccd1 _7892_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8367__A1 _8366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6843_ _6843_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6843_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6378__B1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8423__B _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6917__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8119__A1 _8119_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6774_ _7167_/A _6475_/A _5754_/Y _6694_/B vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8119__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8513_ _8540_/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8513_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5725_ _5722_/Y _4885_/A _5723_/Y _4890_/A _5724_/Y vssd1 vssd1 vccd1 vccd1 _6756_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7327__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8444_ _8444_/A _8444_/B vssd1 vssd1 vccd1 vccd1 _8445_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5656_ _8842_/B _5654_/Y _7529_/B vssd1 vssd1 vccd1 vccd1 _5656_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7342__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5782__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4607_ _4607_/A _4607_/B vssd1 vssd1 vccd1 vccd1 _4841_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_115_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8375_ _8375_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8375_/Y sky130_fd_sc_hd__nand2_1
X_5587_ _5587_/A1 _8368_/A input41/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7326_ _7326_/A vssd1 vssd1 vccd1 vccd1 _7723_/B sky130_fd_sc_hd__buf_6
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8827__C1 _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4538_ _4538_/A vssd1 vssd1 vccd1 vccd1 _4586_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7257_ _6277_/A _7004_/X _6303_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7257_/X
+ sky130_fd_sc_hd__a221o_1
X_4469_ _8166_/A _4466_/Y hold23/A _4468_/Y vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__o211ai_2
X_6208_ _6207_/Y _6173_/Y _8150_/A vssd1 vssd1 vccd1 vccd1 _6209_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6853__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7188_ _5860_/A _7004_/X _5930_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7188_/X
+ sky130_fd_sc_hd__a221o_1
X_6139_ input2/X _4932_/A _6158_/A _4929_/A _6138_/X vssd1 vssd1 vccd1 vccd1 _6185_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6605__A1 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7802__B1 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6118__B _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6369__B1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7030__A1 _7332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4919__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4919__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7333__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8530__A1 _8153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6788__B _6788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5344__A1 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5895__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7097__A1 _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6844__A1 _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6844__B2 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8597__A1 _7800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8597__B2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7021__A1 _6440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7021__B2 _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5032__B1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5510_ _5510_/A vssd1 vssd1 vccd1 vccd1 _5510_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6490_ _6488_/Y _7043_/B _6994_/B vssd1 vssd1 vccd1 vccd1 _6491_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_70_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5441_ _5441_/A vssd1 vssd1 vccd1 vccd1 _5441_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6532__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput403 _8834_/X vssd1 vssd1 vccd1 vccd1 mports_o[133] sky130_fd_sc_hd__buf_12
XANTENNA__5886__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput414 _8070_/X vssd1 vssd1 vccd1 vccd1 mports_o[20] sky130_fd_sc_hd__buf_12
X_8160_ _8160_/A _8172_/B vssd1 vssd1 vccd1 vccd1 _8161_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput425 _8224_/X vssd1 vssd1 vccd1 vccd1 mports_o[30] sky130_fd_sc_hd__buf_12
X_5372_ _5372_/A _6926_/A vssd1 vssd1 vccd1 vccd1 _5372_/Y sky130_fd_sc_hd__nand2_1
Xoutput436 _8326_/X vssd1 vssd1 vccd1 vccd1 mports_o[40] sky130_fd_sc_hd__buf_12
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput447 _8422_/X vssd1 vssd1 vccd1 vccd1 mports_o[50] sky130_fd_sc_hd__buf_12
X_7111_ _5465_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7111_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8285__B1 _7811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput458 _8531_/X vssd1 vssd1 vccd1 vccd1 mports_o[60] sky130_fd_sc_hd__buf_12
X_4323_ _4337_/A vssd1 vssd1 vccd1 vccd1 _8160_/A sky130_fd_sc_hd__buf_8
Xoutput469 _8599_/X vssd1 vssd1 vccd1 vccd1 mports_o[70] sky130_fd_sc_hd__buf_12
X_8091_ _8084_/Y _6500_/X _8085_/Y _7769_/X _8090_/Y vssd1 vssd1 vccd1 vccd1 _8091_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5099__B1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7042_ _7042_/A vssd1 vssd1 vccd1 vccd1 _7042_/X sky130_fd_sc_hd__buf_1
XFILLER_0_129_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4846__B1 hold4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8588__A1 _7765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5123__A _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8588__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7749__S _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7944_ _7944_/A1 _7876_/X _7944_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7944_/Y sky130_fd_sc_hd__o22ai_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7875_ _8174_/A vssd1 vssd1 vccd1 vccd1 _7875_/X sky130_fd_sc_hd__buf_12
XFILLER_0_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6826_ _6825_/X _6899_/B _6968_/A vssd1 vssd1 vccd1 vccd1 _6826_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8760__A1 _7942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6757_ _6432_/X _6756_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6757_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5708_ _6084_/B _6727_/B _5707_/Y _5096_/A _6356_/S vssd1 vssd1 vccd1 vccd1 _5708_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6688_ _6686_/X _6933_/A _6968_/A _6687_/X vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5326__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8427_ _8427_/A _8455_/B vssd1 vssd1 vccd1 vccd1 _8427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_104_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5326__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5639_ _5655_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8358_ _8358_/A _8455_/B vssd1 vssd1 vccd1 vccd1 _8358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7079__A1 _7413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7079__B2 _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7309_ _7510_/B _7309_/B vssd1 vssd1 vccd1 vccd1 _7389_/A sky130_fd_sc_hd__nor2_8
XANTENNA__8815__A2 _8175_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8289_ _8497_/S vssd1 vssd1 vccd1 vccd1 _8349_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5801__A2 _5786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4591__B _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7539__C1 _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7003__A1 _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8200__B1 _8210_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7003__B2 _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5014__B1 _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8751__A1 _8372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7554__A2 _5744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5565__A1 _5562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5565__B2 _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5868__A2 _5928_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8519__A _8519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output449_A _8450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6293__A2 _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7490__A1 _5558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _5274_/X _6061_/A1 _5275_/X input59/X vssd1 vssd1 vccd1 vccd1 _5990_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__5253__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7793__A2 _8272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4941_ input80/X _8706_/B input17/X _4940_/X vssd1 vssd1 vccd1 vccd1 _4941_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7660_ _7660_/A _7660_/B vssd1 vssd1 vccd1 vccd1 _7660_/X sky130_fd_sc_hd__and2_1
X_4872_ _5090_/A vssd1 vssd1 vccd1 vccd1 _8310_/B sky130_fd_sc_hd__buf_6
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5005__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8742__A1 _7869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7545__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8742__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6611_ _6611_/A _8924_/B vssd1 vssd1 vccd1 vccd1 _6611_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7591_ _6820_/Y _7619_/B _7587_/X _7589_/Y _7590_/Y vssd1 vssd1 vccd1 vccd1 _7591_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6542_ _6542_/A _6933_/A vssd1 vssd1 vccd1 vccd1 _6542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7317__B _7372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6473_ _6473_/A vssd1 vssd1 vccd1 vccd1 _6694_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5859__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8212_ _8211_/Y _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _8212_/Y sky130_fd_sc_hd__a21oi_1
X_5424_ _5425_/C vssd1 vssd1 vccd1 vccd1 _7451_/A sky130_fd_sc_hd__inv_2
XFILLER_0_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8143_ _8163_/A _8143_/B vssd1 vssd1 vccd1 vccd1 _8143_/Y sky130_fd_sc_hd__nand2_1
X_5355_ _6621_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _5355_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8429__A _8429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4306_ hold4/X vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__inv_2
X_8074_ _8071_/Y _7013_/A _8072_/Y _5117_/A _8073_/Y vssd1 vssd1 vccd1 vccd1 _8476_/A
+ sky130_fd_sc_hd__a221oi_4
X_5286_ _5013_/Y _5269_/Y _5285_/X _5997_/B vssd1 vssd1 vccd1 vccd1 _5286_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7481__A1 _6679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7025_ _4966_/X _7097_/S _7021_/X _7024_/X vssd1 vssd1 vccd1 vccd1 _7025_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5492__B1 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7685__A1_N _7364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6891__B _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6036__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7233__A1 _7696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8976_ _8976_/CLK _8976_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__7784__A2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4598__A2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7927_ _7922_/Y _6024_/A _7923_/Y _6411_/A _7926_/Y vssd1 vssd1 vccd1 vccd1 _8359_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7858_ _8198_/A _7858_/B vssd1 vssd1 vccd1 vccd1 _7858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5547__A1 _5557_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6809_ _6852_/A _6809_/B vssd1 vssd1 vccd1 vccd1 _6809_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5547__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7789_ _7786_/X _7768_/X _7788_/X _7772_/X _7774_/X vssd1 vssd1 vccd1 vccd1 _7789_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6412__A _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8249__B1 _8252_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5970__B _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4867__A _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4586__B _4793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6275__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7472__B2 _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8421__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5235__B1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7775__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6983__A0 _6982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5786__A1 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5786__B2 _6758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7527__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output399_A _7961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6322__A _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8488__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5140_ _5140_/A vssd1 vssd1 vccd1 vccd1 _5140_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5071_ _5071_/A vssd1 vssd1 vccd1 vccd1 _5071_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7215__A1 _6112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8830_ _8830_/A vssd1 vssd1 vccd1 vccd1 _8830_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_126_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5401__A _5401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8761_ _8824_/S vssd1 vssd1 vccd1 vccd1 _8788_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__5777__A1 _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5973_ _6080_/A _6839_/B _8140_/A vssd1 vssd1 vccd1 vccd1 _5973_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7712_ _7532_/A _6257_/A _7348_/A vssd1 vssd1 vccd1 vccd1 _7712_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4924_ _6212_/A _5108_/A vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__nand2_2
X_8692_ _8217_/X _8581_/A _8219_/X _8583_/A vssd1 vssd1 vccd1 vccd1 _8692_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7518__A2 _5679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5529__A1 _5543_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7643_ _7637_/X _7640_/Y _7641_/X _7642_/X vssd1 vssd1 vccd1 vccd1 _7643_/X sky130_fd_sc_hd__a31o_2
XANTENNA__5529__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4855_ _4855_/A _4863_/C vssd1 vssd1 vccd1 vccd1 _8929_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6726__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8191__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7574_ _7172_/A _7630_/B _5814_/X _7638_/B vssd1 vssd1 vccd1 vccd1 _7574_/X sky130_fd_sc_hd__a22o_1
X_4786_ _4786_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6525_ _6525_/A _6933_/A vssd1 vssd1 vccd1 vccd1 _6525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6456_ _6456_/A _6456_/B vssd1 vssd1 vccd1 vccd1 _6470_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7151__A0 _7150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6886__B _6940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8056__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5407_ _5342_/X _7450_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6645_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5701__A1 _6732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6387_ _6387_/A1 _8706_/B input77/X _4940_/X vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8159__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5701__B2 _7544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8126_ _8123_/Y _7761_/A _8124_/Y _5117_/A _8125_/Y vssd1 vssd1 vccd1 vccd1 _8523_/A
+ sky130_fd_sc_hd__a221oi_4
X_5338_ _5338_/A vssd1 vssd1 vccd1 vccd1 _5338_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8057_ _7975_/X _8451_/A _8053_/X _8056_/X vssd1 vssd1 vccd1 vccd1 _8057_/X sky130_fd_sc_hd__a22o_4
XANTENNA__7454__B2 _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5269_ _6304_/A _6576_/B _5011_/A vssd1 vssd1 vccd1 vccd1 _5269_/Y sky130_fd_sc_hd__o21ai_1
X_7008_ _7008_/A vssd1 vssd1 vccd1 vccd1 _7088_/A sky130_fd_sc_hd__buf_4
XANTENNA__6009__A2 _6868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7510__B _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7206__A1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7757__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8959_ _8978_/CLK _8959_/D fanout732/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4991__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8768__S _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7142__A0 _7141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6288__S _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8890__B1 _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7500__A1_N _5562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6248__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7445__A1 _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7996__A2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7701__A _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8516__B _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8152__A2_N _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5875__B _6809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output683_A _6452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6708__B1 _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4640_ _8264_/A vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__inv_8
XFILLER_0_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7920__A2 _8335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4571_ _5106_/A _4569_/X _4570_/X vssd1 vssd1 vccd1 vccd1 _4571_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6310_ _6299_/A _8516_/B input8/X _4913_/X _6309_/X vssd1 vssd1 vccd1 vccd1 _6310_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7290_ _7289_/X _7750_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7291_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8330__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6241_ _6248_/A1 _8480_/B input5/X _4870_/X _6240_/X vssd1 vssd1 vccd1 vccd1 _6241_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6198__S _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7684__B2 _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5695__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _8978_/CLK sky130_fd_sc_hd__clkbuf_16
X_6172_ _6183_/A1 _5102_/A input3/X _5191_/A _6171_/X vssd1 vssd1 vccd1 vccd1 _7696_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6239__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5123_ _5123_/A _5123_/B vssd1 vssd1 vccd1 vccd1 _5123_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__8633__B1 _7969_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7987__A2 _8772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5054_ _5145_/A vssd1 vssd1 vccd1 vccd1 _5171_/B sky130_fd_sc_hd__inv_8
XANTENNA__7739__A2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8397__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8813_ _8153_/X _8820_/B _8829_/S vssd1 vssd1 vccd1 vccd1 _8813_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6661__S _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5956_ _6031_/A1 _8368_/A input58/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5956_/X sky130_fd_sc_hd__o22a_1
X_8744_ _7867_/Y _8806_/B _8742_/X _8743_/X vssd1 vssd1 vccd1 vccd1 _8744_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_137_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8149__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4907_ _4974_/A _6367_/A vssd1 vssd1 vccd1 vccd1 _5128_/A sky130_fd_sc_hd__nor2_8
X_8675_ _8674_/X _8133_/Y _8689_/S vssd1 vssd1 vccd1 vccd1 _8675_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5887_ _5866_/A _5111_/A _5867_/A _4931_/A _5886_/X vssd1 vssd1 vccd1 vccd1 _5899_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8161__B _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8164__A2 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4838_ _4802_/A _4803_/A _8904_/B vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__o21a_1
X_7626_ _6871_/A _7361_/X _7624_/X _7754_/A _7625_/X vssd1 vssd1 vccd1 vccd1 _7626_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6175__B2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7911__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5922__A1 _5931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7557_ _6767_/Y _7619_/B _7553_/X _7555_/Y _7556_/Y vssd1 vssd1 vccd1 vccd1 _7557_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6897__A _6897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4769_ _4792_/B _4800_/B vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7492__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6508_ _6503_/X _6467_/X _7001_/S _6505_/Y _6507_/Y vssd1 vssd1 vccd1 vccd1 _6508_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7488_ _7488_/A _7680_/B vssd1 vssd1 vccd1 vccd1 _7488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6478__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7505__B _7505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7675__A1 _6102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5135__C1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6439_ _6841_/A _6440_/A vssd1 vssd1 vccd1 vccd1 _6439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8109_ _7975_/X _8499_/A _8105_/X _8108_/X vssd1 vssd1 vccd1 vccd1 _8109_/X sky130_fd_sc_hd__a22o_2
Xinput303 sports_i[43] vssd1 vssd1 vccd1 vccd1 _7910_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8624__B1 _8362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkbuf_4
Xinput314 sports_i[53] vssd1 vssd1 vccd1 vccd1 _8046_/A sky130_fd_sc_hd__clkbuf_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput325 sports_i[63] vssd1 vssd1 vccd1 vccd1 _8210_/B1 sky130_fd_sc_hd__clkbuf_2
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__buf_2
Xinput336 sports_i[73] vssd1 vssd1 vccd1 vccd1 _7841_/A sky130_fd_sc_hd__buf_1
XANTENNA__7978__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput347 sports_i[83] vssd1 vssd1 vccd1 vccd1 _7998_/B1 sky130_fd_sc_hd__clkbuf_4
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput358 sports_i[93] vssd1 vssd1 vccd1 vccd1 _8132_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__6650__A2 _7459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5041__A _6507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4880__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8352__A _8352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8155__A2 _8137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7902__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _7174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7666__A1 _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8863__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5677__B1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5141__A2 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7969__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7431__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8091__B2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6641__A2 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6047__A _6047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5810_ _5810_/A vssd1 vssd1 vccd1 vccd1 _5810_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8952__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6790_ _6511_/A _6789_/X _5824_/X _6908_/B vssd1 vssd1 vccd1 vccd1 _6790_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5741_ _5741_/A _5741_/B vssd1 vssd1 vccd1 vccd1 _5741_/X sky130_fd_sc_hd__and2_1
XANTENNA__4955__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8460_ _8460_/A _8482_/B vssd1 vssd1 vccd1 vccd1 _8460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5672_ _5672_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _5672_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_127_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7354__B1 _7349_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8697__A3 hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7411_ _7630_/B vssd1 vssd1 vccd1 vccd1 _7668_/B sky130_fd_sc_hd__buf_6
XFILLER_0_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4623_ _7398_/A hold7/X vssd1 vssd1 vccd1 vccd1 _8926_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8391_ _8390_/Y _8369_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8392_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7342_ _7340_/Y _7332_/A _7341_/Y vssd1 vssd1 vccd1 vccd1 _7342_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4554_ _4554_/A hold29/X vssd1 vssd1 vccd1 vccd1 _4839_/B sky130_fd_sc_hd__and2_1
XANTENNA__6510__A _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7106__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5380__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7273_ _6342_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7273_/X sky130_fd_sc_hd__a21o_1
X_4485_ _4485_/A _4485_/B vssd1 vssd1 vccd1 vccd1 _8240_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_111_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6224_ _6223_/X _6941_/B _6224_/S vssd1 vssd1 vccd1 vccd1 _6225_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_40_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5132__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6155_ _6593_/A _6118_/A _6154_/Y vssd1 vssd1 vccd1 vccd1 _6156_/A sky130_fd_sc_hd__o21ai_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6880__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7341__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5106_/A _5106_/B vssd1 vssd1 vccd1 vccd1 _5106_/Y sky130_fd_sc_hd__nor2_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6089_/A1 _5192_/X input60/X _5193_/X vssd1 vssd1 vccd1 vccd1 _6086_/X sky130_fd_sc_hd__o22a_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5037_ input85/X _8716_/B input22/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5840__B1 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8385__A2 _8352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6396__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5199__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8172__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6396__B2 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6988_ _6988_/A vssd1 vssd1 vccd1 vccd1 _6988_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__7593__B1 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8790__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8727_ _8320_/X _8806_/B _8721_/X _8726_/X vssd1 vssd1 vccd1 vccd1 _8727_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5939_ _5936_/Y _4890_/A _5937_/Y _4885_/A _5938_/Y vssd1 vssd1 vccd1 vccd1 _6839_/B
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6404__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8137__A2 _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6148__A1 _6183_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6148__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8658_ _8464_/A _8581_/X _8469_/A _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8658_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7609_ _7378_/X _5924_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7609_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8589_ _8589_/A vssd1 vssd1 vccd1 vccd1 _8698_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5036__A _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput100 mports_i[18] vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__buf_4
Xinput111 mports_i[19] vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__clkbuf_4
Xinput122 mports_i[209] vssd1 vssd1 vccd1 vccd1 _6061_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__7251__A _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput133 mports_i[219] vssd1 vssd1 vccd1 vccd1 _6286_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__8073__A1 _8080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput144 mports_i[23] vssd1 vssd1 vccd1 vccd1 _5591_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8073__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput155 mports_i[33] vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__clkbuf_4
Xinput166 mports_i[43] vssd1 vssd1 vccd1 vccd1 _6158_/A sky130_fd_sc_hd__buf_2
Xinput177 mports_i[53] vssd1 vssd1 vccd1 vccd1 _6358_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7820__A1 _7827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput188 mports_i[63] vssd1 vssd1 vccd1 vccd1 _5131_/B2 sky130_fd_sc_hd__buf_2
XANTENNA__7820__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput199 mports_i[73] vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6387__A1 _6387_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6387__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8781__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6314__B _6314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8128__A2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7887__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output479_A _7895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4769__B _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput607 _5680_/X vssd1 vssd1 vccd1 vccd1 sports_o[195] sky130_fd_sc_hd__buf_12
Xoutput618 _5920_/X vssd1 vssd1 vccd1 vccd1 sports_o[204] sky130_fd_sc_hd__buf_12
Xoutput629 _6220_/X vssd1 vssd1 vccd1 vccd1 sports_o[214] sky130_fd_sc_hd__buf_12
XANTENNA__8836__B1 _8240_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5114__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6311__B2 _6310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6862__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7393__A1_N _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8064__A1 _8067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8064__B2 _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7811__A1 _7814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6614__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7960_ _7777_/X _8765_/B _7792_/X vssd1 vssd1 vccd1 vccd1 _7960_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__7811__B2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6911_ _6911_/A _6933_/A vssd1 vssd1 vccd1 vccd1 _6911_/Y sky130_fd_sc_hd__nand2_1
X_7891_ _7888_/Y _7768_/X _7890_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7891_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6842_ _5915_/Y _6912_/B _6838_/X _6840_/Y _6841_/Y vssd1 vssd1 vccd1 vccd1 _6843_/A
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6505__A _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6378__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6773_ _6506_/A _6770_/A _6449_/A vssd1 vssd1 vccd1 vccd1 _6773_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_92_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8119__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5724_ _5274_/A _5792_/A1 _5275_/A input49/X vssd1 vssd1 vccd1 vccd1 _5724_/Y sky130_fd_sc_hd__a22oi_1
X_8512_ _8510_/Y _8511_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8540_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8443_ _8042_/Y _8518_/B _8572_/S vssd1 vssd1 vccd1 vccd1 _8443_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7878__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5655_ _5655_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _7529_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_115_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606_ _5229_/A vssd1 vssd1 vccd1 vccd1 _6102_/B sky130_fd_sc_hd__inv_4
XFILLER_0_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8374_ _8374_/A vssd1 vssd1 vccd1 vccd1 _8374_/X sky130_fd_sc_hd__buf_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5586_ _5585_/X _5562_/X _6356_/S vssd1 vssd1 vccd1 vccd1 _5586_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7325_ _7334_/A vssd1 vssd1 vccd1 vccd1 _7326_/A sky130_fd_sc_hd__buf_8
XANTENNA__7055__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8827__B1 _8219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4537_ hold29/X _8716_/A vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7256_ _7256_/A vssd1 vssd1 vccd1 vccd1 _7256_/X sky130_fd_sc_hd__buf_1
X_4468_ _5185_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4468_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6302__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6207_ _6207_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6207_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6386__S _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7187_ _7187_/A vssd1 vssd1 vccd1 vccd1 _7187_/X sky130_fd_sc_hd__buf_1
X_4399_ _4458_/A _4658_/A _4458_/B vssd1 vssd1 vccd1 vccd1 _4454_/B sky130_fd_sc_hd__nand3_1
X_6138_ _6174_/A1 _4935_/A input64/X _4939_/A vssd1 vssd1 vccd1 vccd1 _6138_/X sky130_fd_sc_hd__o22a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8055__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7802__A1 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6605__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6069_ _6075_/A _4953_/X _6076_/A _4870_/A _6068_/X vssd1 vssd1 vccd1 vccd1 _6913_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__7802__B2 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6369__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7869__B2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8530__A2 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6541__A1 _7383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4589__B _7309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6541__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6844__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8597__A2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5213__B _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7021__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5032__A1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6044__B _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5032__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8521__A2 _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5440_ _5440_/A vssd1 vssd1 vccd1 vccd1 _5440_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6532__A1 _7356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6532__B2 _5159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput404 _8837_/X vssd1 vssd1 vccd1 vccd1 mports_o[134] sky130_fd_sc_hd__buf_12
X_5371_ _5367_/Y _5370_/Y _8842_/B vssd1 vssd1 vccd1 vccd1 _5372_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput415 _8083_/X vssd1 vssd1 vccd1 vccd1 mports_o[21] sky130_fd_sc_hd__buf_12
Xoutput426 _8237_/X vssd1 vssd1 vccd1 vccd1 mports_o[31] sky130_fd_sc_hd__buf_12
Xoutput437 _8329_/X vssd1 vssd1 vccd1 vccd1 mports_o[41] sky130_fd_sc_hd__buf_12
XFILLER_0_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7110_ _7110_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7110_/X sky130_fd_sc_hd__and2_1
XANTENNA__8285__A1 _7809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput448 _8438_/X vssd1 vssd1 vccd1 vccd1 mports_o[51] sky130_fd_sc_hd__buf_12
X_4322_ _4322_/A _7847_/A vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__nand2_1
X_8090_ _8093_/A1 _5780_/X _8093_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _8090_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__8285__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput459 _8534_/X vssd1 vssd1 vccd1 vccd1 mports_o[61] sky130_fd_sc_hd__buf_12
XANTENNA__5099__A1 _6489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6296__B1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7041_ _7040_/Y _7341_/B _7097_/S vssd1 vssd1 vccd1 vccd1 _7042_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8037__A1 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8037__B2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8588__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6599__A1 _5328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7796__B1 _7803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6599__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7943_ _8351_/A _7768_/X _7942_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7943_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7874_ _7874_/A vssd1 vssd1 vccd1 vccd1 _7874_/X sky130_fd_sc_hd__buf_12
XANTENNA__7548__B1 _7359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8745__C1 _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6825_ _5930_/Y _6475_/A _5877_/X _6694_/B vssd1 vssd1 vccd1 vccd1 _6825_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5023__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6756_ _6852_/A _6756_/B vssd1 vssd1 vccd1 vccd1 _6756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6889__B _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ _5707_/A vssd1 vssd1 vccd1 vccd1 _5707_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6687_ _5500_/X _6913_/B _5502_/X _6912_/B vssd1 vssd1 vccd1 vccd1 _6687_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5285__S _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8426_ _8426_/A vssd1 vssd1 vccd1 vccd1 _8426_/Y sky130_fd_sc_hd__inv_2
X_5638_ _5596_/A _4929_/A _5597_/A _4932_/A _5637_/X vssd1 vssd1 vccd1 vccd1 _5655_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5326__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6523__A1 _5161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6523__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8357_ _8376_/A _8323_/X _8355_/X _8356_/X vssd1 vssd1 vccd1 vccd1 _8357_/X sky130_fd_sc_hd__a22o_2
X_5569_ _6212_/A _5558_/X _5108_/A _5568_/Y _5136_/X vssd1 vssd1 vccd1 vccd1 _5569_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7308_ _4876_/X _7753_/B _4899_/Y _7349_/A vssd1 vssd1 vccd1 vccd1 _7308_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8276__A1 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7079__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8276__B2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8288_ _8288_/A vssd1 vssd1 vccd1 vccd1 _8288_/X sky130_fd_sc_hd__buf_1
XANTENNA__6287__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6826__A2 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7239_ _7238_/X _7705_/B _7249_/S vssd1 vssd1 vccd1 vccd1 _7240_/A sky130_fd_sc_hd__mux2_2
XANTENNA__7787__B1 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8200__A1 _8210_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7003__A2 _4408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8200__B2 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5014__A1 _5011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8751__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5565__A2 _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8967__RESET_B input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8519__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8019__A1 _8024_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7490__A2 _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output511_A _6979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5253__A1 _5218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5253__B2 _6578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4940_ _4940_/A vssd1 vssd1 vccd1 vccd1 _4940_/X sky130_fd_sc_hd__buf_8
XFILLER_0_86_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4871_ _4871_/A vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__buf_6
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5005__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5005__B2 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8742__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6610_ _6801_/A _5317_/A _6450_/A vssd1 vssd1 vccd1 vccd1 _6610_/X sky130_fd_sc_hd__o21a_1
XANTENNA__8270__A _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7590_ _7590_/A _7590_/B vssd1 vssd1 vccd1 vccd1 _7590_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5556__A2 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7950__B1 _7958_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6541_ _7383_/A _6475_/X _6540_/X _6851_/B vssd1 vssd1 vccd1 vccd1 _6542_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6472_ _6470_/Y _6471_/Y _6780_/A vssd1 vssd1 vccd1 vccd1 _6472_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4303__A _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8211_ _8211_/A vssd1 vssd1 vccd1 vccd1 _8211_/Y sky130_fd_sc_hd__inv_2
X_5423_ _5466_/A _6875_/B _5422_/X vssd1 vssd1 vccd1 vccd1 _5423_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_152_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5354_ _6870_/S _5245_/X _5353_/Y vssd1 vssd1 vccd1 vccd1 _6621_/A sky130_fd_sc_hd__o21ai_2
X_8142_ _8142_/A vssd1 vssd1 vccd1 vccd1 _8143_/B sky130_fd_sc_hd__inv_2
XFILLER_0_140_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6269__B1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4305_ _5827_/B _4591_/B _4719_/B vssd1 vssd1 vccd1 vccd1 _4305_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8073_ _8080_/A1 _4947_/B _8080_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _8073_/Y sky130_fd_sc_hd__o22ai_2
X_5285_ _5343_/B _5283_/Y _6711_/S vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5134__A _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7024_ _7023_/X _4963_/X _7295_/S vssd1 vssd1 vccd1 vccd1 _7024_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__7481__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5492__A1 _5440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5492__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8445__A _8445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7233__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8975_ _8976_/CLK _8975_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__5244__A1 _5272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5244__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7926_ _7931_/A1 _5145_/A _7931_/B1 _5616_/A vssd1 vssd1 vccd1 vccd1 _7926_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_0_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8718__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7857_ _7851_/Y _7768_/X _7772_/X _7856_/Y _7774_/X vssd1 vssd1 vccd1 vccd1 _7857_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8180__A _8180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6808_ _6807_/Y _5832_/Y _6851_/B vssd1 vssd1 vccd1 vccd1 _6808_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5547__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7941__B1 _7944_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7788_ _7790_/B2 _7299_/A _7790_/A2 _7769_/A _7787_/X vssd1 vssd1 vccd1 vccd1 _7788_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_147_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6739_ _5738_/C _6549_/A _5684_/X _6876_/C vssd1 vssd1 vccd1 vccd1 _6739_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6412__B _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8409_ _8424_/A _8299_/X _8408_/Y _8304_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8409_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7524__A _7524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5180__B1 _5222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8249__A1 _8251_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8249__B2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5979__A _6028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5483__A1 _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4883__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8421__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__A1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6983__A1 _7737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__B1 _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7418__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5219__A _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8488__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7160__A1 _5744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7153__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _5070_/A vssd1 vssd1 vccd1 vccd1 _5070_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8660__A1 _8491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5474__A1 _5697_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5474__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4793__A _4793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8265__A _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7215__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5226__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5226__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8760_ _7942_/Y _8711_/A _8408_/Y _8770_/B vssd1 vssd1 vccd1 vccd1 _8760_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6974__A1 _7729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5972_ _7630_/A _8160_/A _6456_/B _7622_/A vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_149_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7711_ _7711_/A vssd1 vssd1 vccd1 vccd1 _7711_/X sky130_fd_sc_hd__buf_1
X_4923_ _6211_/B vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__inv_2
X_8691_ _8691_/A vssd1 vssd1 vccd1 vccd1 _8691_/X sky130_fd_sc_hd__buf_1
XFILLER_0_87_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8176__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6513__A _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7642_ _6063_/A _7389_/A _6893_/Y _7361_/X vssd1 vssd1 vccd1 vccd1 _7642_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5529__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4854_ _4858_/A _8933_/A vssd1 vssd1 vccd1 vccd1 _4863_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6726__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4785_ _4785_/A _4813_/C vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7573_ _7573_/A vssd1 vssd1 vccd1 vccd1 _7573_/X sky130_fd_sc_hd__buf_1
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6524_ _6899_/B vssd1 vssd1 vccd1 vccd1 _6933_/A sky130_fd_sc_hd__buf_6
XFILLER_0_126_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6455_ _6481_/A _6875_/B _6454_/X vssd1 vssd1 vccd1 vccd1 _6455_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7151__A1 _6743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5406_ _5405_/Y _5389_/Y _7847_/A vssd1 vssd1 vccd1 vccd1 _7450_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6386_ _6382_/X _6385_/Y _6386_/S vssd1 vssd1 vccd1 vccd1 _6386_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5701__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5337_ _5337_/A vssd1 vssd1 vccd1 vccd1 _5337_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8125_ _8132_/A1 _4947_/B _8132_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _8125_/Y sky130_fd_sc_hd__o22ai_2
X_5268_ _5265_/Y _4891_/A _5266_/Y _4886_/A _5267_/Y vssd1 vssd1 vccd1 vccd1 _6576_/B
+ sky130_fd_sc_hd__o221a_4
X_8056_ _7777_/X _8055_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _8056_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__8651__A1 _8036_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7454__A2 _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8651__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5799__A _6771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7007_ _7272_/A _7272_/C vssd1 vssd1 vccd1 vccd1 _7008_/A sky130_fd_sc_hd__and2_1
X_5199_ _5105_/A _5197_/X _8151_/B _5196_/A vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_98_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7206__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6407__B _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5217__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5217__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8958_ _8978_/CLK _8958_/D fanout732/X vssd1 vssd1 vccd1 vccd1 _8958_/Q sky130_fd_sc_hd__dfrtp_4
X_7909_ _7909_/A vssd1 vssd1 vccd1 vccd1 _7909_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8889_ _8886_/Y _8888_/Y _8880_/Y vssd1 vssd1 vccd1 vccd1 _8892_/A sky130_fd_sc_hd__a21o_1
XANTENNA__8167__B1 _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6423__A _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6717__B2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7390__B2 _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4878__A _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7142__A1 _5679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8890__A1 _4661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7693__A2 _7359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8642__A1 _8400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5456__A1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5456__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5208__A1 _5208_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5208__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7602__C1 _7347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6956__A1 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7905__B1 _7905_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7148__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4570_ _4658_/A _8181_/A _7707_/C vssd1 vssd1 vccd1 vccd1 _4570_/X sky130_fd_sc_hd__or3_1
XANTENNA__5392__B1 _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5891__B _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8330__B1 _7903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6240_ _6247_/A1 _8310_/B input68/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6240_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7684__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5695__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6171_ _6182_/A1 _5192_/A input65/X _5193_/A vssd1 vssd1 vccd1 vccd1 _6171_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5122_ _7352_/B vssd1 vssd1 vccd1 vccd1 _5123_/B sky130_fd_sc_hd__inv_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8633__A1 _8404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8633__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5447__A1 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5447__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5053_ _8755_/C vssd1 vssd1 vccd1 vccd1 _7629_/B sky130_fd_sc_hd__buf_8
XANTENNA__7611__B _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5412__A _5412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7103__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8812_ _8145_/Y _8803_/B _8148_/X _8711_/X _8788_/S vssd1 vssd1 vccd1 vccd1 _8812_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4958__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8743_ _8833_/B _7878_/Y _8725_/A vssd1 vssd1 vccd1 vccd1 _8743_/X sky130_fd_sc_hd__o21a_1
X_5955_ _5159_/B _5899_/A _5125_/X _7610_/A _5954_/X vssd1 vssd1 vccd1 vccd1 _5955_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8149__B1 _8148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4906_ _4906_/A vssd1 vssd1 vccd1 vccd1 _6367_/A sky130_fd_sc_hd__inv_2
XFILLER_0_36_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8674_ _8550_/A _8580_/A _8130_/Y _8583_/A vssd1 vssd1 vccd1 vccd1 _8674_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5886_ _5928_/A1 _4934_/A input54/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5886_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5347__A2_N _7422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7625_ _6861_/A _7696_/B _7618_/Y _7700_/B vssd1 vssd1 vccd1 vccd1 _7625_/X sky130_fd_sc_hd__a22o_1
X_4837_ _4837_/A _7511_/B vssd1 vssd1 vccd1 vccd1 _8904_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6175__A2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7556_ _7590_/A _7556_/B vssd1 vssd1 vccd1 vccd1 _7556_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4768_ _4768_/A _4768_/B vssd1 vssd1 vccd1 vccd1 _4792_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6507_ _6801_/A _6507_/B vssd1 vssd1 vccd1 vccd1 _6507_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7124__A1 _5530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4698__A _5130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7487_ _5549_/Y _7668_/B _5580_/X _7638_/B _7753_/B vssd1 vssd1 vccd1 vccd1 _7487_/X
+ sky130_fd_sc_hd__a221o_1
X_4699_ _4699_/A _7272_/B vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6438_ _6462_/A vssd1 vssd1 vccd1 vccd1 _6841_/A sky130_fd_sc_hd__buf_8
XANTENNA__7675__A2 _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6883__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6369_ _6369_/A1 _8480_/B input14/X _4870_/X _6368_/X vssd1 vssd1 vccd1 vccd1 _7743_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8108_ _7777_/A _8107_/Y _7792_/A vssd1 vssd1 vccd1 vccd1 _8108_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__8624__A1 _7929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput304 sports_i[44] vssd1 vssd1 vccd1 vccd1 _7923_/A sky130_fd_sc_hd__buf_1
XANTENNA__8624__B2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput315 sports_i[54] vssd1 vssd1 vccd1 vccd1 _8059_/A sky130_fd_sc_hd__clkbuf_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput326 sports_i[64] vssd1 vssd1 vccd1 vccd1 _4478_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5438__B2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__buf_1
Xinput337 sports_i[74] vssd1 vssd1 vccd1 vccd1 _7877_/B1 sky130_fd_sc_hd__clkbuf_4
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
X_8039_ _8039_/A vssd1 vssd1 vccd1 vccd1 _8468_/A sky130_fd_sc_hd__inv_2
Xinput348 sports_i[84] vssd1 vssd1 vccd1 vccd1 _8011_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__6418__A _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput359 sports_i[94] vssd1 vssd1 vccd1 vccd1 _8150_/B sky130_fd_sc_hd__buf_2
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6938__A1 _6221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6938__B2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8352__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5992__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8560__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_8 _7174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4401__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6323__C1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8615__A1 _7886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5429__A1 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5429__B2 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7431__B _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output424_A _7805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8091__A2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6929__A1 _7683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6063__A _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5740_ _6128_/B _7544_/A _5136_/A vssd1 vssd1 vccd1 vccd1 _5740_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7354__A1 _5150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5671_ _6837_/A _5668_/X _5670_/X vssd1 vssd1 vccd1 vccd1 _6724_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7354__B2 _6514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7410_ _5330_/Y _7619_/B _7406_/X _7408_/Y _7409_/Y vssd1 vssd1 vccd1 vccd1 _7410_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__5365__B1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4622_ _4943_/A vssd1 vssd1 vccd1 vccd1 _7398_/A sky130_fd_sc_hd__buf_8
XFILLER_0_114_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8390_ _8390_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7341_ _7756_/A _7341_/B vssd1 vssd1 vccd1 vccd1 _7341_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4553_ _4837_/A _4553_/B vssd1 vssd1 vccd1 vccd1 _4612_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_53_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7106__A1 _6648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8303__B1 _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4311__A _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8854__A1 _7372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4484_ _4476_/X _4484_/B _8189_/B vssd1 vssd1 vccd1 vccd1 _4485_/B sky130_fd_sc_hd__nand3b_1
X_7272_ _7272_/A _7272_/B _7272_/C vssd1 vssd1 vccd1 vccd1 _7272_/X sky130_fd_sc_hd__and3_1
XANTENNA__5668__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6223_ _6222_/X _7696_/A _6356_/S vssd1 vssd1 vccd1 vccd1 _6223_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6154_ _6154_/A _6593_/A vssd1 vssd1 vccd1 vccd1 _6154_/Y sky130_fd_sc_hd__nand2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8606__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7341__B _7341_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A vssd1 vssd1 vccd1 vccd1 _5106_/B sky130_fd_sc_hd__inv_2
X_6085_ _5096_/A _6912_/A _6083_/X _5715_/B _6084_/X vssd1 vssd1 vccd1 vccd1 _6085_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8082__A2 _8081_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6093__A1 _6104_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6093__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5036_ _7311_/A vssd1 vssd1 vccd1 vccd1 _7536_/B sky130_fd_sc_hd__clkbuf_16
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5840__A1 _5827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5840__B2 _5803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5796__B _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8172__B _8172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6987_ _6986_/X _6358_/X _7001_/S vssd1 vssd1 vccd1 vccd1 _6988_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7593__A1 _7532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8790__B1 _8469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8726_ _8833_/B _8317_/X _8725_/X vssd1 vssd1 vccd1 vccd1 _8726_/X sky130_fd_sc_hd__o21a_1
X_5938_ _5274_/A _5962_/A1 _5275_/A input55/X vssd1 vssd1 vccd1 vccd1 _5938_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_137_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8657_ _8657_/A vssd1 vssd1 vccd1 vccd1 _8657_/X sky130_fd_sc_hd__buf_1
X_5869_ _5866_/Y _4886_/A _5867_/Y _4891_/A _5868_/Y vssd1 vssd1 vccd1 vccd1 _5930_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6148__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7608_ _7683_/B _7606_/B _7605_/X _7606_/X _7607_/Y vssd1 vssd1 vccd1 vccd1 _7608_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6701__A _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8588_ _7765_/X _8581_/X _7771_/X _8583_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8588_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7539_ _6733_/A _7696_/B _7537_/X _7538_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7539_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6420__B _6528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5317__A _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7532__A _7532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput101 mports_i[190] vssd1 vssd1 vccd1 vccd1 _5497_/A1 sky130_fd_sc_hd__buf_2
Xinput112 mports_i[1] vssd1 vssd1 vccd1 vccd1 _4956_/A sky130_fd_sc_hd__buf_2
XANTENNA__6608__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput123 mports_i[20] vssd1 vssd1 vccd1 vccd1 _5510_/A sky130_fd_sc_hd__clkbuf_4
Xinput134 mports_i[21] vssd1 vssd1 vccd1 vccd1 _5505_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8073__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput145 mports_i[24] vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__clkbuf_4
Xinput156 mports_i[34] vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__clkbuf_4
Xinput167 mports_i[44] vssd1 vssd1 vccd1 vccd1 _6183_/A1 sky130_fd_sc_hd__buf_2
Xinput178 mports_i[54] vssd1 vssd1 vccd1 vccd1 _6369_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput189 mports_i[64] vssd1 vssd1 vccd1 vccd1 _5140_/A sky130_fd_sc_hd__buf_2
XANTENNA__7820__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5831__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4891__A _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7033__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6387__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8533__B1 _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7707__A _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6611__A _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput608 _5706_/X vssd1 vssd1 vccd1 vccd1 sports_o[196] sky130_fd_sc_hd__buf_12
XANTENNA__8836__A1 _8239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput619 _5955_/X vssd1 vssd1 vccd1 vccd1 sports_o[205] sky130_fd_sc_hd__buf_12
XANTENNA__8836__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output639_A _6347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8257__B _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8064__A2 _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6058__A _6058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7811__A2 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5822__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6910_ _7668_/A _6475_/X _6082_/X _6851_/B vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__a22o_1
X_7890_ _7884_/Y _6500_/X _7883_/Y _7769_/X _7889_/X vssd1 vssd1 vccd1 vccd1 _7890_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6841_ _6841_/A _6841_/B vssd1 vssd1 vccd1 vccd1 _6841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6378__A2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5586__A0 _5585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4306__A hold4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6772_ _8150_/A _6770_/Y _7558_/A vssd1 vssd1 vccd1 vccd1 _6772_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8511_ _8511_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5723_ _5723_/A vssd1 vssd1 vccd1 vccd1 _5723_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7327__B2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8442_ _8555_/B _8440_/X _8441_/Y vssd1 vssd1 vccd1 vccd1 _8442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7878__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5654_ _6743_/A vssd1 vssd1 vccd1 vccd1 _5654_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4605_ _4605_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4610_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8373_ _8367_/X _8372_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8374_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5585_ _5096_/A _5574_/X _5582_/X _5715_/B _5584_/Y vssd1 vssd1 vccd1 vccd1 _5585_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8827__A1 _8217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7324_ _7715_/S vssd1 vssd1 vccd1 vccd1 _7334_/A sky130_fd_sc_hd__inv_2
XFILLER_0_130_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4536_ _8584_/B vssd1 vssd1 vccd1 vccd1 _8716_/A sky130_fd_sc_hd__inv_6
XFILLER_0_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6838__B1 _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7255_ _7254_/Y _7720_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7256_/A sky130_fd_sc_hd__mux2_2
XANTENNA__4976__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6667__S _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6302__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4467_ _4482_/A vssd1 vssd1 vccd1 vccd1 _5185_/A sky130_fd_sc_hd__buf_8
XFILLER_0_68_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7352__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6206_ _6227_/A _8335_/B input4/X _4913_/A _6205_/X vssd1 vssd1 vccd1 vccd1 _6207_/A
+ sky130_fd_sc_hd__o221a_4
X_7186_ _7185_/X _5885_/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7187_/A sky130_fd_sc_hd__mux2_4
X_4398_ _4398_/A hold40/A vssd1 vssd1 vccd1 vccd1 _4458_/B sky130_fd_sc_hd__nand2_1
XANTENNA__7071__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6137_ _6075_/A _4929_/A _6076_/A _4932_/A _6136_/X vssd1 vssd1 vccd1 vccd1 _6908_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8055__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7802__A2 _7802_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6068_ _6136_/A1 _5090_/A input62/X _4874_/A vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5019_ _5019_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _5060_/B sky130_fd_sc_hd__nand2_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5600__A _5666_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6369__A2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5577__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8709_ _8709_/A _8709_/B vssd1 vssd1 vccd1 vccd1 _8712_/A sky130_fd_sc_hd__nor2_2
XANTENNA__7318__A1 _4942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6431__A _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7869__A2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7246__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6541__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8818__A1 _8157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4886__A _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8358__A _8358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5501__B1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__A1 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__B2 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5213__C _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5510__A _5510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8821__A _8821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5032__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output589_A _5203_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6532__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput405 _8840_/X vssd1 vssd1 vccd1 vccd1 mports_o[135] sky130_fd_sc_hd__buf_12
X_5370_ _6611_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5370_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5740__B1 _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput416 _8096_/X vssd1 vssd1 vccd1 vccd1 mports_o[22] sky130_fd_sc_hd__buf_12
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput427 _8242_/X vssd1 vssd1 vccd1 vccd1 mports_o[32] sky130_fd_sc_hd__buf_12
Xoutput438 _8332_/X vssd1 vssd1 vccd1 vccd1 mports_o[42] sky130_fd_sc_hd__buf_12
X_4321_ _4321_/A _4321_/B vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8285__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8268__A _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput449 _8450_/X vssd1 vssd1 vccd1 vccd1 mports_o[52] sky130_fd_sc_hd__buf_12
XANTENNA__6296__A1 _6309_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5099__A2 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6296__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7040_ _7040_/A vssd1 vssd1 vccd1 vccd1 _7040_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7796__A1 _4566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6599__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7796__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7942_ _7935_/Y _7769_/X _7936_/Y _6500_/X _7941_/Y vssd1 vssd1 vccd1 vccd1 _7942_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7873_ _7869_/Y _7768_/X _7871_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7873_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8745__B1 _7890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5559__B1 _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6824_ _5860_/A _6913_/B _5864_/Y _6912_/B vssd1 vssd1 vccd1 vccd1 _6824_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_147_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6755_ _6755_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6755_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_135_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7347__A _7347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5706_ _5031_/X _5655_/A _5696_/X _5705_/X vssd1 vssd1 vccd1 vccd1 _5706_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6686_ _6724_/A _5517_/Y _5549_/Y _6475_/X vssd1 vssd1 vccd1 vccd1 _6686_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8425_ _8423_/Y _8424_/Y _8481_/S vssd1 vssd1 vccd1 vccd1 _8426_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_104_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5637_ _5637_/A1 _4935_/A input44/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5637_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6523__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8965__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8356_ _8564_/B _7945_/Y _8349_/A vssd1 vssd1 vccd1 vccd1 _8356_/X sky130_fd_sc_hd__o21a_1
X_5568_ _5568_/A vssd1 vssd1 vccd1 vccd1 _5568_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7307_ _7347_/A _7678_/A vssd1 vssd1 vccd1 vccd1 _7349_/A sky130_fd_sc_hd__nor2_8
X_4519_ _8240_/A _4436_/A _4518_/Y _4517_/B vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__a31o_1
X_8287_ _8286_/X _7807_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8288_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8178__A _8192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5499_ _5557_/A1 _5090_/A input40/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5499_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6287__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8681__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7238_ _6207_/A _7026_/X _7237_/X vssd1 vssd1 vccd1 vccd1 _7238_/X sky130_fd_sc_hd__o21a_1
X_7169_ _7168_/X _5772_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7170_/A sky130_fd_sc_hd__mux2_2
XANTENNA__6039__A1 _6047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6039__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7787__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7787__B2 _7791_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8736__B1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8200__A2 _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6161__A _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5505__A _5505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8019__A2 _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7720__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8535__B _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5240__A _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5253__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4461__A0 _8180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ _4870_/A vssd1 vssd1 vccd1 vccd1 _4870_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5005__A2 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7950__A1 _7958_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6753__A2 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7167__A _7167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6540_ _6539_/X _5146_/Y _6837_/A vssd1 vssd1 vccd1 vccd1 _6540_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6471_ _6231_/C _4899_/A _7829_/A vssd1 vssd1 vccd1 vccd1 _6471_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8210_ _8210_/A1 _6102_/B _8210_/B1 _5106_/A _8209_/X vssd1 vssd1 vccd1 vccd1 _8211_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_42_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5422_ _6634_/A _8188_/S hold23/A vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8141_ _8141_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _8141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5353_ _5353_/A _6870_/S vssd1 vssd1 vccd1 vccd1 _5353_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6269__A1 _6286_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6269__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4304_ hold45/X vssd1 vssd1 vccd1 vccd1 _4719_/B sky130_fd_sc_hd__inv_2
X_8072_ _8072_/A vssd1 vssd1 vccd1 vccd1 _8072_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5284_ _6166_/B vssd1 vssd1 vccd1 vccd1 _6711_/S sky130_fd_sc_hd__inv_4
X_7023_ _7138_/A vssd1 vssd1 vccd1 vccd1 _7023_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5492__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4973__B _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8974_ _8976_/CLK _8974_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__5150__A _5150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5244__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7925_ _7922_/Y _7013_/A _7923_/Y _5116_/A _7924_/Y vssd1 vssd1 vccd1 vccd1 _8345_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__8718__B1 _8303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7856_ _7856_/A vssd1 vssd1 vccd1 vccd1 _7856_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6807_ _6837_/A _6807_/B vssd1 vssd1 vccd1 vccd1 _6807_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7787_ _5185_/A _7791_/B1 _6500_/A _7791_/A1 vssd1 vssd1 vccd1 vccd1 _7787_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_81_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4999_ input83/X _8716_/B input20/X _4917_/X vssd1 vssd1 vccd1 vccd1 _4999_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7941__A1 _7944_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7941__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4755__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6738_ _7153_/A _6475_/A _5693_/X _6694_/B vssd1 vssd1 vccd1 vccd1 _6738_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6669_ _6852_/A _6669_/B vssd1 vssd1 vccd1 vccd1 _6669_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8408_ _8300_/B _8354_/A _8407_/Y vssd1 vssd1 vccd1 vccd1 _8408_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7524__B _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5180__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8339_ _8567_/B _8337_/Y _8338_/X vssd1 vssd1 vccd1 vccd1 _8339_/X sky130_fd_sc_hd__o21a_1
XANTENNA__8249__A2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5180__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5979__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8421__A2 _8012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5060__A _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4994__A1 _4978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7932__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8488__A2 _8081_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output454_A _8509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7448__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7999__B2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6120__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8660__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output719_A _6822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7450__A _7450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5474__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5226__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5971_ _5971_/A vssd1 vssd1 vccd1 vccd1 _7622_/A sky130_fd_sc_hd__inv_2
X_7710_ _7709_/X _6248_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7711_/A sky130_fd_sc_hd__mux2_1
X_4922_ _8716_/A _7876_/A vssd1 vssd1 vccd1 vccd1 _6211_/B sky130_fd_sc_hd__nor2_4
X_8690_ _8689_/X _8200_/X _8690_/S vssd1 vssd1 vccd1 vccd1 _8691_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8176__A1 _8175_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7641_ _7542_/A _6016_/A _7326_/A vssd1 vssd1 vccd1 vccd1 _7641_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_129_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4853_ _8977_/D _8976_/D vssd1 vssd1 vccd1 vccd1 _8933_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6187__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7572_ _7571_/X _5772_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7573_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4784_ _4784_/A _4786_/B vssd1 vssd1 vccd1 vccd1 _4813_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6523_ _5161_/X _6475_/X _5163_/X _6851_/B vssd1 vssd1 vccd1 vccd1 _6525_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6454_ _4876_/X _8188_/S _6544_/B _6593_/A vssd1 vssd1 vccd1 vccd1 _6454_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_113_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5405_ _6079_/A _6646_/B vssd1 vssd1 vccd1 vccd1 _5405_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6385_ _6385_/A vssd1 vssd1 vccd1 vccd1 _6385_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5145__A _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8124_ _8124_/A vssd1 vssd1 vccd1 vccd1 _8124_/Y sky130_fd_sc_hd__inv_2
X_5336_ _7432_/B vssd1 vssd1 vccd1 vccd1 _5336_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8100__B2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8055_ _8045_/Y _7874_/X _8046_/Y _7875_/X _8054_/Y vssd1 vssd1 vccd1 vccd1 _8055_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__4984__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5267_ _4893_/A input92/X _4896_/A input29/X vssd1 vssd1 vccd1 vccd1 _5267_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__8651__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7360__A _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7006_ _6080_/A _8755_/C hold40/A _4408_/B vssd1 vssd1 vccd1 vccd1 _7272_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5198_ _8181_/A vssd1 vssd1 vccd1 vccd1 _8151_/B sky130_fd_sc_hd__buf_6
X_8957_ _8976_/CLK hold17/X fanout733/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7908_ _7760_/X _8346_/A _7904_/X _7907_/X vssd1 vssd1 vccd1 vccd1 _7908_/X sky130_fd_sc_hd__a22o_2
X_8888_ _8888_/A vssd1 vssd1 vccd1 vccd1 _8888_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8167__A1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7839_ _7760_/X _7821_/Y _7833_/X _7838_/Y vssd1 vssd1 vccd1 vccd1 _7839_/X sky130_fd_sc_hd__a22o_2
XANTENNA__6423__B _7372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7914__B2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7390__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6350__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4894__A _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5456__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5208__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7602__B1 _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4967__A1 _4966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6169__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7905__A1 _7905_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6708__A2 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7905__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5392__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8951__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7669__B1 _7385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8330__A1 _7901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8330__B2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5695__A2 _7524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6170_ _6170_/A _6170_/B vssd1 vssd1 vccd1 vccd1 _6170_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5121_ _5131_/A2 _4929_/A _5131_/B2 _4932_/A _5120_/X vssd1 vssd1 vccd1 vccd1 _7352_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__8633__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7180__A _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5447__A2 _7105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5052_ hold39/A vssd1 vssd1 vccd1 vccd1 _8755_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5412__B _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8397__A1 _7983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8397__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8811_ _8811_/A vssd1 vssd1 vccd1 vccd1 _8811_/X sky130_fd_sc_hd__buf_1
XFILLER_0_95_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4958__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8742_ _7869_/Y _8803_/B _7871_/Y _8711_/X _8820_/B vssd1 vssd1 vccd1 vccd1 _8742_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4958__B2 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5954_ _6128_/B _6827_/A _5136_/A _5953_/X vssd1 vssd1 vccd1 vccd1 _5954_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6524__A _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8149__A1 _8145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8149__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _5055_/A _5672_/A vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8673_ _8519_/A _8686_/B _8671_/X _8672_/X vssd1 vssd1 vccd1 vccd1 _8673_/X sky130_fd_sc_hd__a22o_1
X_5885_ _5871_/A _5111_/A _5872_/A _4931_/A _5884_/X vssd1 vssd1 vccd1 vccd1 _5885_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7624_ _6002_/Y _7660_/B _7621_/X _7622_/Y _7623_/Y vssd1 vssd1 vccd1 vccd1 _7624_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_7_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4836_ hold10/X _8919_/A _4833_/Y _4835_/X vssd1 vssd1 vccd1 vccd1 _8976_/D sky130_fd_sc_hd__a31o_2
XFILLER_0_145_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7555_ _7556_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7555_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4767_ _4767_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _4768_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5574__S _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6506_ _6506_/A vssd1 vssd1 vccd1 vccd1 _6801_/A sky130_fd_sc_hd__buf_8
X_7486_ _7486_/A vssd1 vssd1 vccd1 vccd1 _7486_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8321__A1 _8320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4698_ _5130_/A _4719_/B vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5135__A1 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6437_ _6724_/A _4960_/A _6436_/Y vssd1 vssd1 vccd1 vccd1 _6437_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6332__B1 _6336_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5135__B2 _6497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6883__A1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6883__B2 _6879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6368_ _6368_/A1 _8310_/B input76/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6368_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8107_ _8097_/Y _7875_/X _8098_/Y _7874_/X _8106_/Y vssd1 vssd1 vccd1 vccd1 _8107_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5319_ _5317_/Y _5318_/Y _8150_/A vssd1 vssd1 vccd1 vccd1 _5320_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8624__A2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6299_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6299_/Y sky130_fd_sc_hd__inv_2
Xinput305 sports_i[45] vssd1 vssd1 vccd1 vccd1 _7936_/A sky130_fd_sc_hd__buf_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkbuf_4
Xinput316 sports_i[55] vssd1 vssd1 vccd1 vccd1 _8072_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__5438__A2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__buf_2
Xinput327 sports_i[65] vssd1 vssd1 vccd1 vccd1 _8234_/B2 sky130_fd_sc_hd__clkbuf_2
X_8038_ _8028_/Y _5185_/A _8029_/Y _5077_/A _8037_/X vssd1 vssd1 vccd1 vccd1 _8039_/A
+ sky130_fd_sc_hd__a221o_2
Xinput338 sports_i[75] vssd1 vssd1 vccd1 vccd1 _7881_/A sky130_fd_sc_hd__clkbuf_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput349 sports_i[85] vssd1 vssd1 vccd1 vccd1 _8024_/B1 sky130_fd_sc_hd__buf_2
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4646__B1 _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5322__B _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6938__A2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7596__C1 _7595_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6434__A _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8560__A1 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4889__A _5130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5484__S _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7265__A _7265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8312__A1 _7788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 _7174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5126__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8795__S _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5126__B2 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4401__B _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8863__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6874__A1 _6866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5677__A2 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7431__C _7432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output417_A _8109_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8379__B2 _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8543__B _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6929__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7051__A1 _6507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6063__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7339__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5670_ _6780_/A _5670_/B vssd1 vssd1 vccd1 vccd1 _5670_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7354__A2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5365__A1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4621_ hold20/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4943_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_115_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5365__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7340_ _5064_/B _7723_/B _7339_/X vssd1 vssd1 vccd1 vccd1 _7340_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4552_ _4552_/A _4552_/B vssd1 vssd1 vccd1 vccd1 _4553_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8303__A1 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7106__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8303__B2 _7798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7271_ _7271_/A vssd1 vssd1 vccd1 vccd1 _7271_/X sky130_fd_sc_hd__buf_1
X_4483_ _4478_/Y _4480_/Y _4481_/Y _4482_/Y _7852_/A vssd1 vssd1 vccd1 vccd1 _4484_/B
+ sky130_fd_sc_hd__a41o_1
XANTENNA__4311__B _8180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6222_ _6937_/A _6234_/B _6221_/Y _5128_/A vssd1 vssd1 vccd1 vccd1 _6222_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_122_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6865__A1 _6028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6865__B2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8067__B1 _8067_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7622__B _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6153_ _6149_/Y _6152_/Y _7852_/A vssd1 vssd1 vccd1 vccd1 _6154_/A sky130_fd_sc_hd__mux2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8606__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5139_/A _8271_/A _5140_/A _4913_/A _5103_/X vssd1 vssd1 vccd1 vccd1 _5105_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7814__B1 _7814_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6084_ _6891_/A _6084_/B vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__and2_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6093__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5035_ _5046_/A _8335_/B _5047_/A _4913_/A _5034_/X vssd1 vssd1 vccd1 vccd1 _5064_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6953__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5840__A2 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8453__B _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6254__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6986_ _6355_/X _6467_/X _6985_/X vssd1 vssd1 vccd1 vccd1 _6986_/X sky130_fd_sc_hd__o21a_1
XANTENNA__8790__A1 _8464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7593__A2 _6809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8790__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5937_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5937_/Y sky130_fd_sc_hd__inv_2
X_8725_ _8725_/A vssd1 vssd1 vccd1 vccd1 _8725_/X sky130_fd_sc_hd__buf_4
XFILLER_0_119_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8656_ _8655_/X _8451_/A _8690_/S vssd1 vssd1 vccd1 vccd1 _8657_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5868_ _5274_/X _5928_/A1 _5275_/X input54/X vssd1 vssd1 vccd1 vccd1 _5868_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8542__A1 _8190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8542__B2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7607_ _8759_/A _7607_/B vssd1 vssd1 vccd1 vccd1 _7607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4819_ _4819_/A _4821_/A _4819_/C vssd1 vssd1 vccd1 vccd1 _8887_/A sky130_fd_sc_hd__nand3_1
X_8587_ _8621_/S vssd1 vssd1 vccd1 vccd1 _8685_/B sky130_fd_sc_hd__buf_4
XFILLER_0_8_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5799_ _6771_/A vssd1 vssd1 vccd1 vccd1 _6762_/A sky130_fd_sc_hd__inv_2
XFILLER_0_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7538_ _7535_/X _7512_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _7538_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5317__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7469_ _5465_/Y _7542_/A _7694_/A _5454_/B _7468_/Y vssd1 vssd1 vccd1 vccd1 _7469_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7532__B _7532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput102 mports_i[191] vssd1 vssd1 vccd1 vccd1 _5543_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__5333__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput113 mports_i[200] vssd1 vssd1 vccd1 vccd1 _5792_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput124 mports_i[210] vssd1 vssd1 vccd1 vccd1 _6089_/A1 sky130_fd_sc_hd__buf_2
Xinput135 mports_i[220] vssd1 vssd1 vccd1 vccd1 _6309_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput146 mports_i[25] vssd1 vssd1 vccd1 vccd1 _5596_/A sky130_fd_sc_hd__clkbuf_4
Xinput157 mports_i[35] vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__clkbuf_4
Xinput168 mports_i[45] vssd1 vssd1 vccd1 vccd1 _6227_/A sky130_fd_sc_hd__buf_2
Xinput179 mports_i[55] vssd1 vssd1 vccd1 vccd1 _6388_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5044__B1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8781__A1 _8423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7336__A2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8533__A1 _8175_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7707__B _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6611__B _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6103__S _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4412__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput609 _5717_/X vssd1 vssd1 vccd1 vccd1 sports_o[197] sky130_fd_sc_hd__buf_12
XFILLER_0_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8836__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8257__C _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5822__A2 _5772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7024__A1 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8221__B1 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6840_ _6432_/X _6839_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6840_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6074__A _6074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5586__A1 _5562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6771_ _6771_/A _7536_/B vssd1 vssd1 vccd1 vccd1 _7558_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6783__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8510_ _8510_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8510_/Y sky130_fd_sc_hd__nand2_1
X_5722_ _5722_/A vssd1 vssd1 vccd1 vccd1 _5722_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7327__A2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8441_ _8441_/A _8441_/B vssd1 vssd1 vccd1 vccd1 _8441_/Y sky130_fd_sc_hd__nand2_1
X_5653_ _5661_/A _4929_/A _5662_/A _4932_/A _5652_/X vssd1 vssd1 vccd1 vccd1 _6743_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7907__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4604_ _4604_/A _4612_/B _4612_/C vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8372_ _8441_/B _8346_/A _8414_/A _8759_/B vssd1 vssd1 vccd1 vccd1 _8372_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5584_ _6284_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5584_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7323_ _7323_/A vssd1 vssd1 vccd1 vccd1 _7323_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4535_ _4535_/A vssd1 vssd1 vccd1 vccd1 _4535_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7254_ _7254_/A vssd1 vssd1 vccd1 vccd1 _7254_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4466_ _8189_/B _4461_/X _4465_/X vssd1 vssd1 vccd1 vccd1 _4466_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6205_ _6229_/A2 _8271_/B input66/X _4917_/A vssd1 vssd1 vccd1 vccd1 _6205_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7352__B _7352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7185_ _6828_/A _7138_/X _7183_/X _7184_/X vssd1 vssd1 vccd1 vccd1 _7185_/X sky130_fd_sc_hd__o22a_2
X_4397_ _4397_/A _7683_/B vssd1 vssd1 vccd1 vccd1 _4398_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6136_ _6136_/A1 _4935_/A input62/X _4939_/A vssd1 vssd1 vccd1 vccd1 _6136_/X sky130_fd_sc_hd__o22a_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6224_/S _6058_/A _6057_/X _6066_/X vssd1 vssd1 vccd1 vccd1 _6067_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8464__A _8464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5018_ _7852_/A vssd1 vssd1 vccd1 vccd1 _8189_/A sky130_fd_sc_hd__buf_8
XFILLER_0_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8212__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout732_A input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5577__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _6467_/X _6310_/X _6450_/A vssd1 vssd1 vccd1 vccd1 _6969_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8708_ _8829_/S vssd1 vssd1 vccd1 vccd1 _8806_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8639_ _8390_/A _8577_/X _8637_/X _8638_/X vssd1 vssd1 vccd1 vccd1 _8639_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6431__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5328__A _5328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7435__A2_N _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8358__B _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5501__A1 _6679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5501__B2 _5500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5998__A _6852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8069__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7006__A1 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8203__B1 _8210_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7006__B2 _4408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8754__A1 _8379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7557__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8821__B _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6622__A _6622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5238__A _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7190__A0 _7189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5740__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput406 _7974_/X vssd1 vssd1 vccd1 vccd1 mports_o[13] sky130_fd_sc_hd__buf_12
XFILLER_0_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput417 _8109_/X vssd1 vssd1 vccd1 vccd1 mports_o[23] sky130_fd_sc_hd__buf_12
XFILLER_0_50_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput428 _8254_/X vssd1 vssd1 vccd1 vccd1 mports_o[33] sky130_fd_sc_hd__buf_12
X_4320_ _4320_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _4321_/B sky130_fd_sc_hd__nand2_1
Xoutput439 _8342_/X vssd1 vssd1 vccd1 vccd1 mports_o[43] sky130_fd_sc_hd__buf_12
XANTENNA__4796__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6296__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7172__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7796__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7941_ _7944_/A1 _5780_/X _7944_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7941_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__6516__B _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7872_ _7872_/A vssd1 vssd1 vccd1 vccd1 _7872_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4317__A _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8745__A1 _7888_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5559__A1 _5558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6823_ _6941_/A _5893_/A _8574_/B vssd1 vssd1 vccd1 vccd1 _6835_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__5559__B2 _5544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6220__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6754_ _5744_/X _6908_/B _6746_/Y _6512_/X _6753_/X vssd1 vssd1 vccd1 vccd1 _6754_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5705_ _6212_/A _5625_/A _5108_/A _5704_/Y _5136_/X vssd1 vssd1 vccd1 vccd1 _5705_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6685_ _6681_/Y _6683_/X _6684_/X _5530_/X _6429_/S vssd1 vssd1 vccd1 vccd1 _6685_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6508__B1 _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5636_ _5591_/A _4929_/A _5592_/A _4932_/A _5635_/X vssd1 vssd1 vccd1 vccd1 _5644_/A
+ sky130_fd_sc_hd__o221a_4
X_8424_ _8424_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8424_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7181__A0 _7179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8355_ _7942_/Y _8299_/X _8354_/Y _8304_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8355_/X
+ sky130_fd_sc_hd__a221o_1
X_5567_ _6689_/S _5560_/Y _5566_/Y vssd1 vssd1 vccd1 vccd1 _5568_/A sky130_fd_sc_hd__a21o_1
XANTENNA__5731__A1 _5011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4987__A _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5731__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7306_ _7306_/A vssd1 vssd1 vccd1 vccd1 _7678_/A sky130_fd_sc_hd__inv_2
X_4518_ _4518_/A _6342_/A vssd1 vssd1 vccd1 vccd1 _4518_/Y sky130_fd_sc_hd__nor2_1
X_8286_ _8567_/B _8284_/Y _8285_/X vssd1 vssd1 vccd1 vccd1 _8286_/X sky130_fd_sc_hd__o21a_1
X_5498_ _5435_/A _5191_/A _5436_/A _5102_/A _5497_/X vssd1 vssd1 vccd1 vccd1 _5498_/X
+ sky130_fd_sc_hd__o221a_4
XANTENNA__8178__B _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6287__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7484__A1 _5544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7237_ _6234_/A _7004_/X _6944_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7237_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7484__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4449_ _4449_/A vssd1 vssd1 vccd1 vccd1 _4449_/Y sky130_fd_sc_hd__inv_2
X_7168_ _6770_/A _7138_/X _7166_/X _7167_/X vssd1 vssd1 vccd1 vccd1 _7168_/X sky130_fd_sc_hd__o22a_2
XANTENNA__6039__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6119_ _6875_/B _6041_/X _6118_/Y vssd1 vssd1 vccd1 vccd1 _6119_/Y sky130_fd_sc_hd__o21ai_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4926__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8194__A _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7099_ _7451_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7099_/X sky130_fd_sc_hd__and2_1
XANTENNA__7787__A2 _7791_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6426__B _6511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8736__A1 _7837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7539__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6747__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6442__A _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8369__A _8369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7475__A1 _6671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8672__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7475__B2 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8976__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7720__B _7720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6617__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7212__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__A1 _5825_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4461__A1 _4312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8727__A1 _8320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5410__B1 _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7167__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6470_ _6470_/A _6470_/B vssd1 vssd1 vccd1 vccd1 _6470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7163__B1 _7162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7702__A2 _7359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5421_ _5465_/A _6017_/A _5077_/A _6648_/B vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_152_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8140_ _8140_/A _8151_/A vssd1 vssd1 vccd1 vccd1 _8141_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5352_ _5352_/A vssd1 vssd1 vccd1 vccd1 _5353_/A sky130_fd_sc_hd__inv_2
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6269__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4303_ _4303_/A vssd1 vssd1 vccd1 vccd1 _4591_/B sky130_fd_sc_hd__buf_4
X_8071_ _8071_/A vssd1 vssd1 vccd1 vccd1 _8071_/Y sky130_fd_sc_hd__inv_2
X_5283_ _7829_/A _6576_/B _5282_/Y vssd1 vssd1 vccd1 vccd1 _5283_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7022_ _7089_/A vssd1 vssd1 vccd1 vccd1 _7138_/A sky130_fd_sc_hd__inv_6
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7630__B _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8973_ _8976_/CLK _8973_/D fanout733/X vssd1 vssd1 vccd1 vccd1 _8973_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7924_ _7931_/A1 _4946_/A _7931_/B1 _5119_/A vssd1 vssd1 vccd1 vccd1 _7924_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_78_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8718__A1 _7771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8718__B2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7855_ _7840_/Y _5780_/A _7841_/Y _5079_/A _7854_/X vssd1 vssd1 vccd1 vccd1 _7856_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7358__A _7372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6806_ _6795_/X _6450_/X _6800_/Y _6801_/X _6805_/X vssd1 vssd1 vccd1 vccd1 _6806_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_19_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4998_ _6356_/S vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__buf_8
X_7786_ _7791_/A1 _6513_/A _7791_/B1 _5171_/B _7785_/X vssd1 vssd1 vccd1 vccd1 _7786_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__7941__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5952__A1 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6737_ _6737_/A vssd1 vssd1 vccd1 vccd1 _7153_/A sky130_fd_sc_hd__inv_2
XANTENNA__5952__B2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6668_ _6668_/A _6694_/B vssd1 vssd1 vccd1 vccd1 _6668_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7154__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8407_ _8407_/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8407_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5619_ _5659_/A _7299_/A _6281_/S _7524_/A vssd1 vssd1 vccd1 vccd1 _5619_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8189__A _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6599_ _5328_/A _6510_/A _5330_/Y _6512_/X vssd1 vssd1 vccd1 vccd1 _6599_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5180__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8338_ _8352_/A _8304_/A _7916_/Y _8299_/A _8269_/A vssd1 vssd1 vccd1 vccd1 _8338_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7457__A1 _6648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8269_ _8269_/A vssd1 vssd1 vccd1 vccd1 _8496_/S sky130_fd_sc_hd__buf_6
XANTENNA__8654__B1 _8455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7457__B2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5468__B1 _5511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7821__A _7821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6680__A2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5341__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7090__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4994__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7917__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7932__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4404__B _8968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5516__A _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7207__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7448__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8645__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output447_A _8422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7999__A2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6120__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7450__B _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6959__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8955__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5970_ _5970_/A _7847_/A vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _6181_/B vssd1 vssd1 vccd1 vccd1 _6212_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_48_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8176__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4852_ _8967_/D _8966_/D vssd1 vssd1 vccd1 vccd1 _4858_/A sky130_fd_sc_hd__nor2_1
XANTENNA__6187__A1 _6908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7640_ _7640_/A _7640_/B _7640_/C vssd1 vssd1 vccd1 vccd1 _7640_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__6187__B2 _7683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5395__C1 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7571_ _6770_/A _7389_/A _7569_/X _7326_/A _7570_/Y vssd1 vssd1 vccd1 vccd1 _7571_/X
+ sky130_fd_sc_hd__a221o_1
X_4783_ _4783_/A _4786_/A vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5934__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6522_ _6694_/B vssd1 vssd1 vccd1 vccd1 _6851_/B sky130_fd_sc_hd__buf_6
XANTENNA__8501__S _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6453_ _8189_/A _6443_/A _4973_/Y vssd1 vssd1 vccd1 vccd1 _6481_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7687__B2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5404_ _5401_/Y _4885_/A _5402_/Y _4890_/A _5403_/Y vssd1 vssd1 vccd1 vccd1 _6646_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4330__A _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6384_ _6388_/A1 _8516_/B input15/X _4913_/X _6383_/X vssd1 vssd1 vccd1 vccd1 _6385_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8123_ _8123_/A vssd1 vssd1 vccd1 vccd1 _8123_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_100_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5335_ _6711_/S vssd1 vssd1 vccd1 vccd1 _6837_/A sky130_fd_sc_hd__buf_6
XANTENNA__8100__A2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8054_ _8054_/A1 _7876_/X _8054_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _8054_/Y sky130_fd_sc_hd__o22ai_2
X_5266_ _5266_/A vssd1 vssd1 vccd1 vccd1 _5266_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6111__A1 _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7005_ _7059_/A vssd1 vssd1 vccd1 vccd1 _7272_/A sky130_fd_sc_hd__inv_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5197_ _7311_/A vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__buf_8
XFILLER_0_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8956_ _8976_/CLK _8956_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5622__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7907_ _7777_/X _7906_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _7907_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8887_ _8887_/A _8887_/B vssd1 vssd1 vccd1 vccd1 _8888_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8167__A2 _8172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7088__A _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7838_ _7837_/X _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _7838_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7914__A2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7769_ _7769_/A vssd1 vssd1 vccd1 vccd1 _7769_/X sky130_fd_sc_hd__buf_12
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7127__B1 _7126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8324__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5336__A _7432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6350__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5153__A2 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6350__B2 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8890__A3 _8264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8627__B1 _8386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6638__C1 _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7551__A _7551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8978__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7850__A1 _7840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7850__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5861__B1 _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7602__A1 _5930_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7602__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6956__A3 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6169__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7905__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5916__A1 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__B2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8321__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6630__A _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8866__B1 _7372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8330__A2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8618__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ input86/X _4935_/A input24/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8094__B2 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5051_ _5008_/A _5050_/Y _6470_/B vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8397__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8810_ _8809_/X _8525_/Y _8829_/S vssd1 vssd1 vccd1 vccd1 _8811_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8741_ _7862_/A _8725_/X _8740_/X vssd1 vssd1 vccd1 vccd1 _8741_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_149_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4958__A2 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5953_ _5944_/X _5715_/B _6356_/S _5952_/X vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8149__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4904_ _5174_/A vssd1 vssd1 vccd1 vccd1 _5672_/A sky130_fd_sc_hd__inv_2
X_5884_ _5902_/A1 _4934_/A input53/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__o22a_1
X_8672_ _8698_/B _8515_/A _8590_/X vssd1 vssd1 vccd1 vccd1 _8672_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7623_ _7694_/A _7623_/B vssd1 vssd1 vccd1 vccd1 _7623_/Y sky130_fd_sc_hd__nor2_1
X_4835_ _4436_/A _8240_/A _6980_/B _4834_/X _7384_/A vssd1 vssd1 vccd1 vccd1 _4835_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_117_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4766_ _8240_/A _6980_/B _4765_/Y _4764_/B vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__a31o_1
X_7554_ _7378_/X _5744_/X _7683_/C vssd1 vssd1 vccd1 vccd1 _7556_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6505_ _6924_/A _6505_/B vssd1 vssd1 vccd1 vccd1 _6505_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7485_ _7484_/X _5530_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7486_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4697_ _4697_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4751_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6332__A1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5135__A2 _6499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6436_ _6436_/A vssd1 vssd1 vccd1 vccd1 _6436_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6332__B2 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6367_ _6367_/A _6367_/B vssd1 vssd1 vccd1 vccd1 _6367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5318_ _5356_/B _6868_/B vssd1 vssd1 vccd1 vccd1 _5318_/Y sky130_fd_sc_hd__nand2_1
X_8106_ _8106_/A1 _7876_/X _8106_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _8106_/Y sky130_fd_sc_hd__o22ai_4
X_6298_ _7729_/B _6059_/B _7733_/B _8857_/B _7725_/B vssd1 vssd1 vccd1 vccd1 _6298_/X
+ sky130_fd_sc_hd__a221o_1
Xinput306 sports_i[46] vssd1 vssd1 vccd1 vccd1 _7949_/A sky130_fd_sc_hd__clkbuf_1
Xinput317 sports_i[56] vssd1 vssd1 vccd1 vccd1 _8084_/A sky130_fd_sc_hd__buf_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _6584_/A _6181_/B vssd1 vssd1 vccd1 vccd1 _5249_/Y sky130_fd_sc_hd__nand2_1
X_8037_ _6500_/A _8031_/Y _8030_/Y _7769_/A vssd1 vssd1 vccd1 vccd1 _8037_/X sky130_fd_sc_hd__a22o_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput328 sports_i[66] vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__buf_4
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xinput339 sports_i[76] vssd1 vssd1 vccd1 vccd1 _7905_/B1 sky130_fd_sc_hd__clkbuf_4
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4646__A1 _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4646__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6399__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8939_ hold42/X vssd1 vssd1 vccd1 vccd1 _8965_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__6434__B _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7899__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8560__A2 _8222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6450__A _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6571__A1 _6567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6571__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6323__A1 _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5126__A2 _7345_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7281__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8076__B2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6609__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8379__A2 _7912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7051__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8000__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4620_ hold18/X vssd1 vssd1 vccd1 vccd1 _4824_/B sky130_fd_sc_hd__clkinv_4
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5365__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4551_ _4554_/A _4551_/B _7707_/C vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8303__A2 _7832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7270_ _7269_/Y _7733_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7271_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_52_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4482_ _4482_/A _4566_/A vssd1 vssd1 vccd1 vccd1 _4482_/Y sky130_fd_sc_hd__nand2_1
X_6221_ _6221_/A vssd1 vssd1 vccd1 vccd1 _6221_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6865__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4876__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7191__A _7191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4876__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6152_ _6192_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6152_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8067__A1 _8067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8067__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5103_ input87/X _8271_/B input25/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__o22a_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7814__A1 _7814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6083_ _5999_/B _7209_/A _6082_/X _5174_/A vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__a22o_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7814__B2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ input84/X _8716_/B input21/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__o22a_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7578__B1 _7576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6985_ _6349_/X _6994_/B _7278_/A _6989_/B _7000_/S vssd1 vssd1 vccd1 vccd1 _6985_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8790__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8724_ _8724_/A vssd1 vssd1 vccd1 vccd1 _8725_/A sky130_fd_sc_hd__inv_2
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _5936_/A vssd1 vssd1 vccd1 vccd1 _5936_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8655_ _8654_/X _8055_/Y _8689_/S vssd1 vssd1 vccd1 vccd1 _8655_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5867_ _5867_/A vssd1 vssd1 vccd1 vccd1 _5867_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8542__A2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7366__A _7686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7606_ _7606_/A _7606_/B vssd1 vssd1 vccd1 vccd1 _7606_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4818_ _4818_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _8877_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8586_ _8689_/S vssd1 vssd1 vccd1 vccd1 _8621_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5798_ _7570_/B _6211_/B vssd1 vssd1 vccd1 vccd1 _5798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7537_ _7536_/B _6733_/A _7535_/X _7536_/Y vssd1 vssd1 vccd1 vccd1 _7537_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4749_ _4770_/C vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__inv_2
XANTENNA__4502__B hold10/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7502__B1 _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7468_ _7468_/A _7640_/B vssd1 vssd1 vccd1 vccd1 _7468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6419_ _8174_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _6528_/A sky130_fd_sc_hd__nand2_4
X_7399_ _7701_/A _6567_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7401_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput103 mports_i[192] vssd1 vssd1 vccd1 vccd1 _5557_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__7805__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6608__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5333__B _5333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput114 mports_i[201] vssd1 vssd1 vccd1 vccd1 _5787_/A1 sky130_fd_sc_hd__buf_2
Xinput125 mports_i[211] vssd1 vssd1 vccd1 vccd1 _6104_/A1 sky130_fd_sc_hd__buf_2
Xinput136 mports_i[221] vssd1 vssd1 vccd1 vccd1 _6315_/B sky130_fd_sc_hd__clkbuf_4
Xinput147 mports_i[26] vssd1 vssd1 vccd1 vccd1 _5661_/A sky130_fd_sc_hd__clkbuf_4
Xinput158 mports_i[36] vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__clkbuf_4
Xinput169 mports_i[46] vssd1 vssd1 vccd1 vccd1 _6248_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7569__B1 _6779_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7033__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5044__A1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6241__B1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6792__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8533__A2 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6180__A _6180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7707__C _7707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4412__B _6411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7723__B _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8049__A1 _8054_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7257__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5283__A1 _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8221__A1 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7024__A2 _4963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8221__B2 _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5035__A1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5035__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6770_ _6770_/A vssd1 vssd1 vccd1 vccd1 _6770_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6783__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7980__B1 _7985_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ _5738_/C _5827_/B _7297_/B vssd1 vssd1 vccd1 vccd1 _5721_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6802__B _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8440_ _8439_/Y _8412_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8440_/X sky130_fd_sc_hd__mux2_1
X_5652_ _5697_/A1 _4935_/A input46/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5652_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4603_ _4603_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _4612_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8371_ _8371_/A vssd1 vssd1 vccd1 vccd1 _8414_/A sky130_fd_sc_hd__inv_2
XANTENNA__4322__B _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5583_ _6697_/B vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__inv_2
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7322_ _7321_/X _4966_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7323_/A sky130_fd_sc_hd__mux2_1
X_4534_ _4839_/A _4534_/B vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6838__A2 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7253_ _6287_/X _7138_/A _7252_/X vssd1 vssd1 vccd1 vccd1 _7254_/A sky130_fd_sc_hd__o21ai_1
X_4465_ _4482_/A _4318_/B _4658_/A _5077_/A vssd1 vssd1 vccd1 vccd1 _4465_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5434__A _6646_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6204_ _7707_/B _6099_/Y _6203_/Y vssd1 vssd1 vccd1 vccd1 _6204_/Y sky130_fd_sc_hd__o21ai_1
X_7184_ _6811_/B _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7184_/X sky130_fd_sc_hd__a21o_1
X_4396_ _4425_/B _4425_/C _4407_/C vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__nand3_1
X_6135_ _6132_/X _6133_/Y _6134_/X _6170_/A _6102_/A vssd1 vssd1 vccd1 vccd1 _6135_/X
+ sky130_fd_sc_hd__a32o_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7799__B1 _4566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6266_/A _6060_/Y _6064_/Y _6065_/X vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__o211a_1
XANTENNA__8464__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5017_ _6284_/A _5019_/A vssd1 vssd1 vccd1 vccd1 _5017_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6471__B1 _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__A1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8480__A _8480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5577__A2 _5587_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6774__A1 _7167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6968_ _6968_/A _6968_/B vssd1 vssd1 vccd1 vccd1 _6968_/X sky130_fd_sc_hd__or2_1
XANTENNA__7971__B1 _7971_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6774__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8707_ _8724_/A vssd1 vssd1 vccd1 vccd1 _8829_/S sky130_fd_sc_hd__buf_6
X_5919_ _6128_/B _6828_/A _5136_/X _5918_/Y vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6899_ _6899_/A _6899_/B vssd1 vssd1 vccd1 vccd1 _6899_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5609__A _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8638_ _8698_/B _8772_/B _8590_/X vssd1 vssd1 vccd1 vccd1 _8638_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_118_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8569_ _4661_/A _8323_/X _8568_/X vssd1 vssd1 vccd1 vccd1 _8569_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7487__C1 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7035__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5501__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8203__A1 _8210_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7006__A2 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8754__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8390__A _8390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5519__A _5519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4423__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7190__A1 _5899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5740__A2 _7544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput407 _7988_/X vssd1 vssd1 vccd1 vccd1 mports_o[14] sky130_fd_sc_hd__buf_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput418 _8122_/X vssd1 vssd1 vccd1 vccd1 mports_o[24] sky130_fd_sc_hd__buf_12
Xoutput429 _8267_/X vssd1 vssd1 vccd1 vccd1 mports_o[34] sky130_fd_sc_hd__buf_12
XFILLER_0_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8690__A1 _8200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8442__A1 _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8284__B _8284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7940_ _7935_/Y _6965_/A _7936_/Y _8163_/A _7939_/Y vssd1 vssd1 vccd1 vccd1 _8351_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7871_ _7864_/Y _7769_/X _7865_/Y _6500_/X _7870_/Y vssd1 vssd1 vccd1 vccd1 _7871_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__4317__B _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6205__B1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8504__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6822_ _6813_/Y _6450_/X _6815_/X _6817_/Y _6821_/X vssd1 vssd1 vccd1 vccd1 _6822_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__5559__A2 _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6813__A _6813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6753_ _6747_/X _6924_/A _6748_/X _6752_/Y vssd1 vssd1 vccd1 vccd1 _6753_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5704_ _5704_/A vssd1 vssd1 vccd1 vccd1 _5704_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6508__A1 _6503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6684_ _6801_/A _5544_/X _6450_/A vssd1 vssd1 vccd1 vccd1 _6684_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_115_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8423_ _8423_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8423_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5148__B _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5635_ _5635_/A1 _4935_/A input42/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5635_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5716__C1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7181__A1 _5853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8354_ _8354_/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8354_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5566_ _6689_/S _5566_/B vssd1 vssd1 vccd1 vccd1 _5566_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4987__B _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7305_ _7532_/A _7364_/A vssd1 vssd1 vccd1 vccd1 _7306_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_130_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4517_ _4517_/A _4517_/B vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__nand2_1
X_5497_ _5497_/A1 _5192_/A input38/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5497_/X sky130_fd_sc_hd__o22a_1
X_8285_ _7809_/X _8304_/A _7811_/X _8299_/A _8496_/S vssd1 vssd1 vccd1 vccd1 _8285_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7236_ _7236_/A vssd1 vssd1 vccd1 vccd1 _7236_/X sky130_fd_sc_hd__buf_1
XANTENNA__7484__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8681__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4448_ _4453_/A hold32/X vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5495__A1 _5497_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5495__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8475__A _8475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4379_ _4300_/Y _4377_/X _8917_/S vssd1 vssd1 vccd1 vccd1 _4380_/B sky130_fd_sc_hd__a21oi_1
X_7167_ _7167_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7167_/X sky130_fd_sc_hd__and2_1
XFILLER_0_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6118_ _6118_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _6118_/Y sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7098_/A vssd1 vssd1 vccd1 vccd1 _7098_/X sky130_fd_sc_hd__buf_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _5274_/X _6104_/A1 _5275_/X input61/X vssd1 vssd1 vccd1 vccd1 _6049_/Y sky130_fd_sc_hd__a22oi_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8197__B1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8736__A2 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6747__A1 _7544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7944__B1 _7944_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6747__B2 _5765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6869__S _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8369__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5074__A _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8672__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7475__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6617__B _7094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8188__A0 _8180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8945__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8727__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7729__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6738__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output594_A _5332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5410__A1 _5011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5961__A2 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7163__A1 _6771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5420_ _5401_/A _4868_/A _5402_/A _5089_/A _5419_/X vssd1 vssd1 vccd1 vccd1 _6648_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6910__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7183__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5351_ _6622_/A _8151_/B _5197_/X _5317_/A vssd1 vssd1 vccd1 vccd1 _5352_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8112__B1 _8119_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4302_ _6312_/A vssd1 vssd1 vccd1 vccd1 _5827_/B sky130_fd_sc_hd__inv_6
XANTENNA__8663__A1 _8476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8070_ _7975_/X _8491_/A _8066_/X _8069_/X vssd1 vssd1 vccd1 vccd1 _8070_/X sky130_fd_sc_hd__a22o_2
X_5282_ _7071_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5282_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5477__A1 _5718_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5477__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7021_ _6440_/A _7019_/X _6456_/A _7288_/B _7012_/S vssd1 vssd1 vccd1 vccd1 _7021_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6674__B1 _6672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8295__A _8295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _8967_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__8415__A1 _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6019__S _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8972_ _8976_/CLK _8972_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__4988__B1 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7923_ _7923_/A vssd1 vssd1 vccd1 vccd1 _7923_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__8718__A2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7854_ _7852_/Y _7853_/Y hold23/A vssd1 vssd1 vccd1 vccd1 _7854_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6543__A _6543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7926__B1 _7931_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6805_ _5853_/X _6510_/A _6804_/Y _6512_/A vssd1 vssd1 vccd1 vccd1 _6805_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7785_ _6079_/A _7790_/A2 _7304_/A _7790_/B2 vssd1 vssd1 vccd1 vccd1 _7785_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_92_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _4997_/A vssd1 vssd1 vccd1 vccd1 _4997_/X sky130_fd_sc_hd__buf_1
XFILLER_0_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5159__A _5159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6736_ _6506_/A _7544_/A _6449_/A vssd1 vssd1 vccd1 vccd1 _6736_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_147_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5952__A2 _5860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6689__S _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4998__A _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6667_ _6642_/Y _6666_/Y _6870_/S vssd1 vssd1 vccd1 vccd1 _6667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7154__A1 _5738_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8406_ _8406_/A vssd1 vssd1 vccd1 vccd1 _8407_/A sky130_fd_sc_hd__inv_2
XFILLER_0_131_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5165__B1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5618_ _5909_/B _5595_/Y _5617_/Y _5997_/B vssd1 vssd1 vccd1 vccd1 _5618_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6598_ _7415_/B _6925_/B vssd1 vssd1 vccd1 vccd1 _6598_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8189__B _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5606__B _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8337_ _8337_/A vssd1 vssd1 vccd1 vccd1 _8337_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4510__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5549_ _5549_/A vssd1 vssd1 vccd1 vccd1 _5549_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7457__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8268_ _8567_/B vssd1 vssd1 vccd1 vccd1 _8269_/A sky130_fd_sc_hd__inv_2
XANTENNA__8654__B2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5468__A1 _5510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5468__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6665__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7219_ _6913_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7219_/X sky130_fd_sc_hd__a21o_1
X_8199_ _8194_/A _8209_/A2 _8845_/C _8198_/X vssd1 vssd1 vccd1 vccd1 _8199_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4632__A1_N hold10/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5341__B _7094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4979__B1 _4674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__A1 _5640_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7917__B1 _7916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__A _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7393__B2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7145__A1 _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6900__B _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8645__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7448__A2 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5459__A1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5459__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6120__A2 _6141_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6959__A1 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7459__A _7459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4920_ _6312_/A _7309_/B vssd1 vssd1 vccd1 vccd1 _6181_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ _4866_/A _4863_/B vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6187__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7570_ _7673_/A _7570_/B vssd1 vssd1 vccd1 vccd1 _7570_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5934__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4782_ _4782_/A _4788_/B vssd1 vssd1 vccd1 vccd1 _4783_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6521_ _7356_/B _6908_/B _5124_/X _6512_/X _6520_/X vssd1 vssd1 vccd1 vccd1 _6521_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7136__A1 _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6452_ _4966_/X _6429_/S _6445_/X _6451_/X vssd1 vssd1 vccd1 vccd1 _6452_/X sky130_fd_sc_hd__a22o_2
XANTENNA__7687__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__A1 _5661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5403_ _5274_/X input98/X _5275_/X input36/X vssd1 vssd1 vccd1 vccd1 _5403_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_141_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6383_ _6387_/A1 _8716_/B input77/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6383_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_24_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4330__B _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7922__A _7922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8122_ _7975_/X _8519_/A _8118_/X _8121_/X vssd1 vssd1 vccd1 vccd1 _8122_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_11_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5334_ _5011_/Y _5333_/Y _5013_/Y vssd1 vssd1 vccd1 vccd1 _5334_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6647__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8053_ _8455_/A _7954_/X _8458_/A _7826_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _8053_/X
+ sky130_fd_sc_hd__a221o_1
X_5265_ _5265_/A vssd1 vssd1 vccd1 vccd1 _5265_/Y sky130_fd_sc_hd__inv_2
X_7004_ _7059_/A vssd1 vssd1 vccd1 vccd1 _7004_/X sky130_fd_sc_hd__buf_6
X_5196_ _5196_/A vssd1 vssd1 vccd1 vccd1 _7368_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8955_ _8967_/CLK _8955_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7906_ _7896_/Y _7874_/A _7897_/Y _8174_/A _7905_/Y vssd1 vssd1 vccd1 vccd1 _7906_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_149_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8886_ _8886_/A _8899_/A _8899_/B vssd1 vssd1 vccd1 vccd1 _8886_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_66_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7837_ _7827_/Y _5230_/B _7834_/X _7707_/C _7836_/Y vssd1 vssd1 vccd1 vccd1 _7837_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7768_ _7954_/A vssd1 vssd1 vccd1 vccd1 _7768_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6719_ _6717_/X _6933_/A _6968_/A _6718_/X vssd1 vssd1 vccd1 vccd1 _6719_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_135_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7127__A1 _5558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6720__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8324__B1 _7871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7699_ _7378_/X _6941_/B _7683_/C vssd1 vssd1 vccd1 vccd1 _7701_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8627__A1 _8384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8627__B2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7551__B _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput590 _7109_/X vssd1 vssd1 vccd1 vccd1 sports_o[17] sky130_fd_sc_hd__buf_12
XANTENNA__7850__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5861__A1 _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7602__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6810__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6169__A2 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8563__B1 _8232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7118__A1 _5496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6630__B _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7669__A2 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8079__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8618__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8094__A2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5050_ _5050_/A vssd1 vssd1 vccd1 vccd1 _5050_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5852__A1 _5881_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5852__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8960__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7054__B1 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5604__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8740_ _8315_/A _8820_/B _8829_/S _8739_/X vssd1 vssd1 vccd1 vccd1 _8740_/X sky130_fd_sc_hd__a211o_1
X_5952_ _6084_/B _5860_/A _6854_/B _5096_/A vssd1 vssd1 vccd1 vccd1 _5952_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4903_ _5485_/A _5145_/A vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__nor2_8
X_8671_ _8510_/A _8581_/A _8117_/Y _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8671_/X
+ sky130_fd_sc_hd__a221o_1
X_5883_ _5880_/X _6801_/B _6386_/S vssd1 vssd1 vccd1 vccd1 _5883_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7622_ _7622_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7622_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5368__B1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8512__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4834_ _4420_/Y _4449_/Y _4760_/A vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_63_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7553_ _7552_/X _5765_/X _7749_/S vssd1 vssd1 vccd1 vccd1 _7553_/X sky130_fd_sc_hd__mux2_1
X_4765_ hold32/A _4871_/A vssd1 vssd1 vccd1 vccd1 _4765_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7128__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6504_ _6528_/A vssd1 vssd1 vccd1 vccd1 _6924_/A sky130_fd_sc_hd__buf_6
X_7484_ _5544_/X _7696_/B _7482_/X _7326_/A _7483_/Y vssd1 vssd1 vccd1 vccd1 _7484_/X
+ sky130_fd_sc_hd__a221o_1
X_4696_ _4696_/A _4696_/B vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7419__A1_N _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _6435_/A vssd1 vssd1 vccd1 vccd1 _6436_/A sky130_fd_sc_hd__buf_6
XFILLER_0_141_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6332__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5540__B1 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6366_ input76/X _8579_/C _6368_/A1 _8713_/C _6365_/X vssd1 vssd1 vccd1 vccd1 _6367_/B
+ sky130_fd_sc_hd__a221oi_4
X_8105_ _8503_/A _7954_/X _8104_/Y _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8105_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5317_ _5317_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _5317_/Y sky130_fd_sc_hd__nand2_1
X_6297_ _6299_/A _8491_/B input8/X _4933_/A _6296_/X vssd1 vssd1 vccd1 vccd1 _7725_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6096__A1 _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5172__A _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput307 sports_i[47] vssd1 vssd1 vccd1 vccd1 _7963_/A sky130_fd_sc_hd__clkbuf_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_8036_ _8444_/B vssd1 vssd1 vccd1 vccd1 _8036_/Y sky130_fd_sc_hd__inv_2
Xinput318 sports_i[57] vssd1 vssd1 vccd1 vccd1 _8097_/A sky130_fd_sc_hd__clkbuf_1
X_5248_ _5248_/A vssd1 vssd1 vccd1 vccd1 _6584_/A sky130_fd_sc_hd__inv_2
Xinput329 sports_i[67] vssd1 vssd1 vccd1 vccd1 _8251_/B2 sky130_fd_sc_hd__buf_2
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5843__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4646__A2 _4927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8483__A _8483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5179_ input91/X _8709_/B input28/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_97_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8793__B1 _8480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7099__A _7451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7596__B2 _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8938_ hold41/X _4694_/A _8938_/S vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8869_ hold30/X _8869_/B vssd1 vssd1 vccd1 vccd1 _8872_/A sky130_fd_sc_hd__or2_1
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7827__A _7827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6731__A _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7899__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6571__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5066__B _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6323__A2 _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8945__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8076__A2 _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6087__A1 _6020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6087__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5834__A1 _5011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5834__B2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6906__A _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5810__A _5810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8233__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5598__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7339__B2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8536__B1 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7737__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8000__A2 _7999_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6011__A1 _6089_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6011__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5257__A _7422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550_ hold12/X vssd1 vssd1 vccd1 vccd1 _7707_/C sky130_fd_sc_hd__inv_6
XANTENNA__5770__B1 _5723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4481_ _5077_/A _4481_/B vssd1 vssd1 vccd1 vccd1 _4481_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6220_ _6202_/Y _6402_/A _6211_/Y _6212_/X _6219_/X vssd1 vssd1 vccd1 vccd1 _6220_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__4876__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6151_ input2/X _4870_/A _6158_/A _4953_/X _6150_/X vssd1 vssd1 vccd1 vccd1 _6192_/A
+ sky130_fd_sc_hd__o221a_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8067__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7275__A0 _7274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5102_ _5102_/A vssd1 vssd1 vccd1 vccd1 _8271_/A sky130_fd_sc_hd__buf_8
XANTENNA__6078__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6082_ _6081_/X _7638_/A _6711_/S vssd1 vssd1 vccd1 vccd1 _6082_/X sky130_fd_sc_hd__mux2_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7814__A2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5825__A1 _5825_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5825__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5046_/A _4930_/X _5047_/A _4933_/X _5032_/X vssd1 vssd1 vccd1 vccd1 _7341_/B
+ sky130_fd_sc_hd__o221a_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6816__A _6828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7578__A1 _6788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7578__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4336__A _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6984_ _6984_/A vssd1 vssd1 vccd1 vccd1 _6984_/X sky130_fd_sc_hd__buf_1
XFILLER_0_94_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8723_ _8782_/A vssd1 vssd1 vccd1 vccd1 _8833_/B sky130_fd_sc_hd__buf_4
XFILLER_0_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5935_ _6024_/A _6852_/B vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_137_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8527__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8654_ _8696_/A _8482_/A _8455_/A _8581_/A vssd1 vssd1 vccd1 vccd1 _8654_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6551__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5866_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5866_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7605_ _6827_/A _7696_/B _7602_/X _7603_/X _7604_/Y vssd1 vssd1 vccd1 vccd1 _7605_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4817_ _4817_/A _4817_/B vssd1 vssd1 vccd1 vccd1 _4818_/A sky130_fd_sc_hd__nand2_1
X_8585_ _8589_/A vssd1 vssd1 vccd1 vccd1 _8689_/S sky130_fd_sc_hd__clkinv_4
XFILLER_0_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8968__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5797_ _6689_/S _5791_/X _5796_/Y vssd1 vssd1 vccd1 vccd1 _7570_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7536_ _7536_/A _7536_/B vssd1 vssd1 vccd1 vccd1 _7536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _4786_/B _4748_/B vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7467_ _7110_/A _7668_/B _6668_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _7468_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_98_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4679_ _4693_/A _4693_/B _4694_/A vssd1 vssd1 vccd1 vccd1 _4680_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__7502__A1 _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6305__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7382__A _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6418_ _6925_/B vssd1 vssd1 vccd1 vccd1 _6506_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7398_ _7398_/A vssd1 vssd1 vccd1 vccd1 _7683_/C sky130_fd_sc_hd__buf_4
XFILLER_0_12_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6349_ _6358_/A1 _8480_/B input13/X _4870_/X _6348_/X vssd1 vssd1 vccd1 vccd1 _6349_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6069__A1 _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6069__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput104 mports_i[193] vssd1 vssd1 vccd1 vccd1 _5587_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__7805__A2 _7796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput115 mports_i[202] vssd1 vssd1 vccd1 vccd1 _5825_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput126 mports_i[212] vssd1 vssd1 vccd1 vccd1 _6136_/A1 sky130_fd_sc_hd__buf_2
Xinput137 mports_i[222] vssd1 vssd1 vccd1 vccd1 _6336_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput148 mports_i[27] vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__buf_4
X_8019_ _8024_/A1 _5145_/A _8024_/B1 _5616_/A vssd1 vssd1 vccd1 vccd1 _8019_/Y sky130_fd_sc_hd__o22ai_4
Xinput159 mports_i[37] vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8417__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7321__S _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7569__A1 _7167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7569__B2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6241__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6792__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7741__A1 _6358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7707__D _7707_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5077__A _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5201__C1 _6359_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8297__A2 _8364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5805__A _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8049__A2 _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5807__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output422_A _8197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5283__A2 _6576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6480__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5035__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6232__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7980__A1 _7985_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7980__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5720_ _6743_/A _7316_/A _8924_/B _5741_/A vssd1 vssd1 vccd1 vccd1 _5720_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5651_ _5644_/A _6059_/B _8924_/B _5679_/A vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4602_ _4602_/A _4602_/B vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5743__B1 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8370_ _8369_/Y _8345_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8371_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_142_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5582_ _5580_/X _8755_/C _6837_/A _5999_/B _5581_/Y vssd1 vssd1 vccd1 vccd1 _5582_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7321_ _7320_/X _4963_/X _7749_/S vssd1 vssd1 vccd1 vccd1 _7321_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4533_ _4557_/B _4591_/B _8584_/B vssd1 vssd1 vccd1 vccd1 _4534_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7252_ _7251_/Y _7059_/A _6272_/X _7088_/A _7089_/A vssd1 vssd1 vccd1 vccd1 _7252_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _8166_/A _8189_/B vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_68_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6203_ _6212_/B _7707_/B vssd1 vssd1 vccd1 vccd1 _6203_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_110_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7183_ _7183_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7183_/X sky130_fd_sc_hd__and2_1
X_4395_ _4395_/A _4395_/B vssd1 vssd1 vccd1 vccd1 _4407_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6134_ _6284_/A _6913_/A _6261_/A vssd1 vssd1 vccd1 vccd1 _6134_/X sky130_fd_sc_hd__o21a_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7799__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7799__B2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6212_/A _6063_/A _4949_/A vssd1 vssd1 vccd1 vccd1 _6065_/X sky130_fd_sc_hd__o21a_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6471__A1 _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5016_ _5003_/A _4870_/A _5004_/A _4953_/X _5015_/X vssd1 vssd1 vccd1 vccd1 _5019_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_84_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8212__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8761__A _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6223__A1 _7696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8480__B _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6967_ _6277_/A _6841_/A _6278_/Y _6854_/A _6966_/X vssd1 vssd1 vccd1 vccd1 _6968_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__7971__A1 _7971_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6774__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7971__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5918_ _5918_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _5918_/Y sky130_fd_sc_hd__nand2_1
X_8706_ _8759_/A _8706_/B vssd1 vssd1 vccd1 vccd1 _8724_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6898_ _6897_/Y _6475_/X _6054_/X _6694_/B vssd1 vssd1 vccd1 vccd1 _6899_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_118_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8637_ _8394_/A _8581_/X _7983_/Y _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8637_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5609__B _5609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _5849_/A vssd1 vssd1 vccd1 vccd1 _6818_/A sky130_fd_sc_hd__inv_2
XFILLER_0_134_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8568_ _8567_/B _4607_/A _8497_/S _8567_/Y vssd1 vssd1 vccd1 vccd1 _8568_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5734__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7519_ _7700_/B _7520_/B _5628_/A _7754_/A vssd1 vssd1 vccd1 vccd1 _7519_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_121_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8499_ _8499_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5625__A _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8684__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5360__A _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8739__B1 _7851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8203__A2 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6214__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8390__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5973__B1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7226__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput408 _8001_/X vssd1 vssd1 vccd1 vccd1 mports_o[15] sky130_fd_sc_hd__buf_12
Xoutput419 _8135_/X vssd1 vssd1 vccd1 vccd1 mports_o[25] sky130_fd_sc_hd__buf_12
XFILLER_0_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6150__B1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7750__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5270__A _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6453__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8581__A _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7870_ _7877_/A1 _5780_/X _7877_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7870_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__6205__A1 _6229_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6205__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6821_ _5885_/X _6510_/A _6820_/Y _6512_/A vssd1 vssd1 vccd1 vccd1 _6821_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_89_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6813__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7953__B2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4614__A _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6752_ _5707_/A _6854_/A _6467_/X _6749_/Y _6751_/Y vssd1 vssd1 vccd1 vccd1 _6752_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5703_ _6689_/S _5701_/X _5702_/Y vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6683_ _6924_/A _7476_/A vssd1 vssd1 vccd1 vccd1 _6683_/X sky130_fd_sc_hd__or2_1
XANTENNA__4333__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6508__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8422_ _8323_/X _8415_/Y _8420_/X _8421_/X vssd1 vssd1 vccd1 vccd1 _8422_/X sky130_fd_sc_hd__a22o_2
XANTENNA__4519__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8520__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5634_ _6212_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _5634_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8353_ _8351_/Y _8352_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8354_/A sky130_fd_sc_hd__mux2_1
X_5565_ _5562_/X _7311_/A _8151_/B _5634_/B vssd1 vssd1 vccd1 vccd1 _5566_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7136__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7469__B1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7304_ _7304_/A _8755_/C vssd1 vssd1 vccd1 vccd1 _7364_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4516_ _4516_/A vssd1 vssd1 vccd1 vccd1 _4517_/B sky130_fd_sc_hd__inv_2
X_8284_ _8284_/A _8284_/B vssd1 vssd1 vccd1 vccd1 _8284_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5496_ _5435_/A _4933_/X _5436_/A _4930_/X _5495_/X vssd1 vssd1 vccd1 vccd1 _5496_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_110_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8130__B2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7235_ _7234_/Y _6941_/B _7249_/S vssd1 vssd1 vccd1 vccd1 _7236_/A sky130_fd_sc_hd__mux2_2
X_4447_ _4760_/A _4502_/A vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__nor2_1
XANTENNA__8681__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7660__A _7660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5495__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6692__A1 _5548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7166_ _5803_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7166_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_95_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4378_ hold40/X hold4/X vssd1 vssd1 vccd1 vccd1 _8917_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6117_ _8189_/A _6115_/Y _6116_/X vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__o21ai_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7096_/X _5367_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7098_/A sky130_fd_sc_hd__mux2_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7641__B1 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6048_ _6048_/A vssd1 vssd1 vccd1 vccd1 _6048_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6995__A2 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8491__A _8491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8197__B2 _8821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7944__A1 _7944_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7999_ _7989_/Y _7875_/X _7990_/Y _7874_/X _7998_/Y vssd1 vssd1 vccd1 vccd1 _7999_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__6747__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7944__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5955__B1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7835__A _7835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5183__A1 _5195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6380__B1 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5183__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8672__A2 _8515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7570__A _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8409__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5090__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4418__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6986__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6914__A _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8188__A1 _8192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7729__B _7729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6633__B _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6738__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5946__B1 _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4434__A _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5249__B _6181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output587_A _5138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7699__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7163__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6371__B1 _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6910__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5350_ _5337_/A _8271_/A _5338_/A _5191_/X _5349_/X vssd1 vssd1 vccd1 vccd1 _6622_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_2_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8112__A1 _8119_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8112__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4301_ _8971_/Q vssd1 vssd1 vccd1 vccd1 _6312_/A sky130_fd_sc_hd__buf_12
XFILLER_0_50_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5281_ _7829_/A _5333_/B _5280_/Y vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__o21ai_1
X_7020_ _7088_/A vssd1 vssd1 vccd1 vccd1 _7288_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__5477__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6674__B2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8971_ _8978_/CLK _8971_/D fanout732/X vssd1 vssd1 vccd1 vccd1 _8971_/Q sky130_fd_sc_hd__dfrtp_1
X_7922_ _7922_/A vssd1 vssd1 vccd1 vccd1 _7922_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7853_ _8166_/A _7859_/B vssd1 vssd1 vccd1 vccd1 _7853_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7639__B _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6543__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7926__A1 _7931_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6804_ _6804_/A vssd1 vssd1 vccd1 vccd1 _6804_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4344__A _5130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7784_ _7791_/A1 _5117_/A _7791_/B1 _5359_/B _7783_/X vssd1 vssd1 vccd1 vccd1 _7784_/X
+ sky130_fd_sc_hd__a221o_4
X_4996_ _4993_/X _7332_/B _6224_/S vssd1 vssd1 vccd1 vccd1 _4997_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5159__B _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6735_ _6729_/Y _6450_/X _6731_/X _6733_/Y _6734_/X vssd1 vssd1 vccd1 vccd1 _6735_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6666_ _6666_/A vssd1 vssd1 vccd1 vccd1 _6666_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7154__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7374__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5165__A1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8405_ _8403_/Y _8404_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8406_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5617_ _5617_/A _7431_/B vssd1 vssd1 vccd1 vccd1 _5617_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5165__B2 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6362__B1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6597_ _6924_/A _6597_/B vssd1 vssd1 vccd1 vccd1 _6597_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8189__C _8189_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8336_ _8334_/Y _8335_/Y _8336_/S vssd1 vssd1 vccd1 vccd1 _8337_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5548_ _5505_/A _4930_/X _5506_/A _4933_/X _5547_/X vssd1 vssd1 vccd1 vccd1 _5548_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_131_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8103__A1 _8106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8103__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8267_ _8267_/A vssd1 vssd1 vccd1 vccd1 _8267_/X sky130_fd_sc_hd__buf_1
X_5479_ _5764_/A1 _4871_/A input48/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5479_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5468__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6665__A1 _7470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7218_ _7668_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7218_/X sky130_fd_sc_hd__and2_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6665__B2 _5498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8198_ _8198_/A _8198_/B vssd1 vssd1 vccd1 vccd1 _8198_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7149_ _6727_/B _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7149_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7614__B1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7090__A1 _5094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7090__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7917__A1 _8352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7917__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7145__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5156__A1 _5195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5156__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8645__A2 _8012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5813__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5459__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6656__A1 _5465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6656__B2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6628__B _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5959__S _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6959__A2 _6261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7081__A1 _5328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__B1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7459__B _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7908__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5919__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4850_ _4850_/A _4850_/B hold19/A vssd1 vssd1 vccd1 vccd1 _8929_/B sky130_fd_sc_hd__nand3_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5395__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4781_ _4788_/A _8904_/A vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6592__B1 _5280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5395__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6520_ _5108_/B _6924_/A _6517_/Y _6518_/X _6519_/X vssd1 vssd1 vccd1 vccd1 _6520_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6451_ _6958_/B _4963_/X _6450_/X vssd1 vssd1 vccd1 vccd1 _6451_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__B _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5147__B2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6344__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5698__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5402_ _5402_/A vssd1 vssd1 vccd1 vccd1 _5402_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6382_ _5715_/B _6379_/Y _5128_/Y _6994_/C vssd1 vssd1 vccd1 vccd1 _6382_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8121_ _7777_/A _8515_/A _7792_/A vssd1 vssd1 vccd1 vccd1 _8121_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_140_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5333_ _6304_/A _5333_/B vssd1 vssd1 vccd1 vccd1 _5333_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5723__A _5723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6647__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7844__B1 hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8052_ _8045_/Y _7769_/A _8046_/Y _6500_/A _8051_/Y vssd1 vssd1 vccd1 vccd1 _8458_/A
+ sky130_fd_sc_hd__a221oi_4
X_5264_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5264_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7003_ _7384_/A _4408_/B _7769_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _7059_/A sky130_fd_sc_hd__a22o_4
XANTENNA__7634__A1_N _6867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5195_ _5195_/A1 _8271_/A _5195_/B1 _5191_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _5196_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7072__A1 _6566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8954_ _8967_/CLK _8954_/D fanout733/X vssd1 vssd1 vccd1 vccd1 _8954_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5083__B1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5622__A2 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7905_ _7905_/A1 _7876_/X _7905_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7905_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8885_ _8894_/C vssd1 vssd1 vccd1 vccd1 _8899_/A sky130_fd_sc_hd__inv_2
XFILLER_0_149_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7836_ _7836_/A _7836_/B vssd1 vssd1 vccd1 vccd1 _7836_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__8572__A1 _8244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4979_ _4977_/Y _4978_/Y _4674_/C vssd1 vssd1 vccd1 vccd1 _4979_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_19_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7767_ _7767_/A _8550_/B _7826_/A vssd1 vssd1 vccd1 vccd1 _7954_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6718_ _7524_/A _6549_/A _5620_/X _6876_/C vssd1 vssd1 vccd1 vccd1 _6718_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8324__A1 _7869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7127__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7698_ _7695_/X _7754_/A _7697_/Y vssd1 vssd1 vccd1 vccd1 _7698_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8324__B2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5138__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5617__B _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6335__B1 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6649_ _6644_/Y _6876_/C _6645_/Y _6647_/Y _6648_/Y vssd1 vssd1 vccd1 vccd1 _6649_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4897__B1 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8088__B1 _8093_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8319_ _7784_/X hold31/A _8759_/B vssd1 vssd1 vccd1 vccd1 _8319_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8627__A2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6729__A _6729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput580 _7757_/Y vssd1 vssd1 vccd1 vccd1 sports_o[170] sky130_fd_sc_hd__buf_12
Xoutput591 _5214_/X vssd1 vssd1 vccd1 vccd1 sports_o[180] sky130_fd_sc_hd__buf_12
XANTENNA__7063__A1 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8260__B1 _7771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6810__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8563__A1 _8230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8563__B2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5377__A1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5377__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6911__B _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5808__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7669__A3 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8079__B1 _8480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8618__A2 _7906_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output452_A _8489_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6629__A1 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5262__B _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5852__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8251__B1 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5604__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5951_ _6875_/B _5862_/A _5950_/Y vssd1 vssd1 vccd1 vccd1 _6854_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4902_ _5999_/B vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8670_ _8499_/A _8577_/X _8668_/X _8669_/X vssd1 vssd1 vccd1 vccd1 _8670_/X sky130_fd_sc_hd__a22o_1
X_5882_ _5804_/A _8271_/A _5805_/A _5191_/X _5881_/X vssd1 vssd1 vccd1 vccd1 _6801_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8554__A1 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7357__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5368__A1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4833_ _4833_/A _4833_/B vssd1 vssd1 vccd1 vccd1 _4833_/Y sky130_fd_sc_hd__nand2_1
X_7621_ _7620_/Y _7297_/B _7575_/A _7385_/Y vssd1 vssd1 vccd1 vccd1 _7621_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5368__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7552_ _5781_/A _7680_/B _7550_/X _7348_/A _7551_/X vssd1 vssd1 vccd1 vccd1 _7552_/X
+ sky130_fd_sc_hd__a221o_2
X_4764_ _4764_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _4768_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6503_ _6495_/X _6498_/Y _6502_/Y vssd1 vssd1 vccd1 vccd1 _6503_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7483_ _7673_/A _7483_/B vssd1 vssd1 vccd1 vccd1 _7483_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4695_ _4714_/A _4695_/B vssd1 vssd1 vccd1 vccd1 _4696_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6434_ _7384_/A _6434_/B vssd1 vssd1 vccd1 vccd1 _6435_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ _8444_/A _6369_/A1 _8257_/C input14/X vssd1 vssd1 vccd1 vccd1 _6365_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5540__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6549__A _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8104_ _8097_/Y _6500_/X _8098_/Y _7769_/X _8103_/Y vssd1 vssd1 vccd1 vccd1 _8104_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5316_ _6102_/B vssd1 vssd1 vccd1 vccd1 _6868_/B sky130_fd_sc_hd__buf_6
X_6296_ _6309_/A1 _8368_/A input71/X _4940_/A vssd1 vssd1 vccd1 vccd1 _6296_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput308 sports_i[48] vssd1 vssd1 vccd1 vccd1 _7976_/A sky130_fd_sc_hd__buf_1
X_8035_ _8028_/Y _5171_/B _8029_/Y _7304_/A _8034_/X vssd1 vssd1 vccd1 vccd1 _8444_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6096__A2 _6094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5247_ _5245_/X _5246_/X _6689_/S vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6983__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput319 sports_i[58] vssd1 vssd1 vccd1 vccd1 _8111_/A sky130_fd_sc_hd__buf_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5208_/A1 _4953_/X _5208_/B1 _4870_/A _5177_/X vssd1 vssd1 vccd1 vccd1 _6550_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__8483__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7045__A1 _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6284__A _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8242__B1 _4662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8793__A1 _8483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7596__A2 _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7099__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8937_ _8936_/A _4713_/B hold27/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8868_ _8868_/A _8868_/B vssd1 vssd1 vccd1 vccd1 _8971_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8545__A1 _8133_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7819_ _7817_/Y _7818_/Y _8845_/C vssd1 vssd1 vccd1 vccd1 _7819_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8799_ _8490_/A _8806_/B _8797_/X _8798_/X vssd1 vssd1 vccd1 vccd1 _8799_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5628__A _5628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6223__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6308__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7843__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5531__A1 _5587_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5531__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5363__A _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7808__B1 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6087__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8233__B1 _8232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8784__A1 _8445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5598__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6795__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4426__B _5827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7339__A2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8536__A1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8536__B2 _8137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7737__B _7737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6011__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4442__A hold10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5257__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5770__A1 _5722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8839__A2 _8252_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5770__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4480_ _6500_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4480_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6150_ _6174_/A1 _5090_/A input64/X _4874_/A vssd1 vssd1 vccd1 vccd1 _6150_/X sky130_fd_sc_hd__o22a_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6078__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5101_ _5136_/A vssd1 vssd1 vccd1 vccd1 _6402_/A sky130_fd_sc_hd__buf_6
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7275__A1 _7737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6122_/A _6080_/Y _6081_/S vssd1 vssd1 vccd1 vccd1 _6081_/X sky130_fd_sc_hd__mux2_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8472__B1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5032_ input84/X _8706_/B input21/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5825__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7578__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5589__A1 _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6983_ _6982_/X _7737_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6984_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4336__B _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8722_ _8824_/S vssd1 vssd1 vccd1 vccd1 _8782_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5934_ _5931_/Y _4885_/A _5932_/Y _4890_/A _5933_/Y vssd1 vssd1 vccd1 vccd1 _6852_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8527__A1 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8653_ _8439_/A _8577_/X _8651_/X _8652_/X vssd1 vssd1 vccd1 vccd1 _8653_/X sky130_fd_sc_hd__a22o_1
X_5865_ _5865_/A vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__inv_2
XFILLER_0_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7735__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4816_ _4816_/A _7511_/B vssd1 vssd1 vccd1 vccd1 _4817_/B sky130_fd_sc_hd__nand2_1
X_7604_ _7673_/A _7604_/B vssd1 vssd1 vccd1 vccd1 _7604_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4352__A hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8584_ _8584_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _8589_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_8_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5796_ _6761_/A _6689_/S vssd1 vssd1 vccd1 vccd1 _5796_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6978__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4747_ _4786_/B _8584_/B vssd1 vssd1 vccd1 vccd1 _4747_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5761__A1 _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7535_ _6727_/B _7348_/A _7531_/Y _7534_/Y vssd1 vssd1 vccd1 vccd1 _7535_/X sky130_fd_sc_hd__a2bb2o_2
XANTENNA__8759__A _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7466_ _7466_/A _7700_/B vssd1 vssd1 vccd1 vccd1 _7466_/X sky130_fd_sc_hd__and2_1
XFILLER_0_114_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4678_ _4713_/A vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__inv_2
XANTENNA__6305__A3 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6417_ _6434_/B _7309_/B vssd1 vssd1 vccd1 vccd1 _6925_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_102_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5513__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7397_ _6566_/B _7696_/B _7395_/X _7326_/A _7396_/Y vssd1 vssd1 vccd1 vccd1 _7397_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6348_ _6357_/A1 _8310_/B input75/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6348_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6069__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput105 mports_i[194] vssd1 vssd1 vccd1 vccd1 _5635_/A1 sky130_fd_sc_hd__buf_2
X_6279_ _6315_/B _8310_/B _6314_/B _5091_/X vssd1 vssd1 vccd1 vccd1 _6279_/X sky130_fd_sc_hd__o22a_1
Xinput116 mports_i[203] vssd1 vssd1 vccd1 vccd1 _5881_/A1 sky130_fd_sc_hd__buf_2
Xinput127 mports_i[213] vssd1 vssd1 vccd1 vccd1 _6140_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput138 mports_i[223] vssd1 vssd1 vccd1 vccd1 _4800_/B sky130_fd_sc_hd__buf_6
X_8018_ _8015_/Y _7013_/A _8016_/Y _5117_/A _8017_/Y vssd1 vssd1 vccd1 vccd1 _8433_/A
+ sky130_fd_sc_hd__a221oi_4
Xinput149 mports_i[28] vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8215__B1 _8222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7569__A2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6241__A2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7224__A_N _7678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8388__B _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7257__A1 _6277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7257__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8608__S _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5807__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7009__A1 _4876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7009__B2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6480__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8206__B1 _8210_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4437__A _4437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output415_A _8083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8757__A1 _7932_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6232__A2 _6944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8509__A1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7980__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5991__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5650_ _5622_/X _6402_/A _5633_/Y _5634_/X _5649_/X vssd1 vssd1 vccd1 vccd1 _5650_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7193__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7732__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _4601_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _8846_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5743__A1 _5764_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _6695_/B vssd1 vssd1 vccd1 vccd1 _5581_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5743__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7483__A _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7320_ _6440_/A _7347_/A _6456_/A _7349_/A vssd1 vssd1 vccd1 vccd1 _7320_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4532_ _4532_/A _4532_/B vssd1 vssd1 vccd1 vccd1 _4557_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_142_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7251_ _8919_/A _7251_/B vssd1 vssd1 vccd1 vccd1 _7251_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5715__B _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8693__B1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4463_ _5780_/A vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__inv_2
XANTENNA__7496__B2 _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6099__A _6180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6202_ _6202_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _6202_/Y sky130_fd_sc_hd__nand2_1
X_7182_ _7182_/A vssd1 vssd1 vccd1 vccd1 _7182_/X sky130_fd_sc_hd__buf_1
XFILLER_0_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4394_ _4394_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7248__A1 _6261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6133_ _6133_/A _6133_/B vssd1 vssd1 vccd1 vccd1 _6133_/Y sky130_fd_sc_hd__nand2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6827__A _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7799__A2 _7803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6892_/B _6211_/B vssd1 vssd1 vccd1 vccd1 _6064_/Y sky130_fd_sc_hd__nand2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5015_ input83/X _5090_/A input20/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5015_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6471__A2 _4899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5877__S _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _6303_/Y _6475_/A _6965_/Y _6694_/B _6994_/B vssd1 vssd1 vccd1 vccd1 _6966_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5431__B1 _5386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7971__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8705_ _8244_/X _8686_/B _8703_/X _8704_/X vssd1 vssd1 vccd1 vccd1 _8705_/X sky130_fd_sc_hd__a22o_1
X_5917_ _5715_/B _5907_/X _5909_/Y _5916_/X vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__a31o_2
XFILLER_0_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6897_ _6897_/A vssd1 vssd1 vccd1 vccd1 _6897_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8636_ _8636_/A vssd1 vssd1 vccd1 vccd1 _8636_/X sky130_fd_sc_hd__buf_1
XFILLER_0_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7184__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5848_ _5772_/X _7316_/A _8194_/A _5824_/X vssd1 vssd1 vccd1 vccd1 _5849_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5734__A1 _7551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8567_ _8567_/A _8567_/B vssd1 vssd1 vccd1 vccd1 _8567_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5734__B2 _6758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5779_ _5159_/B _5744_/X _5766_/X _6402_/A _5778_/X vssd1 vssd1 vccd1 vccd1 _5779_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7518_ _7510_/B _5679_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7520_/B sky130_fd_sc_hd__o21ai_1
X_8498_ _8498_/A vssd1 vssd1 vccd1 vccd1 _8498_/X sky130_fd_sc_hd__buf_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8684__B1 _8190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7487__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7449_ _7606_/A _7449_/B vssd1 vssd1 vccd1 vccd1 _7449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5498__B1 _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7239__A1 _7705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8428__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6737__A _6737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6456__B _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7568__A _7686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6214__A2 _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5973__A1 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7175__A0 _7174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8911__A1 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7714__A2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5725__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7478__A1 _5496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput409 _8014_/X vssd1 vssd1 vccd1 vccd1 mports_o[16] sky130_fd_sc_hd__buf_12
XFILLER_0_120_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6150__A1 _6174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6150__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8958__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6205__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6820_ _6820_/A vssd1 vssd1 vccd1 vccd1 _6820_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_147_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5413__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7953__A2 _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6751_ _6751_/A _6899_/B vssd1 vssd1 vccd1 vccd1 _6751_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5702_ _5702_/A _6689_/S vssd1 vssd1 vccd1 vccd1 _5702_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6682_ _5498_/X _7536_/B _7707_/B _5544_/X vssd1 vssd1 vccd1 vccd1 _7476_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7166__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8902__A1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8421_ _8564_/B _8012_/Y _8497_/S vssd1 vssd1 vccd1 vccd1 _8421_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5716__A1 _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5633_ _6720_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _5633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5716__B2 _5715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5726__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5564_ _5591_/A _5102_/A _5592_/A _5191_/X _5563_/X vssd1 vssd1 vccd1 vccd1 _5634_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__4630__A _4760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8352_ _8352_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8352_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4515_ _4515_/A _4515_/B vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__nand2_1
X_7303_ _7630_/B vssd1 vssd1 vccd1 vccd1 _7532_/A sky130_fd_sc_hd__inv_2
XFILLER_0_130_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8666__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8283_ _8283_/A vssd1 vssd1 vccd1 vccd1 _8283_/X sky130_fd_sc_hd__buf_1
X_5495_ _5497_/A1 _8706_/B input38/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5495_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8130__A2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6141__A1 _6141_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4446_ _4446_/A _4446_/B vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__nand2_1
X_7234_ _7234_/A vssd1 vssd1 vccd1 vccd1 _7234_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7660__B _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7165_ _7165_/A vssd1 vssd1 vccd1 vccd1 _7165_/X sky130_fd_sc_hd__buf_1
XANTENNA__6692__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4377_ _4392_/A _5485_/A vssd1 vssd1 vccd1 vccd1 _4377_/X sky130_fd_sc_hd__and2_1
X_6116_ _6281_/S _6116_/B vssd1 vssd1 vccd1 vccd1 _6116_/X sky130_fd_sc_hd__or2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _6622_/A _7023_/X _7095_/X vssd1 vssd1 vccd1 vccd1 _7096_/X sky130_fd_sc_hd__o21a_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6047_/A vssd1 vssd1 vccd1 vccd1 _6047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6991__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7641__A1 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8491__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ _7998_/A1 _7876_/X _7998_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7998_/Y sky130_fd_sc_hd__o22ai_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7944__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5955__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6949_ _7705_/B _6908_/B _6947_/B _6940_/Y vssd1 vssd1 vccd1 vccd1 _6949_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8619_ _8346_/A _8577_/X _8617_/X _8618_/X vssd1 vssd1 vccd1 vccd1 _8619_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_64_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6380__A1 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5183__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6380__B2 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5355__B _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8121__A2 _8515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7851__A _7851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6132__A1 _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6132__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7880__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7298__A _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5946__A1 _5931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4434__B hold10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5946__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8621__S _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7699__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8896__B1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6371__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8954__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8112__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7761__A _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4300_ _4300_/A _4389_/A vssd1 vssd1 vccd1 vccd1 _4300_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6123__A1 _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5280_ _5280_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5280_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6674__A2 _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7871__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5882__B1 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8970_ _8978_/CLK _8970_/D fanout732/X vssd1 vssd1 vccd1 vccd1 _8970_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7921_ _7760_/X _7912_/Y _7917_/X _7920_/X vssd1 vssd1 vccd1 vccd1 _7921_/X sky130_fd_sc_hd__a22o_2
XANTENNA__4988__A2 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7852_ _7852_/A _7858_/B vssd1 vssd1 vccd1 vccd1 _7852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7926__A2 _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6803_ _6906_/A _5891_/A _6802_/Y vssd1 vssd1 vccd1 vccd1 _6804_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7783_ _7761_/A _7790_/A2 _7316_/A _7790_/B2 vssd1 vssd1 vccd1 vccd1 _7783_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4344__B _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4995_ _4975_/A _4930_/X _4976_/A _4933_/X _4994_/X vssd1 vssd1 vccd1 vccd1 _7332_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_86_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6734_ _6743_/A _6510_/A _5657_/X _6512_/X vssd1 vssd1 vccd1 vccd1 _6734_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6665_ _7470_/A _7311_/A _8151_/B _5498_/X vssd1 vssd1 vccd1 vccd1 _6666_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8404_ _8404_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8404_/Y sky130_fd_sc_hd__nand2_1
X_5616_ _5616_/A vssd1 vssd1 vccd1 vccd1 _7431_/B sky130_fd_sc_hd__buf_8
XANTENNA__5165__A2 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6362__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6596_ _6592_/X _6933_/A _6968_/A _6595_/X vssd1 vssd1 vccd1 vccd1 _6596_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8335_ _8335_/A _8335_/B vssd1 vssd1 vccd1 vccd1 _8335_/Y sky130_fd_sc_hd__nand2_1
X_5547_ _5557_/A1 _8706_/B input40/X _4940_/X vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_42_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8103__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6114__A1 _6141_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6114__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5478_ _5685_/A _5089_/A _5686_/A _4868_/A _5477_/X vssd1 vssd1 vccd1 vccd1 _5738_/C
+ sky130_fd_sc_hd__o221a_4
X_8266_ _8262_/X _8263_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8267_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7217_ _7217_/A vssd1 vssd1 vccd1 vccd1 _7217_/X sky130_fd_sc_hd__buf_1
XANTENNA__6665__A2 _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4429_ _4453_/A _8709_/A vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8197_ _8184_/X _8191_/Y _7760_/X _8821_/A vssd1 vssd1 vccd1 vccd1 _8197_/X sky130_fd_sc_hd__a2bb2o_2
XANTENNA__5191__A _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5873__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7148_ _7148_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7148_/X sky130_fd_sc_hd__and2_1
XANTENNA__7075__C1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7614__A1 _6841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7079_ _7413_/A _7059_/X _5280_/A _7246_/B _7061_/X vssd1 vssd1 vccd1 vccd1 _7079_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7090__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7917__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__A1 _5928_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8327__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7057__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5156__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6353__A1 _6349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6353__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7581__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6105__A1 _6047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6105__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6656__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5813__B _7171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4429__B _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7066__C1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7605__A1 _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5092__A1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5092__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7908__A2 _8346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5919__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5975__S _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7756__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4780_ _4747_/Y _4802_/A _4803_/A vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__B2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6450_ _6450_/A vssd1 vssd1 vccd1 vccd1 _6450_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5147__A2 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6344__A1 _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5401_ _5401_/A vssd1 vssd1 vccd1 vccd1 _5401_/Y sky130_fd_sc_hd__inv_2
X_6381_ _6388_/A1 _8444_/A input15/X _8257_/C _6380_/X vssd1 vssd1 vccd1 vccd1 _6994_/C
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6895__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8587__A _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8120_ _8110_/Y _7874_/A _8111_/Y _8174_/A _8119_/Y vssd1 vssd1 vccd1 vccd1 _8515_/A
+ sky130_fd_sc_hd__a221oi_4
X_5332_ _5312_/X _6402_/A _5322_/Y _5324_/Y _5331_/X vssd1 vssd1 vccd1 vccd1 _5332_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5263_ _6593_/A _5253_/X _5262_/Y vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__o21ai_1
X_8051_ _8054_/A1 _5780_/X _8054_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _8051_/Y sky130_fd_sc_hd__o22ai_2
X_7002_ _7002_/A vssd1 vssd1 vccd1 vccd1 _7002_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5194_ input88/X _5192_/X input26/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_76_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7072__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8953_ _8979_/CLK _8953_/D fanout732/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__5083__A1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5083__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7904_ _7901_/Y _7768_/X _7903_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7904_/X
+ sky130_fd_sc_hd__a221o_1
X_8884_ _8884_/A _8884_/B vssd1 vssd1 vccd1 vccd1 _8972_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8021__A1 _8024_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7835_ _7835_/A vssd1 vssd1 vccd1 vccd1 _7836_/B sky130_fd_sc_hd__buf_8
XANTENNA__8021__B2 _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7766_ _8709_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _7826_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_136_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4978_ hold26/A _4978_/B vssd1 vssd1 vccd1 vccd1 _4978_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7780__B1 _4481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6717_ _6724_/A _5617_/A _5600_/Y _6475_/X vssd1 vssd1 vccd1 vccd1 _6717_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7697_ _7673_/A _6211_/A _7696_/Y vssd1 vssd1 vccd1 vccd1 _7697_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8324__A2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5138__A2 _7352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6648_ _6841_/A _6648_/B vssd1 vssd1 vccd1 vccd1 _6648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6579_ _7394_/B _6912_/B _6575_/X _6577_/Y _6578_/Y vssd1 vssd1 vccd1 vccd1 _6580_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4897__A1 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4897__B2 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8088__A1 _8093_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8318_ _8314_/X _8317_/X _8496_/S vssd1 vssd1 vccd1 vccd1 _8318_/X sky130_fd_sc_hd__mux2_1
XANTENNA__8088__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6729__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5633__B _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6638__A2 _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8249_ _8251_/B2 _8163_/A _8252_/B1 _5171_/B _8248_/X vssd1 vssd1 vccd1 vccd1 _8249_/X
+ sky130_fd_sc_hd__a221o_4
Xoutput570 _7717_/X vssd1 vssd1 vccd1 vccd1 sports_o[161] sky130_fd_sc_hd__buf_12
Xoutput581 _4952_/X vssd1 vssd1 vccd1 vccd1 sports_o[171] sky130_fd_sc_hd__buf_12
XANTENNA__5846__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput592 _5234_/X vssd1 vssd1 vccd1 vccd1 sports_o[181] sky130_fd_sc_hd__buf_12
XANTENNA__4964__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8260__A1 _7765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7063__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8260__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6271__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8012__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8563__A2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6574__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4585__B1 _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5096__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6326__A1 _6326_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6326__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6877__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8079__A1 _8483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8079__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output445_A _8411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8251__A1 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7054__A2 _5150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8251__B2 _8251_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6262__B1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5950_ _6001_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _5950_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4901_ _6312_/A _7302_/B vssd1 vssd1 vccd1 vccd1 _5999_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5881_ _5881_/A1 _5192_/X input52/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_29_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7620_ _7620_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7620_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4832_ _8952_/D hold7/X vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5368__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7762__B1 _7779_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7551_ _7551_/A _7660_/B vssd1 vssd1 vccd1 vccd1 _7551_/X sky130_fd_sc_hd__and2_1
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4763_ _4763_/A vssd1 vssd1 vccd1 vccd1 _4764_/B sky130_fd_sc_hd__inv_2
XFILLER_0_56_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6502_ _6543_/A _6841_/A _6501_/X vssd1 vssd1 vccd1 vccd1 _6502_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6317__A1 _6326_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6317__B2 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7482_ _7348_/A _7480_/X _7481_/X vssd1 vssd1 vccd1 vccd1 _7482_/X sky130_fd_sc_hd__a21o_1
X_4694_ _4694_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4695_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6433_ _6456_/A _6488_/B _6432_/X vssd1 vssd1 vccd1 vccd1 _6433_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6364_ _6369_/A1 _8516_/B input14/X _4913_/X _6363_/X vssd1 vssd1 vccd1 vccd1 _6364_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5540__A2 _7120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8103_ _8106_/A1 _5780_/X _8106_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _8103_/Y sky130_fd_sc_hd__o22ai_2
X_5315_ _5294_/A _8271_/A _5295_/A _5191_/X _5314_/X vssd1 vssd1 vccd1 vccd1 _5317_/A
+ sky130_fd_sc_hd__o221a_4
X_6295_ input10/X _4933_/A _6337_/B1 _8523_/B _6294_/X vssd1 vssd1 vccd1 vccd1 _7733_/B
+ sky130_fd_sc_hd__o221a_2
XANTENNA__7293__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8034_ _6024_/A _8030_/Y _6411_/A _8031_/Y vssd1 vssd1 vccd1 vccd1 _8034_/X sky130_fd_sc_hd__a22o_1
X_5246_ _6566_/B _5197_/X _7707_/B _5248_/A vssd1 vssd1 vccd1 vccd1 _5246_/X sky130_fd_sc_hd__a22o_1
Xinput309 sports_i[49] vssd1 vssd1 vccd1 vccd1 _7989_/A sky130_fd_sc_hd__clkbuf_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ input90/X _5090_/A input27/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7160__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7045__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8242__B2 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8936_ _8936_/A hold26/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8867_ _5359_/B _8857_/A _6264_/X _4591_/A vssd1 vssd1 vccd1 vccd1 _8868_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_66_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7396__A _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7818_ _7818_/A _8842_/B vssd1 vssd1 vccd1 vccd1 _7818_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8798_ _8833_/B _8516_/A _8725_/A vssd1 vssd1 vccd1 vccd1 _8798_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6556__B2 _6511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5628__B _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7749_ _7748_/X _6385_/Y _7749_/S vssd1 vssd1 vccd1 vccd1 _7749_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6308__A1 _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7843__B _7859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5644__A _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5531__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7808__A1 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7284__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6492__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6475__A _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8233__A1 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8233__B2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5598__A2 _5637_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8536__A2 _8821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7744__B1 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output395_A _8807_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5770__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7753__B _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4730__B1 _4760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _6233_/B _5076_/X _5095_/Y _6133_/B _5099_/X vssd1 vssd1 vccd1 vccd1 _5100_/X
+ sky130_fd_sc_hd__a221o_1
X_6080_ _6080_/A _6897_/A vssd1 vssd1 vccd1 vccd1 _6080_/Y sky130_fd_sc_hd__nor2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8584__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__A1 _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5031_ _6224_/S vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__clkbuf_8
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8224__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5038__A1 _5070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5038__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6235__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8775__A2 _7999_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6982_ _4793_/A _6467_/X _6981_/X vssd1 vssd1 vccd1 vccd1 _6982_/X sky130_fd_sc_hd__o21a_1
X_8721_ _8309_/X _8803_/B _8313_/X _8711_/X _8820_/B vssd1 vssd1 vccd1 vccd1 _8721_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5933_ _5274_/A _6007_/A1 _5275_/A input57/X vssd1 vssd1 vccd1 vccd1 _5933_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8527__A2 _8133_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8652_ _8698_/B _8042_/Y _8590_/X vssd1 vssd1 vccd1 vccd1 _8652_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5864_ _5864_/A vssd1 vssd1 vccd1 vccd1 _5864_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7735__B1 _6980_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7603_ _7348_/A _5860_/A _7334_/A vssd1 vssd1 vccd1 vccd1 _7603_/X sky130_fd_sc_hd__o21a_1
X_4815_ _4607_/A _4748_/B _4583_/Y _4814_/B vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8583_ _8583_/A vssd1 vssd1 vccd1 vccd1 _8583_/X sky130_fd_sc_hd__buf_4
XFILLER_0_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5795_ _5795_/A vssd1 vssd1 vccd1 vccd1 _6761_/A sky130_fd_sc_hd__inv_2
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7534_ _7532_/Y _7533_/Y _7497_/B vssd1 vssd1 vccd1 vccd1 _7534_/Y sky130_fd_sc_hd__o21ai_1
X_4746_ _4814_/B _4818_/B vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_145_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8759__B _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7465_ _7701_/A _5464_/X _7683_/C vssd1 vssd1 vccd1 vccd1 _7466_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4677_ _4677_/A _4677_/B vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6416_ _4876_/X _6994_/B _4899_/Y _6989_/B vssd1 vssd1 vccd1 vccd1 _6416_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5513__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6710__A1 _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7396_ _7673_/A _7396_/B vssd1 vssd1 vccd1 vccd1 _7396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6710__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6347_ _7737_/B _5031_/X _6346_/X vssd1 vssd1 vccd1 vccd1 _6347_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8463__A1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6278_ _7769_/A _6278_/B vssd1 vssd1 vccd1 vccd1 _6278_/Y sky130_fd_sc_hd__nor2_1
Xinput106 mports_i[195] vssd1 vssd1 vccd1 vccd1 _5640_/A1 sky130_fd_sc_hd__buf_2
Xinput117 mports_i[204] vssd1 vssd1 vccd1 vccd1 _5902_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__5277__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput128 mports_i[214] vssd1 vssd1 vccd1 vccd1 _6174_/A1 sky130_fd_sc_hd__buf_2
X_8017_ _8024_/A1 _4947_/B _8024_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _8017_/Y sky130_fd_sc_hd__o22ai_2
Xinput139 mports_i[224] vssd1 vssd1 vccd1 vccd1 _6357_/A1 sky130_fd_sc_hd__clkbuf_4
X_5229_ _5229_/A vssd1 vssd1 vccd1 vccd1 _7874_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__8215__A1 _4312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8215__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5029__A1 _5028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8919_ _8919_/A hold10/X vssd1 vssd1 vccd1 vccd1 _8922_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5639__A _5655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4543__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5201__A1 _6181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5201__B2 _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8685__A _8820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7257__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5268__B2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7009__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8206__A1 _8210_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8206__B2 _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8979__RESET_B input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6933__A _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output408_A _8001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6768__A1 _5770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6768__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5549__A _5549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6144__S _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5991__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7193__A1 _6841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600_ _4600_/A _4600_/B vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5743__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5580_ _5610_/A _5509_/Y _6081_/S vssd1 vssd1 vccd1 vccd1 _5580_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_14_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8579__B _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ _4531_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _4532_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5284__A _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7250_ _7250_/A vssd1 vssd1 vccd1 vccd1 _7250_/X sky130_fd_sc_hd__buf_1
XANTENNA__7496__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4462_ _8166_/A hold23/A vssd1 vssd1 vccd1 vccd1 _5780_/A sky130_fd_sc_hd__nand2_8
XANTENNA__6099__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6201_ _5845_/B _7686_/B _6133_/B _7694_/B _6200_/X vssd1 vssd1 vccd1 vccd1 _6202_/A
+ sky130_fd_sc_hd__a221o_1
X_7181_ _7179_/X _5853_/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7182_/A sky130_fd_sc_hd__mux2_1
X_4393_ _4393_/A _4393_/B vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6132_ _5013_/Y _6131_/Y _6081_/X _5997_/B vssd1 vssd1 vccd1 vccd1 _6132_/X sky130_fd_sc_hd__a22o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7248__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6827__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5259__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6063_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6892_/B sky130_fd_sc_hd__nand2_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7004__A _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5014_ _5011_/Y _5012_/Y _5013_/Y vssd1 vssd1 vccd1 vccd1 _5014_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4347__B _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6843__A _6843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6562__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6965_ _6965_/A _6965_/B vssd1 vssd1 vccd1 vccd1 _6965_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5431__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5431__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8704_ _8698_/B _8252_/X _8590_/A vssd1 vssd1 vccd1 vccd1 _8704_/X sky130_fd_sc_hd__o21a_1
X_5916_ _6084_/B _5857_/Y _5915_/Y _5096_/A vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6054__S _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7708__B1 _7242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6896_ _6095_/A _6429_/S _6895_/X vssd1 vssd1 vccd1 vccd1 _6896_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8635_ _8634_/X _8375_/A _8690_/S vssd1 vssd1 vccd1 vccd1 _8636_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7184__A1 _6811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5847_ _6128_/B _6788_/B _5136_/A vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_146_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8566_ _8239_/Y _8304_/A _8240_/Y _8299_/A vssd1 vssd1 vccd1 vccd1 _8567_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5778_ _5778_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__and2_1
XANTENNA__5734__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7517_ _7509_/Y _7536_/A _7513_/X _7516_/Y vssd1 vssd1 vccd1 vccd1 _7517_/X sky130_fd_sc_hd__a22o_1
X_4729_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__inv_2
X_8497_ _8494_/Y _8496_/X _8497_/S vssd1 vssd1 vccd1 vccd1 _8498_/A sky130_fd_sc_hd__mux2_2
XANTENNA__4810__B _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8684__A1 _8187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7487__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7448_ _7701_/A _6630_/A _6264_/X vssd1 vssd1 vccd1 vccd1 _7449_/B sky130_fd_sc_hd__o21a_1
XANTENNA__8684__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5498__A1 _5435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5498__B2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7379_ _7378_/X _5211_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7379_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8436__A1 _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8739__A2 _7856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5973__A2 _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7175__A1 _5824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5725__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6922__A1 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6922__B2 _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5816__B _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4720__B _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8675__A1 _8133_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5489__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5489__B2 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6150__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5832__A _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7402__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5413__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6610__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6750_ _5745_/Y _6475_/A _5713_/Y _6694_/B vssd1 vssd1 vccd1 vccd1 _6751_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_147_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5701_ _6732_/A _5197_/X _8151_/B _7544_/A vssd1 vssd1 vccd1 vccd1 _5701_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6681_ _6681_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7166__A1 _5803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8363__B1 _8362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8420_ _8009_/Y _8299_/X _8419_/X _8304_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8420_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5177__B1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4911__A _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5632_ _6870_/S _5566_/B _5631_/Y vssd1 vssd1 vccd1 vccd1 _6720_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5716__A2 _6732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8351_ _8351_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8351_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5726__B _6756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5563_ _5635_/A1 _5192_/X input42/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5563_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8115__B1 _8111_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7302_ _7510_/B _7302_/B vssd1 vssd1 vccd1 vccd1 _7630_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8666__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4514_ _4514_/A _4525_/B _4525_/C vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__nand3_1
XANTENNA__7469__A2 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8282_ _8281_/Y _7796_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8283_/A sky130_fd_sc_hd__mux2_1
X_5494_ _5031_/X _5464_/X _5490_/Y _5493_/X vssd1 vssd1 vccd1 vccd1 _5494_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_130_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7233_ _7696_/A _7138_/A _7232_/X vssd1 vssd1 vccd1 vccd1 _7234_/A sky130_fd_sc_hd__o21ai_2
X_4445_ _4454_/B _8189_/B _4453_/A vssd1 vssd1 vccd1 vccd1 _4446_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7164_ _7163_/X _5770_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7165_/A sky130_fd_sc_hd__mux2_1
X_4376_ _5827_/B _4591_/B vssd1 vssd1 vccd1 vccd1 _4392_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6557__B _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6115_ _6115_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6115_/Y sky130_fd_sc_hd__nand2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _5400_/A _7004_/X _7094_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7095_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6046_/A vssd1 vssd1 vccd1 vccd1 _7639_/A sky130_fd_sc_hd__inv_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7641__A2 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8772__B _8772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5652__A1 _5697_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5652__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6573__A _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _8403_/A _7954_/X _8424_/A _7826_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7997_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5404__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _6948_/A _8857_/B vssd1 vssd1 vccd1 vccd1 _6948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_138_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5955__A2 _5899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6879_ _6016_/A _6841_/A _6876_/Y _6878_/X vssd1 vssd1 vccd1 vccd1 _6879_/X sky130_fd_sc_hd__o211a_2
XFILLER_0_153_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5168__B1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8618_ _8698_/B _7906_/Y _8590_/X vssd1 vssd1 vccd1 vccd1 _8618_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6904__A1 _6094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8549_ _4874_/X _8169_/Y _4870_/X _8206_/X _8548_/X vssd1 vssd1 vccd1 vccd1 _8549_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6380__A2 _6387_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8409__A1 _8424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8409__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7880__A2 _7867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6840__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8593__B1 _7788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5946__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5827__A _5827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6422__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8896__A1 _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7699__A2 _6941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8648__A1 _8782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8857__B _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6658__A _7470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6123__A2 _7678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7320__A1 _6440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7320__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7871__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5882__A1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5882__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7084__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7920_ _7777_/X _8335_/A _7792_/X vssd1 vssd1 vccd1 vccd1 _7920_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7851_ _7851_/A vssd1 vssd1 vccd1 vccd1 _7851_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4625__B _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6802_ _6802_/A _6906_/A vssd1 vssd1 vccd1 vccd1 _6802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5398__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7782_ _7760_/X _7763_/X _7775_/X _7781_/X vssd1 vssd1 vccd1 vccd1 _7782_/X sky130_fd_sc_hd__a22o_2
X_4994_ _4978_/B _8706_/B _4977_/B _4940_/X vssd1 vssd1 vccd1 vccd1 _4994_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6733_ _6733_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6733_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6664_ _5464_/X _6429_/S _6657_/X _6663_/X vssd1 vssd1 vccd1 vccd1 _6664_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8403_ _8403_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8403_/Y sky130_fd_sc_hd__nand2_1
X_5615_ _7304_/A vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6362__A2 _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6595_ _6854_/A _6594_/Y _7413_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6595_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_121_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8334_ _8334_/A _8335_/B vssd1 vssd1 vccd1 vccd1 _8334_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8639__A1 _8390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5546_ _5031_/X _5530_/X _5542_/X _5545_/X vssd1 vssd1 vccd1 vccd1 _5546_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8265_ _8497_/S vssd1 vssd1 vccd1 vccd1 _8572_/S sky130_fd_sc_hd__inv_6
XANTENNA__6114__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5477_ _5718_/A1 _4871_/A input47/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5477_/X sky130_fd_sc_hd__o22a_1
X_7216_ _7215_/X _6094_/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7217_/A sky130_fd_sc_hd__mux2_2
X_4428_ _4526_/A _4526_/B _4591_/B vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__nand3_2
X_8196_ _8189_/C _7761_/A _8196_/B1 _8857_/B _8195_/X vssd1 vssd1 vccd1 vccd1 _8821_/A
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5873__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7147_ _7147_/A vssd1 vssd1 vccd1 vccd1 _7147_/X sky130_fd_sc_hd__buf_1
X_4359_ _4716_/B vssd1 vssd1 vccd1 vccd1 _4360_/B sky130_fd_sc_hd__inv_2
XANTENNA__7614__A2 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7078_ _7078_/A vssd1 vssd1 vccd1 vccd1 _7078_/X sky130_fd_sc_hd__buf_1
X_6029_ _6284_/A _6029_/B vssd1 vssd1 vccd1 vccd1 _6029_/Y sky130_fd_sc_hd__nor2_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6050__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8327__B1 _7890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5647__A _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8948__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6353__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7862__A _7862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7550__B2 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6105__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7073__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7066__B1 _7383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8802__A1 _8499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7605__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6925__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7102__A _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4445__B _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8566__B1 _8240_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7369__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6941__A _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5919__A2 _6828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7756__B _7756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output592_A _5234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6344__A2 _7737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7541__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5400_ _5400_/A vssd1 vssd1 vccd1 vccd1 _7439_/B sky130_fd_sc_hd__inv_2
XFILLER_0_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6380_ _8713_/C _6387_/A1 _8579_/C input77/X vssd1 vssd1 vccd1 vccd1 _6380_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_152_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5331_ _5159_/B _5328_/A _5330_/Y _5125_/X vssd1 vssd1 vccd1 vccd1 _5331_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8050_ _8045_/Y _6079_/A _8046_/Y _6513_/A _8049_/Y vssd1 vssd1 vccd1 vccd1 _8455_/A
+ sky130_fd_sc_hd__a221oi_4
X_5262_ _5262_/A _6593_/A vssd1 vssd1 vccd1 vccd1 _5262_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6501__C1 _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7001_ _7000_/X _7756_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _7002_/A sky130_fd_sc_hd__mux2_1
X_5193_ _5193_/A vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__7057__A0 _7056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6835__B _6940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6327__S _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4843__A2_N _8976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8952_ _8979_/CLK _8952_/D fanout732/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__5083__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6280__A1 _6326_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6280__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7903_ _7896_/Y _7769_/X _7897_/Y _6500_/X _7902_/Y vssd1 vssd1 vccd1 vccd1 _7903_/Y
+ sky130_fd_sc_hd__a221oi_4
X_8883_ _4824_/B _8882_/Y _4818_/A vssd1 vssd1 vccd1 vccd1 _8884_/B sky130_fd_sc_hd__a21o_1
XANTENNA__6518__A1_N _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7834_ _7823_/A _4474_/A _8181_/A vssd1 vssd1 vccd1 vccd1 _7834_/X sky130_fd_sc_hd__mux2_1
XANTENNA__8021__A2 _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6032__A1 _5965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6032__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7765_ _4318_/B _5171_/B _4481_/B _5299_/B _7764_/X vssd1 vssd1 vccd1 vccd1 _7765_/X
+ sky130_fd_sc_hd__a221o_4
X_4977_ _8512_/S _4977_/B vssd1 vssd1 vccd1 vccd1 _4977_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8309__B1 _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7780__A1 _4318_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7780__B2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6716_ _5679_/A _6908_/B _5651_/X _6512_/X _6715_/X vssd1 vssd1 vccd1 vccd1 _6716_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__5791__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7696_ _7696_/A _7696_/B vssd1 vssd1 vccd1 vccd1 _7696_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6997__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6647_ _6432_/X _6646_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6647_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6335__A2 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6578_ _6841_/A _6578_/B vssd1 vssd1 vccd1 vccd1 _6578_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4897__A2 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5914__B _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8317_ _4913_/X _8315_/Y _8336_/S _8284_/Y _8316_/Y vssd1 vssd1 vccd1 vccd1 _8317_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_42_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5529_ _5543_/A1 _8706_/B input39/X _4940_/X vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8088__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5406__S _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8248_ _6965_/A _8251_/A2 _5299_/B _8252_/A1 vssd1 vssd1 vccd1 vccd1 _8248_/X sky130_fd_sc_hd__a22o_1
Xoutput560 _7647_/X vssd1 vssd1 vccd1 vccd1 sports_o[152] sky130_fd_sc_hd__buf_12
Xoutput571 _7721_/Y vssd1 vssd1 vccd1 vccd1 sports_o[162] sky130_fd_sc_hd__buf_12
Xoutput582 _4968_/X vssd1 vssd1 vccd1 vccd1 sports_o[172] sky130_fd_sc_hd__buf_12
Xoutput593 _5290_/X vssd1 vssd1 vccd1 vccd1 sports_o[182] sky130_fd_sc_hd__buf_12
X_8179_ _8179_/A vssd1 vssd1 vccd1 vccd1 _8179_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8260__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6271__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6271__B2 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8452__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8012__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6023__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7068__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7771__A1 _7779_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7771__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4585__A1 _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4585__B2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4712__C _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6326__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7523__B2 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8079__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7287__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5837__A1 _5881_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5837__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5051__S _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6262__A1 _6262_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6262__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8539__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7767__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4900_ hold40/A vssd1 vssd1 vccd1 vccd1 _7302_/B sky130_fd_sc_hd__inv_4
XFILLER_0_48_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6671__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5880_ _5096_/A _5864_/Y _5878_/X _5715_/B _5879_/X vssd1 vssd1 vccd1 vccd1 _5880_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6014__A1 _6061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6014__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4831_ _4850_/B hold19/X vssd1 vssd1 vccd1 vccd1 _8952_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4903__B _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7762__B2 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7550_ _5745_/Y _7630_/B _5727_/Y _8755_/C vssd1 vssd1 vccd1 vccd1 _7550_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_117_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4762_ _4762_/A _4762_/B vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5773__B1 _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6501_ _6500_/X _6543_/A _5062_/D _5185_/A _6854_/A vssd1 vssd1 vccd1 vccd1 _6501_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7481_ _6679_/B _7660_/B _5502_/X _7363_/A vssd1 vssd1 vccd1 vccd1 _7481_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6317__A2 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4693_ _4693_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4713_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6432_ _6432_/A vssd1 vssd1 vccd1 vccd1 _6432_/X sky130_fd_sc_hd__buf_6
XFILLER_0_153_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6363_ _6368_/A1 _8716_/B input76/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6363_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8102_ _8097_/Y _6513_/A _8098_/Y _6080_/A _8101_/Y vssd1 vssd1 vccd1 vccd1 _8503_/A
+ sky130_fd_sc_hd__a221oi_4
X_5314_ input95/X _5192_/X input32/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5314_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_3_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6294_ _6336_/A1 _8368_/A input73/X _4940_/A vssd1 vssd1 vccd1 vccd1 _6294_/X sky130_fd_sc_hd__o22a_1
X_8033_ _8028_/Y _5359_/B _8029_/Y _5237_/A _8032_/X vssd1 vssd1 vccd1 vccd1 _8439_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5245_ _5323_/A _7536_/B _7707_/B _5356_/B vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__a22o_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _5176_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _5176_/Y sky130_fd_sc_hd__nand2_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6565__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8935_ hold11/X _8935_/B vssd1 vssd1 vccd1 vccd1 _8961_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8866_ _8865_/Y _4591_/A _7372_/B vssd1 vssd1 vccd1 vccd1 _8868_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7202__B1 _7201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5909__B _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7817_ _7829_/B _8194_/A vssd1 vssd1 vccd1 vccd1 _7817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8797_ _8511_/A _8803_/B _8091_/Y _8711_/X _8788_/S vssd1 vssd1 vccd1 vccd1 _8797_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5197__A _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7748_ _7640_/B _6379_/Y _7349_/Y _6994_/C vssd1 vssd1 vccd1 vccd1 _7748_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5764__B1 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6308__A2 _7725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7679_ _6115_/A _7686_/A _7347_/A _7678_/Y _7334_/A vssd1 vssd1 vccd1 vccd1 _7679_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8702__B1 _4662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7808__A2 _7813_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5819__A1 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6756__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput390 _8789_/X vssd1 vssd1 vccd1 vccd1 mports_o[121] sky130_fd_sc_hd__buf_12
XANTENNA__7351__S _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6492__A1 _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8233__A2 _8230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6795__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7992__B2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4723__B _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7744__A1 _7349_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output388_A _7947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5507__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8211__A _8211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output722_A _6863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8472__A2 _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__buf_1
XANTENNA__6483__B2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4494__B1 _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8224__A2 _8215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5038__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6235__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6981_ _7272_/B _6989_/B _6980_/Y _6994_/B _7000_/S vssd1 vssd1 vccd1 vccd1 _6981_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7983__B2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5932_ _5932_/A vssd1 vssd1 vccd1 vccd1 _5932_/Y sky130_fd_sc_hd__inv_2
X_8720_ _8293_/X _8806_/B _8718_/X _8719_/Y vssd1 vssd1 vccd1 vccd1 _8720_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4914__A _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8651_ _8036_/Y _8581_/X _8471_/Y _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8651_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5863_ _5863_/A _5863_/B vssd1 vssd1 vccd1 vccd1 _5864_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_146_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7735__A1 _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8932__B1 hold10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7735__B2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7602_ _5930_/Y _7668_/B _6837_/B _7638_/B _7347_/A vssd1 vssd1 vccd1 vccd1 _7602_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4814_ _4814_/A _4814_/B vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5746__B1 _5130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8582_ _8696_/A vssd1 vssd1 vccd1 vccd1 _8583_/A sky130_fd_sc_hd__inv_6
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5794_ _5765_/X _7311_/A _8151_/B _6771_/A vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_145_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7533_ _5682_/Y _8578_/B _8919_/A vssd1 vssd1 vccd1 vccd1 _7533_/Y sky130_fd_sc_hd__a21oi_1
X_4745_ _4745_/A _4745_/B vssd1 vssd1 vccd1 vccd1 _4814_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7464_ _5460_/X _7741_/S _7461_/X _7463_/Y vssd1 vssd1 vccd1 vccd1 _7464_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4676_ _4676_/A vssd1 vssd1 vccd1 vccd1 _4677_/B sky130_fd_sc_hd__inv_2
XFILLER_0_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6415_ _6415_/A _6994_/A vssd1 vssd1 vccd1 vccd1 _6989_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6171__B1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7395_ _5218_/A _7660_/B _7393_/X _7348_/A _7394_/Y vssd1 vssd1 vccd1 vccd1 _7395_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6710__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6346_ _4793_/A _6128_/B _6342_/X _6343_/X _6345_/Y vssd1 vssd1 vccd1 vccd1 _6346_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6576__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6277_ _6277_/A vssd1 vssd1 vccd1 vccd1 _6278_/B sky130_fd_sc_hd__inv_2
Xinput107 mports_i[196] vssd1 vssd1 vccd1 vccd1 _5637_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput118 mports_i[205] vssd1 vssd1 vccd1 vccd1 _5928_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5277__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8016_ _8016_/A vssd1 vssd1 vccd1 vccd1 _8016_/Y sky130_fd_sc_hd__inv_2
X_5228_ _6551_/A _5197_/X _8151_/B _6566_/B vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7671__B1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput129 mports_i[215] vssd1 vssd1 vccd1 vccd1 _6182_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__8215__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5159_ _5159_/A _5159_/B vssd1 vssd1 vccd1 vccd1 _5159_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7974__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6777__A2 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8918_ hold38/X vssd1 vssd1 vccd1 vccd1 _8955_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5985__B1 _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7200__A _7200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5639__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8849_ _8860_/B vssd1 vssd1 vccd1 vccd1 _8850_/B sky130_fd_sc_hd__inv_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5655__A _5655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6162__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7081__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5268__A2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6465__A1 _7332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8206__A2 _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6768__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7965__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8948__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4453__B _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7193__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8579__C _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4530_ _8240_/A _4436_/A _4529_/Y _4528_/B vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4951__A1 _4942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8678__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ _8180_/A _4312_/B _8166_/A vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__mux2_1
XANTENNA__8693__A2 _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6200_ _6304_/A _6931_/A _5715_/B _6199_/X vssd1 vssd1 vccd1 vccd1 _6200_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_110_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7180_ _7295_/S vssd1 vssd1 vccd1 vccd1 _7249_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4392_ _4392_/A _7847_/A vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6131_ _6304_/A _6909_/A _5011_/A vssd1 vssd1 vccd1 vccd1 _6131_/Y sky130_fd_sc_hd__o21ai_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4909__A _4909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _5988_/A _8271_/A _5989_/A _4913_/A _6061_/X vssd1 vssd1 vccd1 vccd1 _6063_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5013_ _7384_/A _6312_/A vssd1 vssd1 vccd1 vccd1 _5013_/Y sky130_fd_sc_hd__nand2_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6759__A2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6843__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7956__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5967__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6964_ _6964_/A vssd1 vssd1 vccd1 vccd1 _6964_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__7020__A _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5431__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8703_ _8247_/Y _8583_/A _8249_/X _8581_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8703_/X
+ sky130_fd_sc_hd__a221o_1
X_5915_ _6875_/B _5839_/X _5914_/Y vssd1 vssd1 vccd1 vccd1 _5915_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4363__B _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6895_ _6889_/Y _6467_/X _6890_/Y _6891_/Y _6894_/Y vssd1 vssd1 vccd1 vccd1 _6895_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__7708__A1 _6241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7708__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5719__B1 _5686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8634_ _8633_/X _7972_/Y _8689_/S vssd1 vssd1 vccd1 vccd1 _8634_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5846_ _5834_/X _5844_/Y _5845_/Y _6170_/A vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__a31o_2
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6916__C1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7184__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5195__A1 _5195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6392__B1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5195__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8565_ _8226_/X _8349_/A _8562_/Y _8564_/X vssd1 vssd1 vccd1 vccd1 _8565_/X sky130_fd_sc_hd__o22a_1
X_5777_ _6906_/A _6802_/A _5776_/Y vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4942__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4728_ _4734_/B _4733_/B vssd1 vssd1 vccd1 vccd1 _4729_/A sky130_fd_sc_hd__nand2_1
X_7516_ _7767_/A _5607_/A _7515_/X vssd1 vssd1 vccd1 vccd1 _7516_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4942__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8496_ _8495_/X _8516_/A _8496_/S vssd1 vssd1 vccd1 vccd1 _8496_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8133__B2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7447_ _7700_/B vssd1 vssd1 vccd1 vccd1 _7606_/A sky130_fd_sc_hd__inv_2
XANTENNA__8684__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4659_ _6941_/A _4657_/X _4658_/X vssd1 vssd1 vccd1 vccd1 _4659_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5498__A2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7378_ _7510_/B vssd1 vssd1 vccd1 vccd1 _7378_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6329_ _6329_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7644__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7947__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8372__B2 _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7584__B _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6383__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5385__A _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6922__A2 _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6135__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6686__B2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7105__A _7105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7635__B1 _7633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output420_A _8155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6944__A _6944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output518_A _7319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7938__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8060__B1 _8067_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5413__A2 _6622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6610__A1 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5700_ _5685_/A _4913_/A _5686_/A _8335_/B _5699_/X vssd1 vssd1 vccd1 vccd1 _7544_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8370__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6680_ _7474_/B _6876_/C _6676_/X _6678_/Y _6679_/Y vssd1 vssd1 vccd1 vccd1 _6681_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8363__A1 _7956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7166__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8363__B2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5177__A1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5631_ _5702_/A _6870_/S vssd1 vssd1 vccd1 vccd1 _5631_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5177__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6374__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8350_ _8344_/Y _8349_/A _8349_/Y vssd1 vssd1 vccd1 vccd1 _8350_/Y sky130_fd_sc_hd__a21oi_4
X_5562_ _5575_/A _5102_/A _5576_/A _5191_/A _5561_/X vssd1 vssd1 vccd1 vccd1 _5562_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_115_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8115__B2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7301_ _7347_/A vssd1 vssd1 vccd1 vccd1 _7753_/B sky130_fd_sc_hd__buf_6
XFILLER_0_41_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4513_ _4455_/A _4455_/B _4456_/B vssd1 vssd1 vccd1 vccd1 _4525_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6126__B1 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8281_ _7803_/Y _8496_/S _8280_/X vssd1 vssd1 vccd1 vccd1 _8281_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5493_ _6202_/B _7470_/A _5136_/X vssd1 vssd1 vccd1 vccd1 _5493_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8666__A2 _8516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7232_ _6221_/Y _7088_/A _6937_/X _7059_/A _7089_/A vssd1 vssd1 vccd1 vccd1 _7232_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4444_ hold23/X vssd1 vssd1 vccd1 vccd1 _8189_/B sky130_fd_sc_hd__clkinv_8
XFILLER_0_123_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7163_ _6771_/A _7023_/X _7162_/X vssd1 vssd1 vccd1 vccd1 _7163_/X sky130_fd_sc_hd__o21a_1
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _8966_/D sky130_fd_sc_hd__buf_2
XANTENNA__6429__A1 _4942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6114_ _6141_/A1 _4953_/X _6141_/B1 _5089_/X _6113_/X vssd1 vssd1 vccd1 vccd1 _6115_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7626__B1 _7624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7094_/A vssd1 vssd1 vccd1 vccd1 _7094_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6547_/A _6041_/X _6044_/Y vssd1 vssd1 vccd1 vccd1 _7648_/B sky130_fd_sc_hd__o21ai_2
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6854__A _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5652__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7929__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7996_ _7989_/Y _6500_/A _7990_/Y _7769_/A _7995_/Y vssd1 vssd1 vccd1 vccd1 _8424_/A
+ sky130_fd_sc_hd__a221oi_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5404__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5189__B _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6947_ _8857_/B _6947_/B vssd1 vssd1 vccd1 vccd1 _6947_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6878_ _6435_/A _6877_/X _5997_/A _6473_/A vssd1 vssd1 vccd1 vccd1 _6878_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5168__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8617_ _7901_/Y _8581_/X _7903_/Y _8583_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8617_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6365__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5168__B2 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4821__B _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5829_ _8160_/A _6231_/C _5829_/C vssd1 vssd1 vccd1 vccd1 _5830_/A sky130_fd_sc_hd__or3_1
XFILLER_0_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6904__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8548_ _8130_/Y hold36/A _8482_/B vssd1 vssd1 vccd1 vccd1 _8548_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_45_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8106__A1 _8106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8106__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8479_ _8479_/A vssd1 vssd1 vccd1 vccd1 _8479_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8409__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5340__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6840__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8593__A1 _7786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8593__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5827__B _5827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8896__A2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5319__S _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output468_A _7880_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7320__A2 _7347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6658__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5331__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5331__B2 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5882__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7084__A1 _7422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8963__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput290 sports_i[31] vssd1 vssd1 vccd1 vccd1 _8234_/A2 sky130_fd_sc_hd__clkbuf_2
X_7850_ _7840_/Y _5146_/A _7841_/Y _7431_/B _7849_/X vssd1 vssd1 vccd1 vccd1 _7851_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__7387__A2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6801_ _6801_/A _6801_/B vssd1 vssd1 vccd1 vccd1 _6801_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5398__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4993_ _4990_/X _4992_/X _6356_/S vssd1 vssd1 vccd1 vccd1 _4993_/X sky130_fd_sc_hd__mux2_1
X_7781_ _7777_/X _8295_/A _7975_/A vssd1 vssd1 vccd1 vccd1 _7781_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__6595__B1 _7413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4922__A _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6732_ _6732_/A vssd1 vssd1 vccd1 vccd1 _6733_/A sky130_fd_sc_hd__inv_2
XFILLER_0_86_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5737__B _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6663_ _7470_/A _6801_/A _6450_/A _6662_/Y vssd1 vssd1 vccd1 vccd1 _6663_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8402_ _8555_/B _8454_/A _8441_/B _8376_/A vssd1 vssd1 vccd1 vccd1 _8402_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5614_ _6837_/A _5608_/X _5613_/X vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6898__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6594_ _6547_/A _5306_/X _6593_/X vssd1 vssd1 vccd1 vccd1 _6594_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5545_ _6202_/B _5544_/X _5136_/X vssd1 vssd1 vccd1 vccd1 _5545_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8333_ _8333_/A vssd1 vssd1 vccd1 vccd1 _8334_/A sky130_fd_sc_hd__inv_2
XANTENNA__5570__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8639__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8264_ _8264_/A _8574_/B vssd1 vssd1 vccd1 vccd1 _8497_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_42_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5476_ _7524_/A _7299_/A _6281_/S _6727_/B vssd1 vssd1 vccd1 vccd1 _5674_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput720 _6836_/X vssd1 vssd1 vccd1 vccd1 sports_o[91] sky130_fd_sc_hd__buf_12
XFILLER_0_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4427_ _4427_/A hold40/A vssd1 vssd1 vccd1 vccd1 _4526_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7215_ _6112_/B _7026_/X _7214_/X vssd1 vssd1 vccd1 vccd1 _7215_/X sky130_fd_sc_hd__o21a_1
X_8195_ _8193_/Y _8194_/Y hold44/A vssd1 vssd1 vccd1 vccd1 _8195_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5873__A2 _5902_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7146_ _7145_/X _5655_/A _7175_/S vssd1 vssd1 vccd1 vccd1 _7147_/A sky130_fd_sc_hd__mux2_1
X_4358_ hold45/X hold39/X vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__nor2_2
XANTENNA__7075__A1 _6578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7075__B2 _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7077_ _7076_/X _5239_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__mux2_1
X_6028_ _6028_/A vssd1 vssd1 vccd1 vccd1 _6029_/B sky130_fd_sc_hd__inv_2
XFILLER_0_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7979_ _7976_/Y _5117_/A _7977_/Y _7013_/A _7978_/Y vssd1 vssd1 vccd1 vccd1 _8390_/A
+ sky130_fd_sc_hd__a221oi_4
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6050__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8304__A _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8327__A1 _7888_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8327__B2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8878__A2 _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7550__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5561__A1 _5587_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5561__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7838__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7066__A1 _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8263__B1 _7763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7066__B2 _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6494__A _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8802__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8566__A1 _8239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7369__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8566__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6577__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6941__B _6941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8318__A1 _8317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6592__A3 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7781__B1_N _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7541__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5552__A1 _5591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5552__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6669__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7264__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5330_ _8842_/B _5363_/B _5329_/Y vssd1 vssd1 vccd1 vccd1 _5330_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5292__B _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5261_ _5257_/Y _5260_/Y _7852_/A vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5304__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5304__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6501__B1 _5062_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7000_ _6999_/X _7754_/B _7000_/S vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__mux2_1
X_5192_ _5192_/A vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__7057__A1 _7356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4917__A _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8951_ _8967_/CLK hold25/X fanout733/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__8006__B1 _8011_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6280__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7902_ _7905_/A1 _5780_/X _7905_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7902_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8882_ _4818_/B _4930_/X _4662_/C _8574_/B vssd1 vssd1 vccd1 vccd1 _8882_/Y sky130_fd_sc_hd__o31ai_1
X_7833_ _7825_/X _7826_/X _7832_/Y _7768_/X _7774_/X vssd1 vssd1 vccd1 vccd1 _7833_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6851__B _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5748__A _5829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6032__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7764_ _6080_/A _7779_/B1 _6513_/A _4331_/B vssd1 vssd1 vccd1 vccd1 _7764_/X sky130_fd_sc_hd__a22o_1
X_4976_ _4976_/A vssd1 vssd1 vccd1 vccd1 _4976_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8309__A1 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8309__B2 _7809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7780__A2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6715_ _5628_/A _6467_/X _6713_/X _6714_/X _6450_/A vssd1 vssd1 vccd1 vccd1 _6715_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5791__A1 _6770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5791__B2 _6788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7695_ _6937_/A _7660_/B _6221_/Y _7349_/A _7694_/Y vssd1 vssd1 vccd1 vccd1 _7695_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6646_ _6852_/A _6646_/B vssd1 vssd1 vccd1 vccd1 _6646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5543__A1 _5543_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5543__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6577_ _6432_/X _6576_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6577_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6740__B1 _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8316_ _8316_/A _8364_/A vssd1 vssd1 vccd1 vccd1 _8316_/Y sky130_fd_sc_hd__nand2_1
X_5528_ _5031_/X _5496_/X _5527_/X vssd1 vssd1 vccd1 vccd1 _5528_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5459_ input98/X _8706_/B input36/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__o22a_1
X_8247_ _8247_/A vssd1 vssd1 vccd1 vccd1 _8247_/Y sky130_fd_sc_hd__inv_2
Xoutput550 _7567_/X vssd1 vssd1 vccd1 vccd1 sports_o[143] sky130_fd_sc_hd__buf_12
Xoutput561 _7658_/X vssd1 vssd1 vccd1 vccd1 sports_o[153] sky130_fd_sc_hd__buf_12
Xoutput572 _7726_/Y vssd1 vssd1 vccd1 vccd1 sports_o[163] sky130_fd_sc_hd__buf_12
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput583 _4997_/X vssd1 vssd1 vccd1 vccd1 sports_o[173] sky130_fd_sc_hd__buf_12
Xoutput594 _5332_/X vssd1 vssd1 vccd1 vccd1 sports_o[183] sky130_fd_sc_hd__buf_12
X_8178_ _8192_/A _8181_/A vssd1 vssd1 vccd1 vccd1 _8179_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8245__B1 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7129_ _7129_/A vssd1 vssd1 vccd1 vccd1 _7129_/X sky130_fd_sc_hd__buf_1
XANTENNA__8548__A1 _8130_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6761__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6023__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7220__A1 _6102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5658__A _5658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4562__A _7876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7771__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4585__A2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7523__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7592__B _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6489__A _6489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6001__B _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5837__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7039__A1 _5064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8236__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8787__A1 _8458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6262__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output500_A _8699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8539__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7767__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6671__B _6671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7259__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6014__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7211__A1 _6107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ _4830_/A _7398_/A vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__B1 _5222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7762__A2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4761_ _4761_/A _4770_/A _4770_/B vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__nand3_1
XANTENNA__5773__A1 _5770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5773__B2 _5772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6500_ _6500_/A vssd1 vssd1 vccd1 vccd1 _6500_/X sky130_fd_sc_hd__buf_12
XFILLER_0_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7480_ _7121_/A _7630_/B _5516_/X _7638_/B vssd1 vssd1 vccd1 vccd1 _7480_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_126_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4692_ _4692_/A vssd1 vssd1 vccd1 vccd1 _4692_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_126_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5525__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6431_ _6854_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _6432_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5525__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6362_ _6369_/A1 _8523_/B input14/X _4933_/A _6361_/X vssd1 vssd1 vccd1 vccd1 _7746_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_141_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5313_ _5313_/A vssd1 vssd1 vccd1 vccd1 _6870_/S sky130_fd_sc_hd__clkbuf_8
X_8101_ _8106_/A1 _5146_/A _8106_/B1 _5616_/A vssd1 vssd1 vccd1 vccd1 _8101_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7007__B _7272_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6293_ _6326_/A1 _8523_/B input9/X _4933_/A _6292_/X vssd1 vssd1 vccd1 vccd1 _7729_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5289__B1 _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5244_ _5272_/A _8271_/A _5273_/A _5191_/X _5243_/X vssd1 vssd1 vccd1 vccd1 _5356_/B
+ sky130_fd_sc_hd__o221a_4
X_8032_ _5359_/A _8030_/Y _5116_/A _8031_/Y vssd1 vssd1 vccd1 vccd1 _8032_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6846__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__buf_2
XANTENNA__8227__B1 _8235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6338__S _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4647__A _8958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5175_ _5909_/B _5161_/X _6557_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__a22o_1
XANTENNA__7023__A _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4366__B _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8934_ _8934_/A _8934_/B _8934_/C vssd1 vssd1 vccd1 vccd1 _8935_/B sky130_fd_sc_hd__nand3_1
XANTENNA__5461__A0 _5458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8865_ _8865_/A _8865_/B vssd1 vssd1 vccd1 vccd1 _8865_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6581__B _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6005__A2 _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7169__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7202__A1 _6867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7816_ _7760_/X _7807_/X _7812_/X _7815_/Y vssd1 vssd1 vccd1 vccd1 _7816_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_94_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8796_ _8796_/A vssd1 vssd1 vccd1 vccd1 _8796_/X sky130_fd_sc_hd__buf_1
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7747_ _7745_/X _7332_/A _7746_/Y vssd1 vssd1 vccd1 vccd1 _7747_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__5764__A1 _5764_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4959_ _4956_/Y _8455_/B _4957_/Y _4891_/X _4958_/Y vssd1 vssd1 vccd1 vccd1 _4960_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5764__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7678_ _7678_/A _7678_/B vssd1 vssd1 vccd1 vccd1 _7678_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8702__B2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6629_ _6628_/B _6613_/B _6628_/Y vssd1 vssd1 vccd1 vccd1 _6629_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6102__A _6102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput380 _8758_/X vssd1 vssd1 vccd1 vccd1 mports_o[112] sky130_fd_sc_hd__buf_12
Xoutput391 _8792_/X vssd1 vssd1 vccd1 vccd1 mports_o[122] sky130_fd_sc_hd__buf_12
XANTENNA__6756__B _6756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8218__B1 _4312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5660__B _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6492__A2 _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8029__A _8029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7992__A2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6491__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4292__A _7683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__B1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5755__A1 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5755__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6711__S _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5507__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5507__B2 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6704__B1 _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output450_A _8463_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6947__A _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6468__C1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4494__A1 _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4494__B2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6235__A2 _6207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7778__A _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8373__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6980_ _8919_/A _6980_/B vssd1 vssd1 vccd1 vccd1 _6980_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__7983__A2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6640__C1 _6639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5931_ _5931_/A vssd1 vssd1 vccd1 vccd1 _5931_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5298__A _5333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8650_ _8650_/A vssd1 vssd1 vccd1 vccd1 _8650_/X sky130_fd_sc_hd__buf_1
X_5862_ _5862_/A _6593_/A vssd1 vssd1 vccd1 vccd1 _5863_/B sky130_fd_sc_hd__nand2_1
XANTENNA__7735__A2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7601_ _7510_/B _5899_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7606_/B sky130_fd_sc_hd__o21a_1
X_4813_ _4819_/C _4813_/B _4813_/C vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__nand3_1
X_8581_ _8581_/A vssd1 vssd1 vccd1 vccd1 _8581_/X sky130_fd_sc_hd__buf_4
X_5793_ _5722_/A _5102_/A _5723_/A _5191_/X _5792_/X vssd1 vssd1 vccd1 vccd1 _6771_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5746__B2 _5788_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4930__A _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7532_ _7532_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _7532_/Y sky130_fd_sc_hd__nor2_1
X_4744_ _4744_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _4745_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_145_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7463_ _7463_/A _7691_/B vssd1 vssd1 vccd1 vccd1 _7463_/Y sky130_fd_sc_hd__nand2_1
X_4675_ _4675_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7018__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6414_ _6488_/B vssd1 vssd1 vccd1 vccd1 _6994_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6171__A1 _6182_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6171__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7394_ _7575_/A _7394_/B vssd1 vssd1 vccd1 vccd1 _7394_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_114_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6345_ _6345_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6345_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6276_ _6299_/A _4868_/A input8/X _5089_/A _6275_/X vssd1 vssd1 vccd1 vccd1 _6277_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6576__B _6576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput108 mports_i[197] vssd1 vssd1 vccd1 vccd1 _5697_/A1 sky130_fd_sc_hd__buf_2
X_5227_ _5248_/A _5197_/X _8151_/B _5323_/A vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__a22o_1
X_8015_ _8015_/A vssd1 vssd1 vccd1 vccd1 _8015_/Y sky130_fd_sc_hd__inv_2
Xinput119 mports_i[206] vssd1 vssd1 vccd1 vccd1 _5962_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5158_ _5159_/A _5361_/A vssd1 vssd1 vccd1 vccd1 _6536_/B sky130_fd_sc_hd__nand2_1
XANTENNA__8620__B1 _7916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7423__B2 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5089_ _5089_/A vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__buf_8
XANTENNA__7974__A2 _8375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8917_ _4406_/B _8185_/B _8917_/S vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__mux2_1
XANTENNA__4824__B _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8848_ _8848_/A _8848_/B vssd1 vssd1 vccd1 vccd1 _8860_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5001__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7726__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8779_ _8833_/B _8012_/Y _8725_/A vssd1 vssd1 vccd1 vccd1 _8779_/X sky130_fd_sc_hd__o21a_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6934__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5936__A _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5655__B _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6162__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7111__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5390__B _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7662__A1 _6112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7662__B2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5673__B1 _5011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8611__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7414__B2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7965__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5976__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5976__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7110__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7178__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5728__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4460_ _4460_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7350__B1 _7349_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6677__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4391_ _4406_/A _4405_/A vssd1 vssd1 vccd1 vccd1 _4425_/C sky130_fd_sc_hd__nor2_1
XANTENNA__5900__A1 _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5581__A _6695_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6130_ _5159_/B _6094_/X _5125_/X _6926_/B _6129_/X vssd1 vssd1 vccd1 vccd1 _6130_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6061_/A1 _8271_/B input59/X _4917_/A vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__o22a_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7653__A1 _6107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7653__B2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5055_/A _6474_/A vssd1 vssd1 vccd1 vccd1 _5012_/Y sky130_fd_sc_hd__nor2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5416__B1 _5386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7956__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7301__A _7347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5967__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6963_ _6962_/X _7720_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6964_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_88_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8702_ _8700_/Y _8701_/X _4662_/C _8577_/X vssd1 vssd1 vccd1 vccd1 _8702_/X sky130_fd_sc_hd__a22o_1
X_5914_ _5914_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _5914_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7169__A0 _7168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6894_ _6107_/A _6801_/A _6924_/A _6893_/Y _6450_/A vssd1 vssd1 vccd1 vccd1 _6894_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_146_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7708__A2 _7347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5719__A1 _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8633_ _8404_/A _8581_/A _7969_/Y _8583_/A vssd1 vssd1 vccd1 vccd1 _8633_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5845_ _5845_/A _5845_/B vssd1 vssd1 vccd1 vccd1 _5845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5719__B2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6916__B1 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5195__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8564_ _8564_/A _8564_/B vssd1 vssd1 vccd1 vccd1 _8564_/X sky130_fd_sc_hd__and2_1
XFILLER_0_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6392__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8118__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5776_ _6744_/B _6906_/A vssd1 vssd1 vccd1 vccd1 _5776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8669__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7515_ _7514_/Y _7297_/B _7575_/A _7385_/Y vssd1 vssd1 vccd1 vccd1 _7515_/X sky130_fd_sc_hd__a31o_1
X_4727_ _4732_/B _4731_/A _4727_/C vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__nand3_1
XANTENNA__4942__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8495_ _8511_/A _8304_/A _8091_/Y _8299_/A vssd1 vssd1 vccd1 vccd1 _8495_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8133__A2 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7446_ _7442_/X _7444_/Y _7445_/Y vssd1 vssd1 vccd1 vccd1 _7446_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4658_ _4658_/A _8194_/A _8845_/C vssd1 vssd1 vccd1 vccd1 _4658_/X sky130_fd_sc_hd__or3_1
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 mports_i[180] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8278__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7892__A1 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7377_ _6538_/A _7619_/B _7369_/X _7374_/Y _7376_/Y vssd1 vssd1 vccd1 vccd1 _7377_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4589_ _4589_/A _7309_/B vssd1 vssd1 vccd1 vccd1 _4590_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6328_ _6312_/A _7729_/B _6264_/X vssd1 vssd1 vccd1 vccd1 _6329_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__7644__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6259_ _6262_/A1 _8716_/B input69/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6259_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7947__A2 _8376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6604__C1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8372__A2 _8346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5666__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4570__A _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6383__A1 _6387_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6383__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6135__B2 _6102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8188__S _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6497__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7092__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7635__A1 _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7105__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8832__B1 _8232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7635__B2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output413_A _7794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7399__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7938__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8060__A1 _8067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5949__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4464__B _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6610__A2 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8363__A2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5630_ _5630_/A vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__inv_2
XANTENNA__4480__A _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6374__A1 _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5177__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5561_ _5587_/A1 _5192_/X input41/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_54_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8115__A2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7300_ _7686_/A _7575_/A vssd1 vssd1 vccd1 vccd1 _7347_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4512_ _4605_/B _4611_/B vssd1 vssd1 vccd1 vccd1 _4603_/B sky130_fd_sc_hd__nand2_1
X_5492_ _5440_/A _5102_/A _5441_/A _5191_/A _5491_/X vssd1 vssd1 vccd1 vccd1 _7470_/A
+ sky130_fd_sc_hd__o221a_4
X_8280_ _7798_/X _8429_/A _7800_/X _8299_/A _8269_/A vssd1 vssd1 vccd1 vccd1 _8280_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7231_ _7231_/A vssd1 vssd1 vccd1 vccd1 _7231_/X sky130_fd_sc_hd__buf_1
X_4443_ _4443_/A vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__inv_2
XFILLER_0_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5515__S _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5885__B1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7162_ _6758_/B _7004_/X _7560_/A _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7162_/X
+ sky130_fd_sc_hd__a221o_2
X_4374_ _4307_/X hold40/A _8239_/A _4412_/C _4373_/Y vssd1 vssd1 vccd1 vccd1 _4375_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4639__B _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6113_ _6140_/A1 _8709_/B input63/X _5091_/X vssd1 vssd1 vccd1 vccd1 _6113_/X sky130_fd_sc_hd__o22a_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8823__B1 _8206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7093_ _7093_/A vssd1 vssd1 vccd1 vccd1 _7093_/X sky130_fd_sc_hd__buf_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7626__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6044_ _7632_/B _6547_/A vssd1 vssd1 vccd1 vccd1 _6044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4655__A _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7031__A _7031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7929__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8051__A1 _8054_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8051__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7995_ _7998_/A1 _5780_/A _7998_/B1 _5079_/A vssd1 vssd1 vccd1 vccd1 _7995_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_0_95_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6062__B1 _5989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6601__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6946_ _6945_/X _6207_/A _6946_/S vssd1 vssd1 vccd1 vccd1 _6947_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6877_ _7639_/A _6475_/A _6432_/A vssd1 vssd1 vccd1 vccd1 _6877_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_49_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6081__S _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8616_ _8616_/A vssd1 vssd1 vccd1 vccd1 _8616_/X sky130_fd_sc_hd__buf_1
XANTENNA__6365__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5168__A2 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5828_ _5845_/A _7384_/A vssd1 vssd1 vccd1 vccd1 _5828_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6365__B2 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8547_ _8547_/A vssd1 vssd1 vccd1 vccd1 _8547_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5759_ _5759_/A vssd1 vssd1 vccd1 vccd1 _5760_/A sky130_fd_sc_hd__inv_2
XANTENNA__8106__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6117__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8478_ _8477_/X _8434_/X _8555_/B vssd1 vssd1 vccd1 vccd1 _8479_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7429_ _6613_/B _7619_/B _7425_/X _7427_/Y _7428_/Y vssd1 vssd1 vccd1 vccd1 _7429_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5340__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7617__A1 _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4565__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8042__B2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8593__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7876__A _7876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6780__A _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7553__A0 _7552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8896__A3 _4662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6020__A _6020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5331__A2 _5328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7608__A1 _7683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output628_A _6191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5619__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8281__A1 _7803_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7084__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5095__A1 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6292__B1 _6314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput280 sports_i[22] vssd1 vssd1 vccd1 vccd1 _8085_/A sky130_fd_sc_hd__buf_1
Xinput291 sports_i[32] vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8971__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6800_ _7577_/B _6871_/B vssd1 vssd1 vccd1 vccd1 _6800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5398__A2 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7780_ _4318_/B _5230_/B _4481_/B _5197_/X _7779_/X vssd1 vssd1 vccd1 vccd1 _8295_/A
+ sky130_fd_sc_hd__a221o_4
X_4992_ _4975_/A _8516_/B _4976_/A _4913_/X _4991_/X vssd1 vssd1 vccd1 vccd1 _4992_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6595__B2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6731_ _6924_/A _6731_/B vssd1 vssd1 vccd1 vccd1 _6731_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4922__B _7876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6662_ _6662_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6662_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6347__A1 _7737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8401_ _8400_/Y _8375_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8454_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_128_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5613_ _6780_/A _5613_/B vssd1 vssd1 vccd1 vccd1 _5613_/X sky130_fd_sc_hd__or2_1
XANTENNA__6898__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6593_ _6593_/A _6593_/B vssd1 vssd1 vccd1 vccd1 _6593_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8332_ _8346_/A _8323_/X _8330_/X _8331_/X vssd1 vssd1 vccd1 vccd1 _8332_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5544_ _5510_/A _5102_/A _5511_/A _5191_/A _5543_/X vssd1 vssd1 vccd1 vccd1 _5544_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5570__A2 _5548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8263_ _8574_/A _8215_/X _7763_/X _8264_/A vssd1 vssd1 vccd1 vccd1 _8263_/X sky130_fd_sc_hd__a22o_1
X_5475_ _5661_/A _4953_/X _5662_/A _5089_/X _5474_/X vssd1 vssd1 vccd1 vccd1 _6727_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput710 _6723_/X vssd1 vssd1 vccd1 vccd1 sports_o[82] sky130_fd_sc_hd__buf_12
XFILLER_0_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput721 _6850_/X vssd1 vssd1 vccd1 vccd1 sports_o[92] sky130_fd_sc_hd__buf_12
XANTENNA__7026__A _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7214_ _7660_/A _7004_/X _6897_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7214_/X
+ sky130_fd_sc_hd__a221o_1
X_4426_ _4426_/A _5827_/B vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8194_ _8194_/A _8194_/B vssd1 vssd1 vccd1 vccd1 _8194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7145_ _5625_/A _7023_/X _7144_/X vssd1 vssd1 vccd1 vccd1 _7145_/X sky130_fd_sc_hd__o21a_1
X_4357_ _4422_/B vssd1 vssd1 vccd1 vccd1 _4412_/C sky130_fd_sc_hd__inv_4
XFILLER_0_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7075__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7076_ _5248_/A _7023_/X _7075_/X vssd1 vssd1 vccd1 vccd1 _7076_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5086__A1 _5070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6584__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5086__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6027_ _5999_/B _7630_/A _6026_/X _5174_/A vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4385__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6822__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8024__A1 _8024_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8024__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7232__C1 _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7696__A _7696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7978_ _7985_/A1 _4947_/B _7985_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _7978_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__6586__A1 _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7783__B1 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6929_ _7683_/A _6510_/A _6928_/Y _6512_/A vssd1 vssd1 vccd1 vccd1 _6929_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8327__A2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4551__C _7707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5561__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7838__A1 _7837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7066__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8263__B2 _8264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6274__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4295__A _4408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8566__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6577__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4742__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5552__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6669__B _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _7413_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _5260_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5304__A2 _5280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6501__A1 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6501__B2 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5191_ _5191_/A vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__buf_8
XFILLER_0_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7280__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8254__A1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5068__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6265__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8950_ _8967_/CLK _8950_/D fanout733/X vssd1 vssd1 vccd1 vccd1 _8950_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4815__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7901_ _7896_/Y _6965_/A _7897_/Y _8163_/A _7900_/Y vssd1 vssd1 vccd1 vccd1 _7901_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__8006__A1 _8011_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8006__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8881_ _8879_/Y _4818_/A _8880_/Y vssd1 vssd1 vccd1 vccd1 _8884_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7214__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7832_ _7832_/A vssd1 vssd1 vccd1 vccd1 _7832_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__4933__A _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7765__B1 _4481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7763_ _4318_/B _5359_/B _4481_/B _7316_/A _7762_/X vssd1 vssd1 vccd1 vccd1 _7763_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4975_ _4975_/A vssd1 vssd1 vccd1 vccd1 _4975_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6714_ _5659_/A _6549_/A _5574_/X _6876_/C _7000_/S vssd1 vssd1 vccd1 vccd1 _6714_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5791__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7694_ _7694_/A _7694_/B vssd1 vssd1 vccd1 vccd1 _7694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6645_ _6645_/A _6694_/B vssd1 vssd1 vccd1 vccd1 _6645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8140__A _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5543__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6576_ _6852_/A _6576_/B vssd1 vssd1 vccd1 vccd1 _6576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8315_ _8315_/A vssd1 vssd1 vccd1 vccd1 _8315_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5527_ _6128_/B _5498_/X _5503_/X _5526_/X _6402_/A vssd1 vssd1 vccd1 vccd1 _5527_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8246_ _8251_/A2 _7769_/X _8252_/A1 _5682_/B _8245_/X vssd1 vssd1 vccd1 vccd1 _8247_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5458_ _5455_/X _7459_/A _6356_/S vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__mux2_2
Xoutput540 _7486_/X vssd1 vssd1 vccd1 vccd1 sports_o[134] sky130_fd_sc_hd__buf_12
XFILLER_0_112_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput551 _7573_/X vssd1 vssd1 vccd1 vccd1 sports_o[144] sky130_fd_sc_hd__buf_12
Xoutput562 _7667_/X vssd1 vssd1 vccd1 vccd1 sports_o[154] sky130_fd_sc_hd__buf_12
X_4409_ _4409_/A hold40/A vssd1 vssd1 vccd1 vccd1 _4504_/B sky130_fd_sc_hd__nand2_1
Xoutput573 _7730_/Y vssd1 vssd1 vccd1 vccd1 sports_o[164] sky130_fd_sc_hd__buf_12
Xoutput584 _5030_/X vssd1 vssd1 vccd1 vccd1 sports_o[174] sky130_fd_sc_hd__buf_12
X_8177_ _7975_/X _8157_/X _8170_/X _8176_/Y vssd1 vssd1 vccd1 vccd1 _8177_/X sky130_fd_sc_hd__a22o_2
Xoutput595 _5376_/X vssd1 vssd1 vccd1 vccd1 sports_o[184] sky130_fd_sc_hd__buf_12
X_5389_ _6079_/A _5425_/C vssd1 vssd1 vccd1 vccd1 _5389_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7190__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7128_ _7127_/X _5548_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7129_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8245__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8245__B2 _8251_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7059_ _7059_/A vssd1 vssd1 vccd1 vccd1 _7059_/X sky130_fd_sc_hd__buf_6
XANTENNA__5004__A _5004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6008__B1 _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7205__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8315__A _8315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7220__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5674__A _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8720__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6794__A1_N _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7287__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7039__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8236__A1 _8235_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6247__B1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7995__B1 _7998_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4753__A _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7211__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7762__A3 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4760_ _4760_/A _4760_/B vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5773__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6970__A1 _7725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4691_ _4734_/B _8578_/B vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7275__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5584__A _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6430_ _6430_/A vssd1 vssd1 vccd1 vccd1 _6430_/X sky130_fd_sc_hd__buf_1
XFILLER_0_153_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6722__A1 _5655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6722__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6361_ _6368_/A1 _8368_/A input76/X _4940_/A vssd1 vssd1 vccd1 vccd1 _6361_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_113_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8100_ _8097_/Y _5117_/A _8098_/Y _7013_/A _8099_/Y vssd1 vssd1 vccd1 vccd1 _8499_/A
+ sky130_fd_sc_hd__a221oi_4
X_5312_ _5304_/X _6233_/B _6170_/A _5311_/X vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__a211o_1
X_6292_ _6315_/B _8368_/A _6314_/B _4940_/A vssd1 vssd1 vccd1 vccd1 _6292_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_122_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5289__A1 _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8031_ _8031_/A vssd1 vssd1 vccd1 vccd1 _8031_/Y sky130_fd_sc_hd__inv_2
X_5243_ input94/X _5192_/X input31/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4928__A _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7304__A _7304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8227__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8227__B2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5174_ _5174_/A vssd1 vssd1 vccd1 vccd1 _5997_/B sky130_fd_sc_hd__buf_6
XANTENNA__4647__B hold44/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6238__B1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8778__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8933_ _8933_/A _8933_/B vssd1 vssd1 vccd1 vccd1 _8934_/C sky130_fd_sc_hd__and2_1
XFILLER_0_36_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5461__A1 _5460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8864_ _8862_/Y _6264_/X _8863_/X vssd1 vssd1 vccd1 vccd1 _8970_/D sky130_fd_sc_hd__a21bo_1
XFILLER_0_148_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7815_ _8284_/B _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _7815_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7202__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8795_ _8794_/X _8476_/A _8829_/S vssd1 vssd1 vccd1 vccd1 _8796_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7746_ _7756_/A _7746_/B vssd1 vssd1 vccd1 vccd1 _7746_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4958_ _4893_/A input81/X _4896_/A input18/X vssd1 vssd1 vccd1 vccd1 _4958_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__6961__A1 _6283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5764__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6961__B2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7677_ _7672_/Y _7673_/X _7675_/X _7676_/X vssd1 vssd1 vccd1 vccd1 _7677_/X sky130_fd_sc_hd__a31o_1
X_4889_ _5130_/A vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__inv_6
XFILLER_0_151_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6628_ _6628_/A _6628_/B vssd1 vssd1 vccd1 vccd1 _6628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6559_ _6432_/X _6558_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6559_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6102__B _6102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8229_ _8229_/A _8229_/B vssd1 vssd1 vccd1 vccd1 _8696_/B sky130_fd_sc_hd__nor2_2
Xoutput370 _8727_/X vssd1 vssd1 vccd1 vccd1 mports_o[103] sky130_fd_sc_hd__buf_12
Xoutput381 _8763_/X vssd1 vssd1 vccd1 vccd1 mports_o[113] sky130_fd_sc_hd__buf_12
Xoutput392 _8796_/X vssd1 vssd1 vccd1 vccd1 mports_o[123] sky130_fd_sc_hd__buf_12
XANTENNA__8218__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8218__B2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4557__B _4557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6229__B1 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4292__B _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5204__A1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6401__B1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5204__B2 _4937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6952__A1 _7707_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8154__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5507__A2 _5557_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8209__A1 _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4494__A2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7968__B1 _7971_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5443__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5579__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5930_ _5930_/A vssd1 vssd1 vccd1 vccd1 _5930_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6686__A1_N _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5861_ _5079_/A _5857_/Y _7852_/A _5860_/Y vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7600_ _5926_/B _7619_/B _7596_/Y _7598_/Y _7599_/Y vssd1 vssd1 vccd1 vccd1 _7600_/X
+ sky130_fd_sc_hd__a221o_1
X_4812_ _4789_/A _4789_/B _4837_/A vssd1 vssd1 vccd1 vccd1 _4819_/C sky130_fd_sc_hd__a21oi_1
X_8580_ _8580_/A vssd1 vssd1 vccd1 vccd1 _8581_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5792_ _5792_/A1 _5192_/X input49/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5792_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5746__A2 _5788_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6943__A1 _6941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7531_ _7531_/A _8755_/C vssd1 vssd1 vccd1 vccd1 _7531_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4954__B1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4743_ _8919_/A vssd1 vssd1 vccd1 vccd1 _7266_/B sky130_fd_sc_hd__inv_6
XFILLER_0_22_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7462_ _7701_/A _5460_/X _6264_/X vssd1 vssd1 vccd1 vccd1 _7463_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__7499__A2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6203__A _6212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4674_ _4674_/A _4674_/B _4674_/C vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__nand3_1
X_6413_ _6919_/A _6724_/A vssd1 vssd1 vccd1 vccd1 _6488_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8829__S _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7393_ _7767_/A _5282_/Y _7071_/A _7630_/B vssd1 vssd1 vccd1 vccd1 _7393_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6171__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6344_ _6312_/A _7737_/B _6264_/X vssd1 vssd1 vccd1 vccd1 _6345_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6275_ _6309_/A1 _4871_/A input71/X _5091_/A vssd1 vssd1 vccd1 vccd1 _6275_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4658__A _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8014_ _7975_/X _8412_/A _8010_/X _8013_/X vssd1 vssd1 vccd1 vccd1 _8014_/X sky130_fd_sc_hd__a22o_2
Xinput109 mports_i[198] vssd1 vssd1 vccd1 vccd1 _5718_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__5131__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5226_ input34/X _8335_/B _5326_/B1 _4913_/A _5225_/X vssd1 vssd1 vccd1 vccd1 _5323_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__7671__A2 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5157_ _5359_/A vssd1 vssd1 vccd1 vccd1 _5361_/A sky130_fd_sc_hd__inv_2
XANTENNA__8620__A1 _8352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7423__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8620__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5088_ _5079_/X _6499_/A _4518_/A _5150_/A _5087_/Y vssd1 vssd1 vccd1 vccd1 _5088_/X
+ sky130_fd_sc_hd__o221a_1
X_8916_ _8916_/A vssd1 vssd1 vccd1 vccd1 _8954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5985__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8847_ _8847_/A vssd1 vssd1 vccd1 vccd1 _8848_/B sky130_fd_sc_hd__inv_2
XANTENNA__8384__B1 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8778_ _8418_/Y _7629_/B _8713_/C _8755_/A _8777_/X vssd1 vssd1 vccd1 vccd1 _8778_/X
+ sky130_fd_sc_hd__a41o_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ _7756_/A _7729_/B vssd1 vssd1 vccd1 vccd1 _7729_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8136__B1 _8150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6162__A2 _6183_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7111__A1 _5465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7662__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5673__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8474__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7598__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8611__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7414__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7178__A1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8503__A _8503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8127__B1 _8132_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7119__A _7119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8678__A1 _8148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8678__B2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7350__A1 _6499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7350__B2 _6497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7553__S _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _4390_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8957__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6677__B _7120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4478__A _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _8842_/B _6058_/Y _6059_/Y vssd1 vssd1 vccd1 vccd1 _6060_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__7653__A2 _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5664__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5011_ _5011_/A vssd1 vssd1 vccd1 vccd1 _5011_/Y sky130_fd_sc_hd__inv_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8602__A1 _8320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7405__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5416__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5416__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6962_ _6961_/X _6287_/X _7000_/S vssd1 vssd1 vccd1 vccd1 _6962_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5967__A2 _6031_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5102__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5913_ _5948_/B _5860_/Y _8189_/A vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__mux2_1
X_8701_ _8239_/Y _8581_/A _8240_/Y _8583_/A _8621_/S vssd1 vssd1 vccd1 vccd1 _8701_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7169__A1 _5772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6893_ _8150_/A _6108_/B _6892_/X vssd1 vssd1 vccd1 vccd1 _6893_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__8366__B1 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8632_ _8369_/A _8577_/X _8630_/X _8631_/X vssd1 vssd1 vccd1 vccd1 _8632_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5844_ _7584_/A _6133_/B vssd1 vssd1 vccd1 vccd1 _5844_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5719__A2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6916__A1 _6102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8563_ _8230_/Y _8299_/A _8232_/X _8304_/A vssd1 vssd1 vccd1 vccd1 _8564_/A sky130_fd_sc_hd__a22o_1
XANTENNA__8118__B1 _8117_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5775_ _5741_/A _7316_/A _8194_/A _5744_/X vssd1 vssd1 vccd1 vccd1 _6744_/B sky130_fd_sc_hd__a22o_1
XANTENNA__6392__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7514_ _7514_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7514_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8669__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4726_ _4833_/B _4692_/Y _4833_/A vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8494_ _8494_/A vssd1 vssd1 vccd1 vccd1 _8494_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7445_ _7590_/A _7444_/A _7372_/A _6629_/Y vssd1 vssd1 vccd1 vccd1 _7445_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4657_ _4481_/B _5237_/A _4566_/A _5359_/B _4656_/X vssd1 vssd1 vccd1 vccd1 _4657_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6868__A _6868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput80 mports_i[171] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput91 mports_i[181] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_4
X_7376_ _7590_/A _7376_/B vssd1 vssd1 vccd1 vccd1 _7376_/Y sky130_fd_sc_hd__nor2_1
X_4588_ _7510_/A vssd1 vssd1 vccd1 vccd1 _7309_/B sky130_fd_sc_hd__inv_4
XFILLER_0_141_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6327_ _6324_/X _6326_/X _6386_/S vssd1 vssd1 vccd1 vccd1 _6327_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6896__B1_N _6895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6258_ _6252_/X _6234_/B _7246_/A _5128_/A _6386_/S vssd1 vssd1 vccd1 vccd1 _6258_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7644__A2 _6058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5209_ _5206_/X _6551_/A _6386_/S vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__mux2_1
X_6189_ _6628_/B _6186_/X _6188_/Y vssd1 vssd1 vccd1 vccd1 _6189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5407__A1 _7450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6604__B1 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7801__C1 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6108__A _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5947__A _6002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8323__A _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6907__A1 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5666__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4918__B1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4570__B _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6383__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5682__A _6727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6497__B _6497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5894__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5894__B2 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7096__B1 _7095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8832__A1 _8230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5646__A1 _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7399__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7121__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output406_A _7974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5857__A _6811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4480__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7571__A1 _6770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7571__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5560_ _5560_/A vssd1 vssd1 vccd1 vccd1 _5560_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5582__B1 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4511_ _4511_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5491_ input99/X _5192_/A input37/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5491_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6126__A2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7230_ _7229_/X _6185_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7231_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_151_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4442_ hold10/X vssd1 vssd1 vccd1 vccd1 _4760_/A sky130_fd_sc_hd__inv_2
XANTENNA__5334__B1 _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5885__A1 _5871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5885__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7161_ _7161_/A vssd1 vssd1 vccd1 vccd1 _7161_/X sky130_fd_sc_hd__buf_1
XFILLER_0_22_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ _8936_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6212_/A _6112_/B vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__or2_1
XANTENNA__8823__A1 _8203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7626__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7091_/X _6611_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7093_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5637__A1 _5637_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6834__B1 _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6043_ _8189_/A _6017_/B _6042_/X vssd1 vssd1 vccd1 vccd1 _7632_/B sky130_fd_sc_hd__o21ai_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4936__A _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6627__S _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7312__A _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4655__B _8845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8051__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7994_ _7989_/Y _6513_/A _7990_/Y _6080_/A _7993_/Y vssd1 vssd1 vccd1 vccd1 _8403_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6062__A1 _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6062__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6234_/A _6994_/B _6944_/Y _6989_/B vssd1 vssd1 vccd1 vccd1 _6945_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_135_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5767__A _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8143__A _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6876_ _6876_/A _6876_/B _6876_/C vssd1 vssd1 vccd1 vccd1 _6876_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8615_ _8614_/X _7886_/Y _8686_/B vssd1 vssd1 vccd1 vccd1 _8616_/A sky130_fd_sc_hd__mux2_1
X_5827_ _5827_/A _5827_/B vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7562__A1 _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8546_ _8584_/A _8175_/Y _8211_/Y _8261_/A _8545_/Y vssd1 vssd1 vccd1 vccd1 _8547_/A
+ sky130_fd_sc_hd__a221o_1
X_5758_ _6758_/B _5077_/A _6017_/A _5803_/A vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__a22o_1
XANTENNA__5573__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4709_ hold45/A _4894_/A _7272_/B vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__nor3_1
X_8477_ _8476_/Y _8451_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8477_/X sky130_fd_sc_hd__mux2_1
X_5689_ _6024_/A _6737_/A vssd1 vssd1 vccd1 vccd1 _5689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5325__B1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7428_ _7590_/A _7428_/B vssd1 vssd1 vccd1 vccd1 _7428_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7359_ _7359_/A vssd1 vssd1 vccd1 vccd1 _7619_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__6110__B _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5007__A _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8814__A1 _8137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7222__A _7222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4565__B _7707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8042__A2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7553__A1 _5765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5619__A1 _5659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5619__B2 _7524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8281__A2 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6292__A1 _6315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6292__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput270 sports_i[13] vssd1 vssd1 vccd1 vccd1 _7962_/A sky130_fd_sc_hd__buf_1
Xinput281 sports_i[23] vssd1 vssd1 vccd1 vccd1 _8098_/A sky130_fd_sc_hd__buf_1
Xinput292 sports_i[33] vssd1 vssd1 vccd1 vccd1 _8251_/A2 sky130_fd_sc_hd__buf_2
XANTENNA__6971__A _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8033__A2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7241__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4991_ _4978_/B _8716_/B _4977_/B _4917_/X vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6730_ _5625_/A _7536_/B _7707_/B _6732_/A vssd1 vssd1 vccd1 vccd1 _6731_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_129_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6661_ _6637_/Y _6660_/X _6870_/S vssd1 vssd1 vccd1 vccd1 _6662_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6347__A2 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8400_ _8400_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8400_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5612_ _6470_/B _5609_/Y _7498_/A vssd1 vssd1 vccd1 vccd1 _5613_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6592_ _6590_/X _6591_/X _6694_/B _5280_/A _6475_/X vssd1 vssd1 vccd1 vccd1 _6592_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8972__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8331_ _8564_/B _7906_/Y _8349_/A vssd1 vssd1 vccd1 vccd1 _8331_/X sky130_fd_sc_hd__o21a_1
X_5543_ _5543_/A1 _5192_/A input39/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5543_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_42_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7307__A _7347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8262_ _8255_/X _8260_/X _8567_/B vssd1 vssd1 vccd1 vccd1 _8262_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5307__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5474_ _5697_/A1 _8709_/B input46/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5474_/X sky130_fd_sc_hd__o22a_1
Xoutput700 _6640_/Y vssd1 vssd1 vccd1 vccd1 sports_o[73] sky130_fd_sc_hd__buf_12
XANTENNA__5858__A1 _5928_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput711 _6735_/X vssd1 vssd1 vccd1 vccd1 sports_o[83] sky130_fd_sc_hd__buf_12
X_7213_ _7213_/A vssd1 vssd1 vccd1 vccd1 _7213_/X sky130_fd_sc_hd__buf_1
Xoutput722 _6863_/X vssd1 vssd1 vccd1 vccd1 sports_o[93] sky130_fd_sc_hd__buf_12
XANTENNA__5858__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4425_ _4425_/A _4425_/B _4425_/C vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_100_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8193_ _8193_/A vssd1 vssd1 vccd1 vccd1 _8193_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7741__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4530__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7144_ _7524_/A _7004_/X _5600_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7144_/X
+ sky130_fd_sc_hd__a221o_1
X_4356_ _4684_/A _4684_/B hold46/A vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_10_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7075_ _6578_/B _7059_/X _5292_/A _7246_/B _7061_/X vssd1 vssd1 vccd1 vccd1 _7075_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5261__S _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8138__A _8150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7042__A _7042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5086__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6026_ _5972_/X _7638_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6026_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4385__B _7304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8572__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8024__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7696__B _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7977_ _7977_/A vssd1 vssd1 vccd1 vccd1 _7977_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7783__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7783__B2 _7790_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5794__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6928_ _6928_/A vssd1 vssd1 vccd1 vccd1 _6928_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6859_ _6859_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_147_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8732__B1 _7811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8529_ _8145_/Y _8304_/X _8148_/X _8299_/X _8496_/S vssd1 vssd1 vccd1 vccd1 _8529_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7217__A _7217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7838__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8747__S _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5960__A _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8263__A2 _8215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6274__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7471__B1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4295__B _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7223__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8420__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8511__A _8511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8487__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6501__A2 _6543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5870__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ _6526_/A _5845_/B vssd1 vssd1 vccd1 vccd1 _5190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6177__S _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8254__A2 _8244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4486__A _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk_i clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk_i/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__6265__A1 _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5068__A2 _7341_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7462__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7900_ _7905_/A1 _5146_/A _7905_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _7900_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__8006__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8880_ _8880_/A vssd1 vssd1 vccd1 vccd1 _8880_/Y sky130_fd_sc_hd__inv_2
X_7831_ _7827_/Y _5146_/A _7828_/Y _7431_/B _7830_/X vssd1 vssd1 vccd1 vccd1 _7832_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7765__A1 _4318_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7765__B2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4974_ _4974_/A vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__inv_2
X_7762_ _7761_/Y _5117_/A _4331_/B _7779_/B1 _7761_/A vssd1 vssd1 vccd1 vccd1 _7762_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6713_ _6713_/A _6899_/B vssd1 vssd1 vccd1 vccd1 _6713_/X sky130_fd_sc_hd__and2_1
XFILLER_0_129_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7693_ _6189_/Y _7359_/A _7689_/X _7691_/Y _7692_/Y vssd1 vssd1 vccd1 vccd1 _7693_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5528__B1 _5527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6644_ _6644_/A vssd1 vssd1 vccd1 vccd1 _6644_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_34_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8190__B2 hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6575_ _7767_/A _7829_/A _8185_/B _5283_/Y vssd1 vssd1 vccd1 vccd1 _6575_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8140__B _8151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6740__A2 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7037__A _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8314_ _8309_/X _8304_/A _8313_/X _8299_/A vssd1 vssd1 vccd1 vccd1 _8314_/X sky130_fd_sc_hd__a22o_1
X_5526_ _5526_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _5526_/X sky130_fd_sc_hd__and2_1
XFILLER_0_143_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8245_ _5185_/A _8252_/B1 _6500_/A _8251_/B2 vssd1 vssd1 vccd1 vccd1 _8245_/X sky130_fd_sc_hd__a22o_1
X_5457_ _5401_/A _5102_/A _5402_/A _5191_/A _5456_/X vssd1 vssd1 vccd1 vccd1 _7459_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_2_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput530 _7410_/X vssd1 vssd1 vccd1 vccd1 sports_o[125] sky130_fd_sc_hd__buf_12
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5780__A _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput541 _7493_/X vssd1 vssd1 vccd1 vccd1 sports_o[135] sky130_fd_sc_hd__buf_12
XFILLER_0_140_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput552 _7582_/X vssd1 vssd1 vccd1 vccd1 sports_o[145] sky130_fd_sc_hd__buf_12
X_4408_ _4408_/A _4408_/B vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__nand2_1
Xoutput563 _7677_/X vssd1 vssd1 vccd1 vccd1 sports_o[155] sky130_fd_sc_hd__buf_12
XANTENNA__5700__B1 _5686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8176_ _8175_/Y _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _8176_/Y sky130_fd_sc_hd__a21oi_1
X_5388_ _5385_/Y _4885_/A _5386_/Y _4891_/A _5387_/Y vssd1 vssd1 vccd1 vccd1 _5425_/C
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput574 _7734_/Y vssd1 vssd1 vccd1 vccd1 sports_o[165] sky130_fd_sc_hd__buf_12
XFILLER_0_10_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput585 _5068_/X vssd1 vssd1 vccd1 vccd1 sports_o[175] sky130_fd_sc_hd__buf_12
Xoutput596 _5399_/X vssd1 vssd1 vccd1 vccd1 sports_o[185] sky130_fd_sc_hd__buf_12
X_7127_ _5558_/X _7023_/X _7126_/X vssd1 vssd1 vccd1 vccd1 _7127_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8245__A2 _8252_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4339_ _4338_/Y _4337_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__6256__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7058_ _7058_/A vssd1 vssd1 vccd1 vccd1 _7058_/X sky130_fd_sc_hd__buf_1
X_6009_ _6128_/B _6868_/A _5136_/X vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6008__A1 _5931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6008__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6116__A _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5020__A _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4990__A1 _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6716__C1 _6715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8477__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8961__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6786__A _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8236__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6247__A1 _6247_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6247__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7995__A1 _7998_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7995__B2 _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__B1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output688_A _6493_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6970__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4690_ _4690_/A vssd1 vssd1 vccd1 vccd1 _4833_/B sky130_fd_sc_hd__inv_2
XFILLER_0_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6722__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6360_ _6360_/A vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__buf_1
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5311_ _5845_/B _7413_/A _5310_/Y _6133_/B vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__a22o_1
X_6291_ _6224_/S _7720_/B _6288_/X _6290_/Y vssd1 vssd1 vccd1 vccd1 _6291_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6486__A1 _7341_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8030_ _8030_/A vssd1 vssd1 vccd1 vccd1 _8030_/Y sky130_fd_sc_hd__inv_2
X_5242_ _8151_/B vssd1 vssd1 vccd1 vccd1 _7707_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__5694__C1 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7304__B _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8227__A2 _8235_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5173_ _5163_/X _6590_/B _6780_/A vssd1 vssd1 vccd1 vccd1 _6557_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6238__A1 _6247_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5105__A _5105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6238__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8778__A3 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7986__B2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 mports_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
X_8932_ _4848_/A _4847_/A hold10/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4944__A _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8416__A _8416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8863_ _8857_/A _6059_/B _6264_/X _4618_/A vssd1 vssd1 vccd1 vccd1 _8863_/X sky130_fd_sc_hd__a211o_1
XANTENNA__7738__A1 _7736_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7814_ _7814_/A1 _5230_/B _7814_/B1 _5197_/X _7813_/X vssd1 vssd1 vccd1 vccd1 _8284_/B
+ sky130_fd_sc_hd__a221oi_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8794_ _8793_/X _8081_/Y _8824_/S vssd1 vssd1 vccd1 vccd1 _8794_/X sky130_fd_sc_hd__mux2_1
X_4957_ _4957_/A vssd1 vssd1 vccd1 vccd1 _4957_/Y sky130_fd_sc_hd__inv_2
X_7745_ _6364_/X _7754_/A _7743_/Y _7744_/X vssd1 vssd1 vccd1 vccd1 _7745_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6961__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8151__A _8151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4888_ _4888_/A vssd1 vssd1 vccd1 vccd1 _4888_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7676_ _7683_/B _7674_/X _6928_/Y _7359_/A vssd1 vssd1 vccd1 vccd1 _7676_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6174__B1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6627_ _5367_/Y _6626_/Y _8924_/B vssd1 vssd1 vccd1 vccd1 _6628_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_144_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6558_ _6852_/A _6558_/B vssd1 vssd1 vccd1 vccd1 _6558_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5509_ _6080_/A _5549_/A vssd1 vssd1 vccd1 vccd1 _5509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_131_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6489_ _6489_/A vssd1 vssd1 vccd1 vccd1 _7043_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7674__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8228_ _6500_/A _8234_/B2 _8234_/A2 _7769_/A vssd1 vssd1 vccd1 vccd1 _8229_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_30_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput371 _8730_/X vssd1 vssd1 vccd1 vccd1 mports_o[104] sky130_fd_sc_hd__buf_12
Xoutput382 _8766_/X vssd1 vssd1 vccd1 vccd1 mports_o[114] sky130_fd_sc_hd__buf_12
XFILLER_0_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput393 _8799_/X vssd1 vssd1 vccd1 vccd1 mports_o[124] sky130_fd_sc_hd__buf_12
XANTENNA__8218__A2 _8222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8159_ _8160_/A _8171_/B vssd1 vssd1 vccd1 vccd1 _8159_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6229__A1 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6229__B2 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7426__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6545__S _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6401__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5685__A _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4963__A1 _4956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4963__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8154__A1 _8153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6704__A2 _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7901__B2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6468__B2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8209__A2 _8209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7417__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7968__A1 _7971_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7968__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8090__B1 _8093_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5443__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5579__B _6695_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5860_ _5860_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _5860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _8875_/A _4811_/B vssd1 vssd1 vccd1 vccd1 _8869_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5791_ _6770_/A _7536_/B _7707_/B _6788_/B vssd1 vssd1 vccd1 vccd1 _5791_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_145_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6943__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5595__A _5609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4954__A1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4742_ hold32/X _8578_/B vssd1 vssd1 vccd1 vccd1 _8919_/A sky130_fd_sc_hd__nor2_8
X_7530_ _7683_/B _7528_/B _7527_/X _7528_/X _7529_/Y vssd1 vssd1 vccd1 vccd1 _7530_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4954__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7461_ _7458_/X _7723_/B _7460_/Y vssd1 vssd1 vccd1 vccd1 _7461_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4673_ _4673_/A _4675_/A vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6203__B _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6412_ _6513_/A _8755_/C vssd1 vssd1 vccd1 vccd1 _6724_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5903__B1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7392_ _7590_/A _7379_/Y _7380_/Y _7391_/X vssd1 vssd1 vccd1 vccd1 _7392_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_3_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6343_ _7272_/B _5128_/A _6342_/A _5845_/B _6386_/S vssd1 vssd1 vccd1 vccd1 _6343_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4939__A _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7315__A _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6459__B2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6274_ _6287_/A1 _5080_/A input7/X _4870_/X _6273_/X vssd1 vssd1 vccd1 vccd1 _6283_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__4658__B _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5131__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5225_ input93/X _8271_/B input30/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__o22a_1
X_8013_ _7777_/X _8012_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _8013_/X sky130_fd_sc_hd__o21ba_1
X_5156_ _5195_/A1 _5111_/A _5195_/B1 _4931_/A _5155_/X vssd1 vssd1 vccd1 vccd1 _5159_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_99_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7959__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8620__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8146__A _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5087_ _6489_/A _5185_/A vssd1 vssd1 vccd1 vccd1 _5087_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6631__A1 _7451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6631__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8915_ _4425_/A _6470_/B _8917_/S vssd1 vssd1 vccd1 vccd1 _8916_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8846_ _8846_/A _8846_/B vssd1 vssd1 vccd1 vccd1 _8847_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8384__A1 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8384__B2 _7942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8777_ _8009_/Y _8711_/A _8824_/S vssd1 vssd1 vccd1 vccd1 _8777_/X sky130_fd_sc_hd__a21o_1
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A vssd1 vssd1 vccd1 vccd1 _5989_/Y sky130_fd_sc_hd__inv_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6934__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7728_ _6326_/X _7723_/B _7727_/X vssd1 vssd1 vccd1 vccd1 _7728_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8136__A1 _8151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8136__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7209__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6147__B1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8687__A2 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7659_ _6897_/Y _7668_/B _6082_/X _7638_/B vssd1 vssd1 vccd1 vccd1 _7659_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_133_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6698__A1 _5535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8966__D _8966_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7647__B1 _7643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7111__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8611__A2 _7878_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7178__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8503__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7583__C1 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8127__A1 _8132_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6304__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8127__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6138__B1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8678__A2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7834__S _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7350__A2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6958__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5862__B _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4478__B _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A1 _5070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _6469_/B _5174_/A vssd1 vssd1 vccd1 vccd1 _5010_/Y sky130_fd_sc_hd__nand2_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5664__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8602__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5416__A2 _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7810__B1 _7813_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6961_ _6283_/A _6994_/B _6272_/X _6989_/B vssd1 vssd1 vccd1 vccd1 _6961_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8700_ _4607_/A _8685_/B _8686_/B vssd1 vssd1 vccd1 vccd1 _8700_/Y sky130_fd_sc_hd__a21oi_1
X_5912_ _6841_/B _6544_/B vssd1 vssd1 vccd1 vccd1 _5948_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8366__A1 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6892_ _7707_/B _6892_/B vssd1 vssd1 vccd1 vccd1 _6892_/X sky130_fd_sc_hd__or2_1
XANTENNA__8366__B2 _7932_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8631_ _8698_/B _8765_/B _8590_/X vssd1 vssd1 vccd1 vccd1 _8631_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6377__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5843_ _6547_/A _5839_/X _5842_/Y vssd1 vssd1 vccd1 vccd1 _7584_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6916__A2 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8562_ _8564_/B _8235_/Y _8349_/A vssd1 vssd1 vccd1 vccd1 _8562_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8118__A1 _8510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5774_ _5774_/A vssd1 vssd1 vccd1 vccd1 _6802_/A sky130_fd_sc_hd__inv_2
XFILLER_0_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8118__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7513_ _5659_/A _7542_/A _7694_/A _5620_/X vssd1 vssd1 vccd1 vccd1 _7513_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8669__A2 _8107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4725_ _4725_/A _4725_/B vssd1 vssd1 vccd1 vccd1 _4833_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_72_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6129__B1 _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8493_ _8440_/X _8492_/X _8759_/B vssd1 vssd1 vccd1 vccd1 _8494_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_115_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7877__B1 _7877_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4656_ _5359_/A _4478_/B _5116_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4656_/X sky130_fd_sc_hd__a22o_1
X_7444_ _7444_/A _7691_/B vssd1 vssd1 vccd1 vccd1 _7444_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6868__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput70 mports_i[162] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_2
XFILLER_0_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput81 mports_i[172] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_2
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4587_ _4607_/A _5230_/B _4607_/B _4557_/B vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__a31o_1
X_7375_ _7701_/A vssd1 vssd1 vccd1 vccd1 _7590_/A sky130_fd_sc_hd__buf_8
Xinput92 mports_i[182] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_2
XFILLER_0_40_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6326_ _6326_/A1 _8516_/B input9/X _4913_/X _6325_/X vssd1 vssd1 vccd1 vccd1 _6326_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5104__A1 _5139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5104__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6257_ _6257_/A vssd1 vssd1 vccd1 vccd1 _7246_/A sky130_fd_sc_hd__inv_2
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6301__B1 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5208_ _5208_/A1 _8271_/A _5208_/B1 _5191_/X _5207_/X vssd1 vssd1 vccd1 vccd1 _6551_/A
+ sky130_fd_sc_hd__o221a_4
X_6188_ _6628_/B _6188_/B vssd1 vssd1 vccd1 vccd1 _6188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5139_ _5139_/A vssd1 vssd1 vccd1 vccd1 _5139_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6604__A1 _5356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7801__B1 _7800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8357__A1 _8376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5947__B _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6368__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8829_ _8828_/X _8215_/X _8829_/S vssd1 vssd1 vccd1 vccd1 _8830_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_137_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4918__A1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5666__C _5666_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4918__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8109__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4570__C _7707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7868__B1 _7877_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5682__B _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5894__A2 _5853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4298__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7096__A1 _6622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8293__B1 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7399__A2 _6567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7571__A2 _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4510_ _4510_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _4511_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5490_ _5490_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _5490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4441_ _7510_/A hold1/X vssd1 vssd1 vccd1 vccd1 _8942_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5334__A1 _5011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5885__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7160_ _7159_/X _5744_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7161_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4372_ _4372_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4373_/B sky130_fd_sc_hd__nor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6689_/S _6103_/X _6110_/Y vssd1 vssd1 vccd1 vccd1 _7673_/B sky130_fd_sc_hd__o21ai_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8395__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7091_ _5317_/A _7023_/X _7090_/X vssd1 vssd1 vccd1 vccd1 _7091_/X sky130_fd_sc_hd__o21a_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6042_ _6281_/S _6042_/B vssd1 vssd1 vccd1 vccd1 _6042_/X sky130_fd_sc_hd__or2_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6834__A1 _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7312__B _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7993_ _7998_/A1 _5146_/A _7998_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _7993_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__6062__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6643__S _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6944_ _6944_/A vssd1 vssd1 vccd1 vccd1 _6944_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8424__A _8424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8339__A1 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4671__B _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6875_ _7632_/B _6875_/B vssd1 vssd1 vccd1 vccd1 _6876_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8614_ _8613_/X _8334_/A _8621_/S vssd1 vssd1 vccd1 vccd1 _8614_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5826_ _5809_/A _4953_/A _5810_/A _5089_/A _5825_/X vssd1 vssd1 vccd1 vccd1 _5827_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8545_ _8133_/Y _8336_/S _8364_/Y vssd1 vssd1 vccd1 vccd1 _8545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5573__A1 _5552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5757_ _5788_/A1 _4868_/A _5788_/B1 _5089_/A _5756_/X vssd1 vssd1 vccd1 vccd1 _5803_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_45_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5573__B2 _5659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5783__A _6756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4708_ _8512_/S hold41/A vssd1 vssd1 vccd1 vccd1 _4894_/A sky130_fd_sc_hd__nand2_4
X_8476_ _8476_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8476_/Y sky130_fd_sc_hd__nand2_1
X_5688_ _5685_/Y _4890_/A _5686_/Y _4885_/A _5687_/Y vssd1 vssd1 vccd1 vccd1 _6737_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6598__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5325__A1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7427_ _7428_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7427_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5325__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4639_ hold30/A _8875_/B vssd1 vssd1 vccd1 vccd1 _8264_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7358_ _7372_/A vssd1 vssd1 vccd1 vccd1 _7359_/A sky130_fd_sc_hd__inv_2
XFILLER_0_102_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6309_ _6309_/A1 _8716_/B input71/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6309_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8275__B1 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8814__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7289_ _6385_/A _7138_/A _7287_/X _7288_/X vssd1 vssd1 vccd1 vccd1 _7289_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6825__A1 _5930_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6825__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5958__A _6059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8334__A _8334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5564__A1 _5591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5564__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8805__A2 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7413__A _7413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5619__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4756__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6292__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput260 sports_i[127] vssd1 vssd1 vccd1 vccd1 _8132_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__6029__A _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output516_A _6998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8569__A1 _4661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput271 sports_i[14] vssd1 vssd1 vccd1 vccd1 _7977_/A sky130_fd_sc_hd__buf_1
Xinput282 sports_i[24] vssd1 vssd1 vccd1 vccd1 _8110_/A sky130_fd_sc_hd__buf_1
Xinput293 sports_i[34] vssd1 vssd1 vccd1 vccd1 _4331_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6971__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7241__A1 _6241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4990_ _8578_/B _5185_/A _4973_/Y _4989_/X vssd1 vssd1 vccd1 vccd1 _4990_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6660_ _6658_/Y _6659_/Y _8150_/A vssd1 vssd1 vccd1 vccd1 _6660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8741__A1 _7862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5611_ _5611_/A vssd1 vssd1 vccd1 vccd1 _7498_/A sky130_fd_sc_hd__inv_2
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5555__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6591_ _6837_/A _6591_/B vssd1 vssd1 vccd1 vccd1 _6591_/X sky130_fd_sc_hd__or2_1
XANTENNA__5555__B2 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6752__B1 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8330_ _7901_/Y _8304_/X _7903_/Y _8299_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8330_/X
+ sky130_fd_sc_hd__a221o_1
X_5542_ _5536_/X _5541_/X _6170_/A vssd1 vssd1 vccd1 vccd1 _5542_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5307__A1 _7422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5473_ _5596_/A _5080_/A _5597_/A _5089_/X _5472_/X vssd1 vssd1 vccd1 vccd1 _7524_/A
+ sky130_fd_sc_hd__o221a_4
X_8261_ _8261_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _8567_/B sky130_fd_sc_hd__nand2_8
XANTENNA__5307__B2 _5094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6211__B _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput701 _6652_/X vssd1 vssd1 vccd1 vccd1 sports_o[74] sky130_fd_sc_hd__buf_12
Xoutput712 _6742_/X vssd1 vssd1 vccd1 vccd1 sports_o[84] sky130_fd_sc_hd__buf_12
XANTENNA__5108__A _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5858__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7212_ _7211_/X _6095_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7213_/A sky130_fd_sc_hd__mux2_2
X_4424_ _4424_/A _6312_/A vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__nand2_1
Xoutput723 _6874_/X vssd1 vssd1 vccd1 vccd1 sports_o[94] sky130_fd_sc_hd__buf_12
XFILLER_0_111_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8192_ _8192_/A _8194_/A vssd1 vssd1 vccd1 vccd1 _8193_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7143_ _7143_/A vssd1 vssd1 vccd1 vccd1 _7143_/X sky130_fd_sc_hd__buf_1
X_4355_ hold45/X _5485_/A vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__nor2_1
XANTENNA__4947__A _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7074_ _7074_/A vssd1 vssd1 vccd1 vccd1 _7074_/X sky130_fd_sc_hd__buf_1
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6025_ _5992_/Y _6051_/A _8160_/A vssd1 vssd1 vccd1 vccd1 _7638_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7480__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7232__A1 _6221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7232__B2 _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7976_ _7976_/A vssd1 vssd1 vccd1 vccd1 _7976_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7783__A2 _7790_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5794__A1 _5765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6927_ _6906_/A _6188_/B _6926_/X vssd1 vssd1 vccd1 vccd1 _6928_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5794__B2 _6771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6858_ _6858_/A vssd1 vssd1 vccd1 vccd1 _6859_/A sky130_fd_sc_hd__inv_2
XANTENNA__8732__A1 _7809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5809_ _5809_/A vssd1 vssd1 vccd1 vccd1 _5809_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5546__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6789_ _6818_/A _6765_/A _6906_/A vssd1 vssd1 vccd1 vccd1 _6789_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6402__A _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8528_ _8323_/X _8525_/Y _8526_/X _8527_/X vssd1 vssd1 vccd1 vccd1 _8528_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8459_ _8458_/Y _8423_/Y _8481_/S vssd1 vssd1 vccd1 vccd1 _8460_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5018__A _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8248__B1 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8799__A1 _8490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6274__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7471__B2 _7469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7223__A1 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5785__A1 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5785__B2 _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8511__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6312__A _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8239__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6265__A2 _6263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7462__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7214__A1 _7660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6193__S _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7830_ _7829_/Y _4328_/B _8185_/B vssd1 vssd1 vccd1 vccd1 _7830_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7214__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5225__B1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7765__A2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7761_ _7761_/A _7778_/B vssd1 vssd1 vccd1 vccd1 _7761_/Y sky130_fd_sc_hd__nand2_1
X_4973_ _5022_/B _6017_/A vssd1 vssd1 vccd1 vccd1 _4973_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6712_ _7514_/A _6475_/A _6711_/X _6694_/B vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7692_ _7701_/A _7692_/B vssd1 vssd1 vccd1 vccd1 _7692_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_132_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5528__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6643_ _5353_/A _6642_/Y _6870_/S vssd1 vssd1 vccd1 vccd1 _6643_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8190__A2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6574_ _6547_/A _5253_/X _6573_/X vssd1 vssd1 vccd1 vccd1 _7394_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8313_ _4870_/X _7856_/Y _4874_/X _7811_/X _8312_/X vssd1 vssd1 vccd1 vccd1 _8313_/X
+ sky130_fd_sc_hd__o221a_2
X_5525_ _5909_/B _7115_/A _5524_/Y _5997_/B vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8244_ _8251_/B2 _8857_/B _8252_/B1 _5359_/B _8243_/X vssd1 vssd1 vccd1 vccd1 _8244_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5456_ input98/X _5192_/A input36/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5456_/X sky130_fd_sc_hd__o22a_1
Xoutput520 _7333_/Y vssd1 vssd1 vccd1 vccd1 sports_o[116] sky130_fd_sc_hd__buf_12
XFILLER_0_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput531 _7420_/X vssd1 vssd1 vccd1 vccd1 sports_o[126] sky130_fd_sc_hd__buf_12
Xoutput542 _7502_/Y vssd1 vssd1 vccd1 vccd1 sports_o[136] sky130_fd_sc_hd__buf_12
XFILLER_0_100_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4407_ _4415_/A _4425_/B _4407_/C vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__nand3_1
Xoutput553 _7591_/X vssd1 vssd1 vccd1 vccd1 sports_o[146] sky130_fd_sc_hd__buf_12
XANTENNA__5700__A1 _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8175_ _8175_/A1 _6102_/B _8171_/Y _8173_/Y _8174_/Y vssd1 vssd1 vccd1 vccd1 _8175_/Y
+ sky130_fd_sc_hd__o221ai_4
Xoutput564 _7684_/X vssd1 vssd1 vccd1 vccd1 sports_o[156] sky130_fd_sc_hd__buf_12
X_5387_ _5274_/X input97/X _5275_/X input35/X vssd1 vssd1 vccd1 vccd1 _5387_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__5700__B2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput575 _7738_/Y vssd1 vssd1 vccd1 vccd1 sports_o[166] sky130_fd_sc_hd__buf_12
XFILLER_0_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput586 _5127_/X vssd1 vssd1 vccd1 vccd1 sports_o[176] sky130_fd_sc_hd__buf_12
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput597 _5414_/X vssd1 vssd1 vccd1 vccd1 sports_o[186] sky130_fd_sc_hd__buf_12
XFILLER_0_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ _5500_/X _7004_/X _5549_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7126_/X
+ sky130_fd_sc_hd__a221o_1
X_4338_ _4338_/A _4338_/B vssd1 vssd1 vccd1 vccd1 _4338_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6256__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7453__A1 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7057_ _7056_/X _7356_/B _7097_/S vssd1 vssd1 vccd1 vccd1 _7058_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6892__A _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5464__B1 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6008_ _5931_/A _8335_/B _5932_/A _4913_/A _6007_/X vssd1 vssd1 vccd1 vccd1 _6868_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__7199__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6008__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7205__A1 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7205__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5216__B1 _5222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5301__A _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7948_/Y _7874_/X _7949_/Y _7875_/X _7958_/Y vssd1 vssd1 vccd1 vccd1 _8765_/B
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_38_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8705__A1 _8244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7508__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4990__A2 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5690__B _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6247__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8493__S _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7995__A2 _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5207__B1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7747__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5211__A _5211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__A1 _6758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__B2 _5803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6955__B1 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7904__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7138__A _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6183__A1 _6183_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6042__A _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7572__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5310_ _5310_/A vssd1 vssd1 vccd1 vccd1 _5310_/Y sky130_fd_sc_hd__inv_2
X_6290_ _6290_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6290_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5241_ _6059_/B _6567_/A _5329_/A _8924_/B vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4497__A _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5172_ _6166_/B vssd1 vssd1 vccd1 vccd1 _6780_/A sky130_fd_sc_hd__buf_6
XANTENNA__6238__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5446__A0 _7450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7986__A2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 mports_i[100] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_8931_ hold8/X _8931_/B vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__nand2_1
XANTENNA__4944__B _7372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8416__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8862_ _8855_/A _8861_/Y _4618_/A vssd1 vssd1 vccd1 vccd1 _8862_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6217__A _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7738__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7813_ _7874_/A _7813_/A2 _8174_/A _7813_/B2 vssd1 vssd1 vccd1 vccd1 _7813_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8793_ _8483_/A _8738_/A _8480_/A _8711_/A vssd1 vssd1 vccd1 vccd1 _8793_/X sky130_fd_sc_hd__a22o_1
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7744_ _7349_/Y _6367_/B _7326_/A vssd1 vssd1 vccd1 vccd1 _7744_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4960__A _4960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4956_ _4956_/A vssd1 vssd1 vccd1 vccd1 _4956_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8699__B1 _8226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8151__B _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7675_ _6102_/A _7681_/A _7606_/A _7674_/X vssd1 vssd1 vccd1 vccd1 _7675_/X sky130_fd_sc_hd__o22a_1
X_4887_ _8455_/B vssd1 vssd1 vccd1 vccd1 _8550_/B sky130_fd_sc_hd__buf_8
XFILLER_0_117_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6174__A1 _6174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6626_ _6630_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _6626_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6174__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7371__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5921__A1 _6007_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6557_ _6557_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6557_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5921__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5508_ _5505_/Y _4886_/A _5506_/Y _4891_/A _5507_/Y vssd1 vssd1 vccd1 vccd1 _5549_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6488_ _6488_/A _6488_/B vssd1 vssd1 vccd1 vccd1 _6488_/Y sky130_fd_sc_hd__nand2_1
X_8227_ _5185_/A _8235_/B1 _8235_/A1 _7299_/A vssd1 vssd1 vccd1 vccd1 _8229_/A sky130_fd_sc_hd__a22o_1
XANTENNA__7674__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5439_ _6079_/A _6669_/B vssd1 vssd1 vccd1 vccd1 _5537_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput372 _8734_/X vssd1 vssd1 vccd1 vccd1 mports_o[105] sky130_fd_sc_hd__buf_12
Xoutput383 _8769_/X vssd1 vssd1 vccd1 vccd1 mports_o[115] sky130_fd_sc_hd__buf_12
Xoutput394 _8802_/X vssd1 vssd1 vccd1 vccd1 mports_o[125] sky130_fd_sc_hd__buf_12
X_8158_ _8158_/A vssd1 vssd1 vccd1 vccd1 _8171_/B sky130_fd_sc_hd__inv_2
XANTENNA__6229__A2 _6229_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7426__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7109_ _7109_/A vssd1 vssd1 vccd1 vccd1 _7109_/X sky130_fd_sc_hd__buf_1
X_8089_ _8084_/Y _6513_/A _8085_/Y _6080_/A _8088_/Y vssd1 vssd1 vccd1 vccd1 _8511_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5437__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4660__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6401__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4870__A _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4963__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8154__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6165__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7901__A2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6468__A2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5676__B1 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7417__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5428__B1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7968__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8090__A1 _8093_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8090__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6640__A2 _6511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8917__A1 _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ _4810_/A _4810_/B vssd1 vssd1 vccd1 vccd1 _4811_/B sky130_fd_sc_hd__nand2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _5809_/A _8271_/A _5810_/A _5191_/X _5789_/X vssd1 vssd1 vccd1 vccd1 _6788_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_118_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4741_ _8240_/A _6980_/B _4740_/Y _4738_/B vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__a31o_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4954__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7460_ _7673_/A _6662_/A _7459_/Y vssd1 vssd1 vccd1 vccd1 _7460_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4672_ _4672_/A _4674_/A vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6411_ _6411_/A vssd1 vssd1 vccd1 vccd1 _6513_/A sky130_fd_sc_hd__buf_12
XANTENNA__5903__A1 _5871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7391_ _6565_/A _7361_/X _7388_/Y _7754_/A _7390_/X vssd1 vssd1 vccd1 vccd1 _7391_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5903__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5815__S _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6500__A _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6342_ _6342_/A _8578_/B _8188_/S hold23/A vssd1 vssd1 vccd1 vccd1 _6342_/X sky130_fd_sc_hd__and4_1
XFILLER_0_141_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7315__B _7683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6273_ _6286_/A1 _8310_/B input70/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6273_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8853__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4658__C _8845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8012_ _8002_/Y _7874_/X _8003_/Y _7875_/X _8011_/Y vssd1 vssd1 vccd1 vccd1 _8012_/Y
+ sky130_fd_sc_hd__a221oi_4
X_5224_ _5265_/A _5191_/X _5266_/A _8335_/B _5223_/X vssd1 vssd1 vccd1 vccd1 _5248_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5131__A2 _5131_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5155_ input88/X _4934_/A input26/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8427__A _8427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7331__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7959__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5086_ _5070_/A _5080_/A _5071_/A _4870_/X _5085_/X vssd1 vssd1 vccd1 vccd1 _6489_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__8081__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7050__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6631__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8914_ _8913_/A _4502_/A hold24/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8845_ _8845_/A _8845_/B _8845_/C vssd1 vssd1 vccd1 vccd1 _8848_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8384__A2 _7969_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8951__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8162__A _8162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8776_ _8400_/A _8806_/B _8774_/X _8775_/X vssd1 vssd1 vccd1 vccd1 _8776_/X sky130_fd_sc_hd__a22o_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5988_ _5988_/A vssd1 vssd1 vccd1 vccd1 _5988_/Y sky130_fd_sc_hd__inv_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7727_ _6317_/X _7349_/A _6971_/X _7753_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7727_/X
+ sky130_fd_sc_hd__a221o_1
X_4939_ _4939_/A vssd1 vssd1 vccd1 vccd1 _4940_/A sky130_fd_sc_hd__buf_6
XFILLER_0_136_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8136__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6147__A1 _6182_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7658_ _8574_/B _6095_/X _7654_/X _7656_/Y _7657_/Y vssd1 vssd1 vccd1 vccd1 _7658_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6147__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7895__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6609_ _6609_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6609_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6698__A2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7589_ _7590_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6410__A _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5696__A _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6304__B _6965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8127__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6138__A1 _6174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6138__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8532__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7886__A1 _7881_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7886__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5897__B1 _5937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8835__B1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A2 _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6310__A1 _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8063__B2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7810__A1 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7810__B2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6960_ _6263_/X _6429_/S _6958_/Y _6959_/X vssd1 vssd1 vccd1 vccd1 _6960_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5821__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8966__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5911_ _5936_/A _4870_/A _5937_/A _5080_/A _5910_/X vssd1 vssd1 vccd1 vccd1 _6841_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_76_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6891_ _6891_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6891_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8366__A2 _8765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8630_ _8358_/A _8581_/X _7956_/Y _8583_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8630_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6377__A1 _6387_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5842_ _5842_/A _6547_/A vssd1 vssd1 vccd1 vccd1 _5842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_124_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6377__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8561_ _8215_/X _8323_/X _8559_/X _8560_/X vssd1 vssd1 vccd1 vccd1 _8561_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5773_ _5770_/X _7316_/A _8194_/A _5772_/X vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8118__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7512_ _7512_/A vssd1 vssd1 vccd1 vccd1 _7536_/A sky130_fd_sc_hd__inv_2
X_4724_ _4732_/B _4731_/A vssd1 vssd1 vccd1 vccd1 _4725_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6129__A1 _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8492_ _8490_/Y _8491_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8492_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_133_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7877__A1 _7877_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7443_ _7701_/A _5367_/A _6264_/X vssd1 vssd1 vccd1 vccd1 _7444_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7877__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4655_ _8194_/A _8845_/C vssd1 vssd1 vccd1 vccd1 _5237_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_25_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7326__A _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5888__B1 _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput60 mports_i[153] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
Xinput71 mports_i[163] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_2
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7374_ _7376_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7374_/Y sky130_fd_sc_hd__nand2_1
Xinput82 mports_i[173] vssd1 vssd1 vccd1 vccd1 _4978_/B sky130_fd_sc_hd__buf_2
XFILLER_0_141_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4586_ _4586_/A _4793_/A vssd1 vssd1 vccd1 vccd1 _4607_/B sky130_fd_sc_hd__nor2_1
Xinput93 mports_i[183] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6325_ _6315_/B _8716_/B _6314_/B _4917_/X vssd1 vssd1 vccd1 vccd1 _6325_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_40_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4388__C _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5104__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6256_ _6253_/Y _8455_/B _6254_/Y _4891_/X _6255_/Y vssd1 vssd1 vccd1 vccd1 _6257_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6301__A1 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6301__B2 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5207_ input90/X _5192_/X input27/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__o22a_1
X_6187_ _6908_/A _7316_/A _8924_/B _7683_/A vssd1 vssd1 vccd1 vccd1 _6188_/B sky130_fd_sc_hd__a22o_1
XANTENNA__7061__A _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8054__A1 _8054_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5138_ _5031_/X _7352_/B _5135_/Y _5137_/X vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__a22o_2
XANTENNA__8054__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7801__A1 _7798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6604__A2 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7801__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5069_ _5715_/B vssd1 vssd1 vccd1 vccd1 _6233_/B sky130_fd_sc_hd__buf_6
XFILLER_0_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8357__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8000__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6368__A1 _6368_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6405__A _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8828_ _8222_/X _8782_/A _8827_/X vssd1 vssd1 vccd1 vccd1 _8828_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_149_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7000__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6368__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7565__B1 _6771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4918__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8759_ _8759_/A _8759_/B vssd1 vssd1 vccd1 vccd1 _8759_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__5040__A1 _5131_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8109__A2 _8499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5040__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8514__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7868__A1 _7877_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7868__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7236__A _7236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8293__A1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7096__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8293__B2 _7796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6056__B1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6359__A1 _6358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6315__A hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5582__A2 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4440_ _8584_/B _4748_/B vssd1 vssd1 vccd1 vccd1 _7510_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4371_ _4675_/A _4674_/A _4674_/B vssd1 vssd1 vccd1 vccd1 _4668_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6110_ _6110_/A _6689_/S vssd1 vssd1 vccd1 vccd1 _6110_/Y sky130_fd_sc_hd__nand2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _5094_/A _7059_/X _5336_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7090_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6013_/Y _6040_/Y _8188_/S vssd1 vssd1 vccd1 vccd1 _6041_/X sky130_fd_sc_hd__mux2_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6834__A2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6209__B _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7992_ _7989_/Y _5117_/A _7990_/Y _7013_/A _7991_/Y vssd1 vssd1 vccd1 vccd1 _8400_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7795__B1 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6943_ _6941_/B _6908_/B _6939_/X _6940_/Y _6942_/X vssd1 vssd1 vccd1 vccd1 _6943_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8424__B _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6874_ _6866_/X _6871_/Y _6872_/X _6873_/X vssd1 vssd1 vccd1 vccd1 _6874_/X sky130_fd_sc_hd__a31o_2
XFILLER_0_92_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8613_ _7888_/Y _8581_/A _7890_/Y _8583_/A vssd1 vssd1 vccd1 vccd1 _8613_/X sky130_fd_sc_hd__a22o_1
X_5825_ _5825_/A1 _4871_/A input51/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8544_ _8349_/A _8806_/A _8539_/Y _8543_/X vssd1 vssd1 vccd1 vccd1 _8544_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5756_ _5787_/A1 _5090_/A input50/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_106_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5573__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4707_ _4707_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__nand2_1
X_8475_ _8475_/A vssd1 vssd1 vccd1 vccd1 _8475_/X sky130_fd_sc_hd__buf_1
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5687_ _5274_/A _5718_/A1 _5275_/A input47/X vssd1 vssd1 vccd1 vccd1 _5687_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7426_ _7378_/X _5362_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7428_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__5325__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4638_ hold31/A vssd1 vssd1 vccd1 vccd1 _8875_/B sky130_fd_sc_hd__clkinv_8
XFILLER_0_115_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4399__B _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4533__B1 _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7357_ _7355_/X _7332_/A _7356_/Y vssd1 vssd1 vccd1 vccd1 _7357_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4569_ _4481_/B _7311_/A _4567_/Y _4568_/X vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6308_ _6312_/A _7725_/B _7398_/A vssd1 vssd1 vccd1 vccd1 _6312_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__8275__A1 _7786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8275__B2 _8232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7288_ _6994_/C _7288_/B vssd1 vssd1 vccd1 vccd1 _7288_/X sky130_fd_sc_hd__and2b_1
XANTENNA__6286__B1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6239_ _6248_/A1 _8335_/B input5/X _4913_/A _6238_/X vssd1 vssd1 vccd1 vccd1 _7707_/D
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6825__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__A1 hold10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8027__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7786__B1 _7791_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5958__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8334__B _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7538__B1 _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8735__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8750__A2 _8366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5564__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8496__S _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5913__S _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7413__B _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8018__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput250 sports_i[118] vssd1 vssd1 vccd1 vccd1 _8011_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput261 sports_i[128] vssd1 vssd1 vccd1 vccd1 _8151_/A sky130_fd_sc_hd__clkbuf_4
Xinput272 sports_i[15] vssd1 vssd1 vccd1 vccd1 _7990_/A sky130_fd_sc_hd__buf_1
XANTENNA__8569__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output411_A _8044_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput283 sports_i[25] vssd1 vssd1 vccd1 vccd1 _8123_/A sky130_fd_sc_hd__buf_1
XANTENNA__8525__A _8555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput294 sports_i[35] vssd1 vssd1 vccd1 vccd1 _7791_/A1 sky130_fd_sc_hd__buf_2
XANTENNA_output509_A _6970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7241__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7793__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6201__B1 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5610_ _5610_/A _6081_/S vssd1 vssd1 vccd1 vccd1 _5611_/A sky130_fd_sc_hd__nand2_1
X_6590_ _6780_/A _6590_/B vssd1 vssd1 vccd1 vccd1 _6590_/X sky130_fd_sc_hd__or2_1
XANTENNA__5555__A2 _5500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6699__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5541_ _5539_/X _7629_/B _6837_/A _5540_/Y vssd1 vssd1 vccd1 vccd1 _5541_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_54_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8260_ _7765_/X _8304_/A _7771_/X _8299_/A vssd1 vssd1 vccd1 vccd1 _8260_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5472_ _5637_/A1 _8709_/B input44/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5307__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7211_ _6107_/A _7138_/X _7209_/X _7210_/X vssd1 vssd1 vccd1 vccd1 _7211_/X sky130_fd_sc_hd__o22a_2
Xoutput702 _6664_/X vssd1 vssd1 vccd1 vccd1 sports_o[75] sky130_fd_sc_hd__buf_12
XFILLER_0_112_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput713 _6754_/X vssd1 vssd1 vccd1 vccd1 sports_o[85] sky130_fd_sc_hd__buf_12
X_4423_ _8239_/A _4423_/B vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8191_ _8187_/X _7768_/X _8190_/X _7772_/X _7774_/X vssd1 vssd1 vccd1 vccd1 _8191_/Y
+ sky130_fd_sc_hd__a221oi_1
Xoutput724 _6887_/X vssd1 vssd1 vccd1 vccd1 sports_o[95] sky130_fd_sc_hd__buf_12
XFILLER_0_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7604__A _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7142_ _7141_/X _5679_/A _7175_/S vssd1 vssd1 vccd1 vccd1 _7143_/A sky130_fd_sc_hd__mux2_1
X_4354_ hold39/A vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__inv_2
XANTENNA__4947__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7073_ _7072_/X _6567_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7074_/A sky130_fd_sc_hd__mux2_1
X_6024_ _6024_/A _6074_/A vssd1 vssd1 vccd1 vccd1 _6051_/A sky130_fd_sc_hd__nor2_1
XANTENNA__8009__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7480__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5491__A1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5491__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5778__B _5893_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7232__A2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7975_ _7975_/A vssd1 vssd1 vccd1 vccd1 _7975_/X sky130_fd_sc_hd__buf_6
XANTENNA__5243__A1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5243__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6926_ _6926_/A _6926_/B vssd1 vssd1 vccd1 vccd1 _6926_/X sky130_fd_sc_hd__or2_1
XANTENNA__5794__A2 _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6857_ _6847_/A _7536_/B _7707_/B _6868_/A vssd1 vssd1 vccd1 vccd1 _6858_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7485__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5808_ _6079_/A _5865_/A vssd1 vssd1 vccd1 vccd1 _5904_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_119_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5546__A2 _5530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6788_ _6801_/A _6788_/B vssd1 vssd1 vccd1 vccd1 _6788_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8527_ _8567_/B _8133_/Y _8497_/S vssd1 vssd1 vccd1 vccd1 _8527_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5739_ _5731_/X _5737_/Y _5738_/X _6170_/A vssd1 vssd1 vccd1 vccd1 _5739_/X sky130_fd_sc_hd__a31o_2
XANTENNA__6402__B _7756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8496__A1 _8516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8458_ _8458_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7409_ _7590_/A _7409_/B vssd1 vssd1 vccd1 vccd1 _7409_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6829__S _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8389_ _8349_/A _8379_/X _8382_/Y _8388_/X vssd1 vssd1 vccd1 vccd1 _8389_/X sky130_fd_sc_hd__o22a_2
XFILLER_0_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8248__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8248__B2 _8252_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6259__B1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8799__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7471__A2 _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5969__A _5993_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4873__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8345__A _8345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8420__A1 _8009_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7223__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8420__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5234__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6982__A1 _4793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5785__A2 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8184__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6734__A1 _6743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7931__B1 _7931_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6734__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7408__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8487__A1 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8487__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6498__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output459_A _8534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5643__S _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5170__B1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7998__B1 _7998_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7462__A2 _5460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5473__A1 _5596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5879__A _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5473__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6670__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8411__A1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7214__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__A1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7760_ _7975_/A vssd1 vssd1 vccd1 vccd1 _7760_/X sky130_fd_sc_hd__clkbuf_8
X_4972_ _8166_/A vssd1 vssd1 vccd1 vccd1 _6017_/A sky130_fd_sc_hd__buf_8
XFILLER_0_148_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6973__A1 _6326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6711_ _5670_/B _5580_/X _6711_/S vssd1 vssd1 vccd1 vccd1 _6711_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7691_ _7692_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6642_ _6642_/A vssd1 vssd1 vccd1 vccd1 _6642_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5528__A2 _5496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6573_ _6593_/A _6573_/B vssd1 vssd1 vccd1 vccd1 _6573_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8312_ _7788_/X hold36/A _8482_/B vssd1 vssd1 vccd1 vccd1 _8312_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_42_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5524_ _7829_/A _5517_/Y _5727_/A vssd1 vssd1 vccd1 vccd1 _5524_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8243_ _7761_/A _8251_/A2 _6059_/B _8252_/A1 vssd1 vssd1 vccd1 vccd1 _8243_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5455_ _6084_/B _6648_/B _5447_/X _5715_/B _5454_/Y vssd1 vssd1 vccd1 vccd1 _5455_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput510 _6975_/X vssd1 vssd1 vccd1 vccd1 sports_o[107] sky130_fd_sc_hd__buf_12
XANTENNA__7150__A1 _6732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput521 _7338_/X vssd1 vssd1 vccd1 vccd1 sports_o[117] sky130_fd_sc_hd__buf_12
XANTENNA__6876__C _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7334__A _7334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput532 _7429_/X vssd1 vssd1 vccd1 vccd1 sports_o[127] sky130_fd_sc_hd__buf_12
X_4406_ _4406_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__nor2_1
Xoutput543 _7508_/X vssd1 vssd1 vccd1 vccd1 sports_o[137] sky130_fd_sc_hd__buf_12
XANTENNA__5161__B1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8174_ _8174_/A _8174_/B vssd1 vssd1 vccd1 vccd1 _8174_/Y sky130_fd_sc_hd__nand2_1
Xoutput554 _7600_/X vssd1 vssd1 vccd1 vccd1 sports_o[147] sky130_fd_sc_hd__buf_12
X_5386_ _5386_/A vssd1 vssd1 vccd1 vccd1 _5386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5700__A2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput565 _7693_/X vssd1 vssd1 vccd1 vccd1 sports_o[157] sky130_fd_sc_hd__buf_12
Xoutput576 _7742_/X vssd1 vssd1 vccd1 vccd1 sports_o[167] sky130_fd_sc_hd__buf_12
Xoutput587 _5138_/X vssd1 vssd1 vccd1 vccd1 sports_o[177] sky130_fd_sc_hd__buf_12
X_7125_ _7125_/A vssd1 vssd1 vccd1 vccd1 _7125_/X sky130_fd_sc_hd__buf_1
Xoutput598 _5433_/X vssd1 vssd1 vccd1 vccd1 sports_o[187] sky130_fd_sc_hd__buf_12
X_4337_ _4337_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4338_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7056_ _5105_/A _7026_/X _7054_/Y _7055_/X vssd1 vssd1 vccd1 vccd1 _7056_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5464__A1 _5440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6007_ _6007_/A1 _8271_/B input57/X _4917_/A vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5464__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7205__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8402__B2 _8376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5216__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _7958_/A1 _7876_/X _7958_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7958_/Y sky130_fd_sc_hd__o22ai_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6909_/A vssd1 vssd1 vccd1 vccd1 _7668_/A sky130_fd_sc_hd__inv_2
X_7889_ _5185_/A _7882_/Y _7881_/Y _5682_/B vssd1 vssd1 vccd1 vccd1 _7889_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8705__A2 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6716__A1 _5679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7913__B1 _7918_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6716__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4868__A _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7141__A1 _5628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5152__B1 _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8641__A1 _7999_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__A1 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__B2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5207__A1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5207__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__A2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6955__A1 _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8157__B1 _8162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__C1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6707__A1 _5552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7904__B1 _7903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6707__B2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7132__A1 _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5240_ _8194_/A vssd1 vssd1 vccd1 vccd1 _8924_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__5694__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5694__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5171_ _6024_/A _5171_/B vssd1 vssd1 vccd1 vccd1 _6166_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8632__A1 _8369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8930_ _8934_/A _8934_/B _8930_/C vssd1 vssd1 vccd1 vccd1 _8931_/B sky130_fd_sc_hd__nand3_1
Xinput3 mports_i[101] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5402__A _5402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8861_ _8861_/A _8865_/B vssd1 vssd1 vccd1 vccd1 _8861_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7199__A1 _5923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8396__B1 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7812_ _7809_/X _7768_/X _7811_/X _7772_/X _7774_/X vssd1 vssd1 vccd1 vccd1 _7812_/X
+ sky130_fd_sc_hd__a221o_1
X_8792_ _8491_/A _8806_/B _8790_/X _8791_/X vssd1 vssd1 vccd1 vccd1 _8792_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6946__A1 _6207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7743_ _7743_/A _7753_/B vssd1 vssd1 vccd1 vccd1 _7743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4955_ _4956_/A _4953_/X _4957_/A _4870_/A _4954_/X vssd1 vssd1 vccd1 vccd1 _6440_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8148__B1 _8142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7329__A _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7674_ _7378_/X _6908_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7674_/X sky130_fd_sc_hd__o21a_1
X_4886_ _4886_/A vssd1 vssd1 vccd1 vccd1 _8455_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_129_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8699__B2 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6625_ _6620_/Y _6450_/X _6621_/Y _6623_/Y _6624_/X vssd1 vssd1 vccd1 vccd1 _6625_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6174__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7371__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6556_ _5212_/B _6426_/A _6585_/A _6511_/A _6555_/X vssd1 vssd1 vccd1 vccd1 _6556_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__5921__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5507_ _4893_/A _5557_/A1 _4896_/A input40/X vssd1 vssd1 vccd1 vccd1 _5507_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6487_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6487_/X sky130_fd_sc_hd__buf_1
XANTENNA__7123__A1 _5544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8320__B1 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8226_ _8235_/A1 _6059_/B _8235_/B1 _5359_/B _8225_/X vssd1 vssd1 vccd1 vccd1 _8226_/X
+ sky130_fd_sc_hd__a221o_4
X_5438_ _5435_/Y _4890_/A _5436_/Y _4886_/A _5437_/Y vssd1 vssd1 vccd1 vccd1 _6669_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7674__A2 _6908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput373 _8737_/X vssd1 vssd1 vccd1 vccd1 mports_o[106] sky130_fd_sc_hd__buf_12
XANTENNA__8594__S _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8157_ _8175_/A1 _6626_/B _8162_/A _6941_/A _8156_/X vssd1 vssd1 vccd1 vccd1 _8157_/X
+ sky130_fd_sc_hd__o221a_4
X_5369_ _5294_/A _5111_/A _5295_/A _4932_/A _5368_/X vssd1 vssd1 vccd1 vccd1 _6611_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_11_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput384 _8773_/X vssd1 vssd1 vccd1 vccd1 mports_o[116] sky130_fd_sc_hd__buf_12
Xoutput395 _8807_/Y vssd1 vssd1 vccd1 vccd1 mports_o[126] sky130_fd_sc_hd__buf_12
X_7108_ _7107_/X _5460_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7109_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7426__A2 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8088_ _8093_/A1 _5146_/A _8093_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _8088_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__5437__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7039_ _5064_/B _7138_/A _7038_/X vssd1 vssd1 vccd1 vccd1 _7040_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8387__B1 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4660__A2 _5359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6398__C1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5458__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8614__A1 _8334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7417__A2 _5328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5428__A1 _6634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8090__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4740_ hold32/A _4953_/A vssd1 vssd1 vccd1 vccd1 _4740_/Y sky130_fd_sc_hd__nor2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4671_ _4674_/B _8512_/S vssd1 vssd1 vccd1 vccd1 _4672_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6410_ _6475_/A vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7390_ _6551_/Y _7696_/B _7379_/Y _7700_/B vssd1 vssd1 vccd1 vccd1 _7390_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5903__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6341_ _6224_/S _7733_/B _6338_/X _6340_/Y vssd1 vssd1 vccd1 vccd1 _6341_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6272_ input70/X _8579_/C _6286_/A1 _8713_/C _6271_/X vssd1 vssd1 vccd1 vccd1 _6272_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8011_ _8011_/A1 _7876_/X _8011_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _8011_/Y sky130_fd_sc_hd__o22ai_2
X_5223_ input92/X _5192_/X input29/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_110_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8708__A _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8066__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8605__A1 _7821_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5154_ _5031_/X _7356_/B _5153_/X vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5419__A1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8427__B _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5419__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5085_ input85/X _8310_/B input22/X _4874_/X vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8081__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4674__C _4674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8913_ _8913_/A hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8844_ _8844_/A _8846_/B vssd1 vssd1 vccd1 vccd1 _8861_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5987_ _5159_/B _5924_/A _5125_/X _7619_/A _5986_/X vssd1 vssd1 vccd1 vccd1 _5987_/X
+ sky130_fd_sc_hd__a221o_1
X_8775_ _8833_/B _7999_/Y _8725_/A vssd1 vssd1 vccd1 vccd1 _8775_/X sky130_fd_sc_hd__o21a_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7059__A _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4938_ _4938_/A vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__clkbuf_8
X_7726_ _7724_/Y _7332_/A _7725_/Y vssd1 vssd1 vccd1 vccd1 _7726_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6147__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4869_ _5089_/A vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__buf_8
XFILLER_0_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7344__A1 _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7657_ _7701_/A _7657_/B vssd1 vssd1 vccd1 vccd1 _7657_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__8541__B1 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6608_ _6606_/X _6933_/A _6968_/A _6607_/X vssd1 vssd1 vccd1 vccd1 _6608_/X sky130_fd_sc_hd__a211o_1
XANTENNA__7895__A2 _7886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7588_ _7378_/X _5853_/X _7683_/C vssd1 vssd1 vccd1 vccd1 _7590_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6539_ _7383_/A _8140_/A _5161_/X _5299_/B vssd1 vssd1 vccd1 vccd1 _6539_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5107__B1 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7647__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8209_ _8181_/A _8209_/A2 _8208_/X vssd1 vssd1 vccd1 vccd1 _8209_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6083__A1 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5042__A _5106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6083__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4881__A _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5188__S _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7583__B2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6138__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7335__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8532__B1 _8169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7886__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5897__A1 _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6320__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8835__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5649__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5649__B2 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output441_A _8357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6310__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7432__A _7532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8063__A2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output706_A _6703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5821__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5910_ _5962_/A1 _8709_/B input55/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5910_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_49_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6890_ _7637_/B _6912_/B vssd1 vssd1 vccd1 vccd1 _6890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8220__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5841_ _5841_/A vssd1 vssd1 vccd1 vccd1 _5842_/A sky130_fd_sc_hd__inv_2
XANTENNA__6377__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8771__B1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7574__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5772_ _5788_/A1 _5111_/A _5788_/B1 _4931_/A _5771_/X vssd1 vssd1 vccd1 vccd1 _5772_/X
+ sky130_fd_sc_hd__o221a_4
X_8560_ _8567_/B _8222_/X _8497_/S vssd1 vssd1 vccd1 vccd1 _8560_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7511_ _7511_/A _7511_/B vssd1 vssd1 vccd1 vccd1 _7512_/A sky130_fd_sc_hd__nand2_2
X_4723_ _4762_/A _4800_/B _4762_/B vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__nand3_1
X_8491_ _8491_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8491_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7607__A _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7442_ _6637_/A _7361_/X _7440_/X _7754_/A _7441_/Y vssd1 vssd1 vccd1 vccd1 _7442_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7877__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ hold44/A vssd1 vssd1 vccd1 vccd1 _8845_/C sky130_fd_sc_hd__clkinv_4
XANTENNA__6511__A _6511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5888__A1 _5885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput50 mports_i[144] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5888__B2 _5899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput61 mports_i[154] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7373_ _7700_/B vssd1 vssd1 vccd1 vccd1 _7691_/B sky130_fd_sc_hd__buf_4
XFILLER_0_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput72 mports_i[164] vssd1 vssd1 vccd1 vccd1 _6314_/B sky130_fd_sc_hd__buf_2
X_4585_ _4810_/B _5193_/A _4800_/B _5192_/A _4584_/Y vssd1 vssd1 vccd1 vccd1 _4793_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput83 mports_i[174] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_4
Xinput94 mports_i[184] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_2
X_6324_ _5845_/B _6971_/A _5128_/A _6317_/X _6323_/X vssd1 vssd1 vccd1 vccd1 _6324_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6255_ _4893_/A _6262_/A1 _8579_/C input69/X vssd1 vssd1 vccd1 vccd1 _6255_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__8438__A _8438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6301__A2 _6309_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5206_ _6550_/A _6234_/B _7383_/A _5128_/A vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6186_ _6184_/Y _6185_/Y _8842_/B vssd1 vssd1 vccd1 vccd1 _6186_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4685__B _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5137_ _6202_/B _6507_/B _5136_/X vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__o21a_1
XANTENNA__8054__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6065__A1 _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7801__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5068_ _5031_/X _7341_/B _5067_/X vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5812__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7014__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8827_ _8217_/X _8738_/A _8219_/X _8711_/A _8824_/S vssd1 vssd1 vccd1 vccd1 _8827_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6368__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7565__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8758_ _4930_/X _8345_/A _8829_/S _8757_/X vssd1 vssd1 vccd1 vccd1 _8758_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5040__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7709_ _7707_/D _7681_/A _7707_/X _7708_/X vssd1 vssd1 vccd1 vccd1 _7709_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_118_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8689_ _8688_/X _8211_/A _8689_/S vssd1 vssd1 vccd1 vccd1 _8689_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7868__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8293__A2 _7821_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5500__B1 _5506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6056__A1 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6315__B _6315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8753__B1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8811__A _8811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7308__A1 _4876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7308__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5582__A3 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6531__A2 _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4370_ _4715_/B _4800_/B vssd1 vssd1 vccd1 vccd1 _4674_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8258__A _8429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__B2 _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6040_ _7660_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6040_/Y sky130_fd_sc_hd__nand2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7795__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7991_ _7998_/A1 _4946_/A _7998_/B1 _5119_/A vssd1 vssd1 vccd1 vccd1 _7991_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7795__B2 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6942_ _8857_/B _6939_/X _8574_/B _6941_/X vssd1 vssd1 vccd1 vccd1 _6942_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6873_ _6059_/A _6908_/B _7619_/A _6512_/X vssd1 vssd1 vccd1 vccd1 _6873_/X sky130_fd_sc_hd__a22o_1
X_8612_ _7867_/Y _8577_/X _8610_/X _8611_/X vssd1 vssd1 vccd1 vccd1 _8612_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5824_ _5809_/A _5111_/A _5810_/A _4931_/A _5823_/X vssd1 vssd1 vccd1 vccd1 _5824_/X
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5558__B1 _5506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8543_ _8543_/A _8564_/B vssd1 vssd1 vccd1 vccd1 _8543_/X sky130_fd_sc_hd__and2_1
XFILLER_0_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5755_ _5999_/B _5745_/Y _5754_/Y _5174_/A vssd1 vssd1 vccd1 vccd1 _5755_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4706_ _4706_/A _4706_/B vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__nand2_1
X_5686_ _5686_/A vssd1 vssd1 vccd1 vccd1 _5686_/Y sky130_fd_sc_hd__inv_2
X_8474_ _8473_/X _8491_/A _8572_/S vssd1 vssd1 vccd1 vccd1 _8475_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4637_ _4637_/A vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__clkinv_4
X_7425_ _5356_/B _7696_/B _7423_/X _7326_/A _7424_/X vssd1 vssd1 vccd1 vccd1 _7425_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4533__A1 _4557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4568_ _5229_/A _4478_/B _4597_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__a22o_1
X_7356_ _7756_/A _7356_/B vssd1 vssd1 vccd1 vccd1 _7356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6307_ _6305_/X _6233_/B _6386_/S _6306_/X vssd1 vssd1 vccd1 vccd1 _6307_/X sky130_fd_sc_hd__a211o_1
X_7287_ _6379_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7287_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8275__A2 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4499_ _4499_/A _4499_/B vssd1 vssd1 vccd1 vccd1 _4613_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6286__A1 _6286_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6238_ _6247_/A1 _8271_/B input68/X _4917_/A vssd1 vssd1 vccd1 vccd1 _6238_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6286__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4836__A2 _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8027__A2 _8433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6284_/A _6115_/A _5762_/A _6156_/Y _6168_/Y vssd1 vssd1 vccd1 vccd1 _6170_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6038__A1 _6104_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6038__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7786__A1 _7791_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6589__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7786__B2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7538__A1 _7535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8735__B1 _7832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6210__A1 _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8964__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7710__A1 _6248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5721__B1 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8671__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8018__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput240 sports_i[109] vssd1 vssd1 vccd1 vccd1 _7882_/A sky130_fd_sc_hd__clkbuf_2
Xinput251 sports_i[119] vssd1 vssd1 vccd1 vccd1 _8024_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7226__A0 _7225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput262 sports_i[129] vssd1 vssd1 vccd1 vccd1 _8172_/B sky130_fd_sc_hd__clkbuf_4
Xinput273 sports_i[16] vssd1 vssd1 vccd1 vccd1 _8002_/A sky130_fd_sc_hd__buf_1
Xinput284 sports_i[26] vssd1 vssd1 vccd1 vccd1 _8148_/A1 sky130_fd_sc_hd__buf_2
Xinput295 sports_i[36] vssd1 vssd1 vccd1 vccd1 _4326_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5788__B1 _5788_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output404_A _8837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6985__C1 _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5230__A _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6201__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6752__A2 _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5540_ _6304_/A _7120_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _5540_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5471_ _5466_/Y _5470_/Y _6793_/S vssd1 vssd1 vccd1 vccd1 _7474_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7162__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7210_ _6891_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7210_/X sky130_fd_sc_hd__a21o_1
Xoutput703 _6675_/X vssd1 vssd1 vccd1 vccd1 sports_o[76] sky130_fd_sc_hd__buf_12
X_4422_ _5145_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4423_/B sky130_fd_sc_hd__nor2_1
X_8190_ _8196_/B1 _6500_/X _8188_/X hold23/A _8189_/X vssd1 vssd1 vccd1 vccd1 _8190_/X
+ sky130_fd_sc_hd__a221o_4
Xoutput714 _6769_/X vssd1 vssd1 vccd1 vccd1 sports_o[86] sky130_fd_sc_hd__buf_12
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput725 _6896_/X vssd1 vssd1 vccd1 vccd1 sports_o[96] sky130_fd_sc_hd__buf_12
XFILLER_0_50_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7141_ _5628_/A _7138_/X _7139_/X _7140_/X vssd1 vssd1 vccd1 vccd1 _7141_/X sky130_fd_sc_hd__o22a_2
XANTENNA_hold41_A hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4353_ _4350_/Y _4351_/Y _4674_/C vssd1 vssd1 vccd1 vccd1 _4684_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5405__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6268__B2 _6263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7465__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7072_ _6566_/B _7026_/X _7070_/X _7071_/X vssd1 vssd1 vccd1 vccd1 _7072_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6023_ _6020_/Y _4885_/A _6021_/Y _4890_/A _6022_/Y vssd1 vssd1 vccd1 vccd1 _6074_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__8009__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8716__A _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5491__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5779__B1 _5766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7974_ _7760_/X _8375_/A _7970_/X _7973_/X vssd1 vssd1 vccd1 vccd1 _7974_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5243__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8950__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6925_ _7681_/B _6925_/B vssd1 vssd1 vccd1 vccd1 _6925_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8451__A _8451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6856_ _6856_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_147_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5807_ _5804_/Y _4886_/A _5805_/Y _4891_/A _5806_/Y vssd1 vssd1 vccd1 vccd1 _5865_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6787_ _7570_/B _6871_/B vssd1 vssd1 vccd1 vccd1 _6787_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7940__B2 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8526_ _8550_/A _8304_/X _8130_/Y _8299_/X _8496_/S vssd1 vssd1 vccd1 vccd1 _8526_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5738_ _6312_/A _7297_/B _5738_/C vssd1 vssd1 vccd1 vccd1 _5738_/X sky130_fd_sc_hd__or3_1
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8457_ _8457_/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5669_ _5606_/A _5609_/Y _7829_/A vssd1 vssd1 vccd1 vccd1 _5670_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7408_ _7409_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7408_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8388_ _8388_/A _8564_/B vssd1 vssd1 vccd1 vccd1 _8388_/X sky130_fd_sc_hd__and2_1
XFILLER_0_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7514__B _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7339_ _5050_/Y _7349_/A _7037_/Y _7753_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7339_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6259__A1 _6262_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6259__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7535__A1_N _6727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8345__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8420__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A2 _6567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6982__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8184__A1 _8820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7931__A1 _7931_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6734__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7931__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7144__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6498__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7705__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7695__B1 _6221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5170__A1 _7383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8644__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7998__A1 _7998_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7998__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5473__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6670__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5879__B _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5225__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4971_ _6461_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _5022_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6973__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6710_ _5644_/A _6908_/B _5647_/B _6512_/X _6709_/X vssd1 vssd1 vccd1 vccd1 _6710_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6490__S _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8271__A _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8175__A1 _8175_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7690_ _7378_/X _6185_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7692_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6641_ _7459_/A _8151_/B _5197_/X _6635_/A vssd1 vssd1 vccd1 vccd1 _6642_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5933__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6572_ _6562_/Y _6450_/X _6565_/Y _6566_/X _6571_/X vssd1 vssd1 vccd1 vccd1 _6572_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8311_ _8311_/A vssd1 vssd1 vccd1 vccd1 _8482_/B sky130_fd_sc_hd__inv_2
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5523_ _5523_/A _6081_/S vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8242_ _8238_/Y _8241_/X _4662_/C _7760_/X vssd1 vssd1 vccd1 vccd1 _8242_/X sky130_fd_sc_hd__a22o_2
X_5454_ _5762_/A _5454_/B vssd1 vssd1 vccd1 vccd1 _5454_/Y sky130_fd_sc_hd__nor2_1
Xoutput500 _8699_/X vssd1 vssd1 vccd1 vccd1 mports_o[99] sky130_fd_sc_hd__buf_12
Xoutput511 _6979_/X vssd1 vssd1 vccd1 vccd1 sports_o[108] sky130_fd_sc_hd__buf_12
XANTENNA__7150__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput522 _7342_/Y vssd1 vssd1 vccd1 vccd1 sports_o[118] sky130_fd_sc_hd__buf_12
X_4405_ _4405_/A vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__inv_2
XANTENNA__5161__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput533 _7437_/X vssd1 vssd1 vccd1 vccd1 sports_o[128] sky130_fd_sc_hd__buf_12
X_5385_ _5385_/A vssd1 vssd1 vccd1 vccd1 _5385_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5161__B2 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8173_ _8173_/A hold12/A vssd1 vssd1 vccd1 vccd1 _8173_/Y sky130_fd_sc_hd__nand2_1
Xoutput544 _7521_/X vssd1 vssd1 vccd1 vccd1 sports_o[138] sky130_fd_sc_hd__buf_12
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput555 _7608_/X vssd1 vssd1 vccd1 vccd1 sports_o[148] sky130_fd_sc_hd__buf_12
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput566 _7702_/X vssd1 vssd1 vccd1 vccd1 sports_o[158] sky130_fd_sc_hd__buf_12
XFILLER_0_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput577 _7747_/Y vssd1 vssd1 vccd1 vccd1 sports_o[168] sky130_fd_sc_hd__buf_12
X_7124_ _7123_/X _5530_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7125_/A sky130_fd_sc_hd__mux2_2
X_4336_ _7847_/A _4478_/B vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__nand2_1
Xoutput588 _5154_/X vssd1 vssd1 vccd1 vccd1 sports_o[178] sky130_fd_sc_hd__buf_12
Xoutput599 _5462_/X vssd1 vssd1 vccd1 vccd1 sports_o[188] sky130_fd_sc_hd__buf_12
X_7055_ _7055_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7055_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5464__A2 _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6006_ _6006_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _6006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7957_ _8358_/A _7954_/X _7956_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7957_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8181__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6908_ _6908_/A _6908_/B vssd1 vssd1 vccd1 vccd1 _6908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7888_ _7881_/Y _5299_/B _7882_/Y _5171_/B _7887_/X vssd1 vssd1 vccd1 vccd1 _7888_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7509__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6839_ _6852_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6839_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7913__A1 _7918_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6716__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6413__B _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7913__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8509_ _8323_/X _8502_/Y _8507_/X _8508_/X vssd1 vssd1 vccd1 vccd1 _8509_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7126__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7141__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5152__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7260__A _7260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6652__A1 _5460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__A2 _6648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5207__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7601__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8803__B _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4966__A1 _4956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4966__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8157__A1 _8175_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8157__B2 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7904__A1 _7901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6707__A2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7904__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4778__B _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5170_ _7383_/A _5299_/B _6470_/B _7071_/A vssd1 vssd1 vccd1 vccd1 _6590_/B sky130_fd_sc_hd__a22o_1
XANTENNA__6485__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8093__B1 _8093_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8632__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7170__A _7170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput4 mports_i[102] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8860_ _8893_/A _8860_/B vssd1 vssd1 vccd1 vccd1 _8865_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8396__B2 _8359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7811_ _7814_/A1 _5185_/A _7814_/B1 _7299_/A _7810_/X vssd1 vssd1 vccd1 vccd1 _7811_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8791_ _8833_/B _8068_/Y _8725_/A vssd1 vssd1 vccd1 vccd1 _8791_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8713__B _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7742_ _7742_/A vssd1 vssd1 vccd1 vccd1 _7742_/X sky130_fd_sc_hd__buf_1
XANTENNA__6514__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4954_ input81/X _5090_/A input18/X _4874_/A vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8148__A1 _8148_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8148__B2 _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6159__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6233__B _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7673_ _7673_/A _7673_/B vssd1 vssd1 vccd1 vccd1 _7673_/X sky130_fd_sc_hd__or2_1
X_4885_ _4885_/A vssd1 vssd1 vccd1 vccd1 _4886_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6624_ _5367_/A _6510_/A _5374_/Y _6512_/X vssd1 vssd1 vccd1 vccd1 _6624_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_117_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7371__A2 _5159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5382__A1 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6555_ _6542_/Y _6467_/X _6548_/X _6550_/Y _6554_/X vssd1 vssd1 vccd1 vccd1 _6555_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__7345__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5506_ _5506_/A vssd1 vssd1 vccd1 vccd1 _5506_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6486_ _6485_/X _7341_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6487_/A sky130_fd_sc_hd__mux2_4
XANTENNA__8320__A1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7123__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4688__B _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8320__B2 _7807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8225_ _7761_/A _8234_/A2 _8857_/B _8234_/B2 vssd1 vssd1 vccd1 vccd1 _8225_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6331__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5437_ _5274_/A _5497_/A1 _5275_/X input38/X vssd1 vssd1 vccd1 vccd1 _5437_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5368_ input95/X _4935_/A input32/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5368_/X sky130_fd_sc_hd__o22a_1
Xoutput374 _8741_/Y vssd1 vssd1 vccd1 vccd1 mports_o[107] sky130_fd_sc_hd__buf_12
X_8156_ _8172_/B _4947_/B _8158_/A _5123_/A vssd1 vssd1 vccd1 vccd1 _8156_/X sky130_fd_sc_hd__o22a_1
Xoutput385 _8776_/X vssd1 vssd1 vccd1 vccd1 mports_o[117] sky130_fd_sc_hd__buf_12
Xoutput396 _8811_/X vssd1 vssd1 vccd1 vccd1 mports_o[127] sky130_fd_sc_hd__buf_12
XFILLER_0_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7107_ _7459_/A _7026_/X _7105_/X _7106_/X vssd1 vssd1 vccd1 vccd1 _7107_/X sky130_fd_sc_hd__o22a_2
X_4319_ _4319_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__nand2_1
X_8087_ _8084_/Y _5116_/A _8085_/Y _7013_/A _8086_/Y vssd1 vssd1 vccd1 vccd1 _8490_/A
+ sky130_fd_sc_hd__a221oi_4
X_5299_ _7083_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5299_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5437__A2 _5497_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7038_ _5050_/Y _7088_/A _7037_/Y _7059_/A _7089_/A vssd1 vssd1 vccd1 vccd1 _7038_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4645__B1 _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8387__A1 _8384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8387__B2 _8386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__A _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7898__B1 _7905_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5982__B _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5373__A1 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4879__A _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8785__S _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6873__A1 _6059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6873__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5428__A2 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output686_A _6479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7889__B1 _7881_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4670_ _4670_/A _4670_/B vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_56_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7353__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5364__A1 _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7165__A _7165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6340_ _6340_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6340_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8838__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8302__A1 _7765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6271_ _8444_/A _6287_/A1 _8257_/C input7/X vssd1 vssd1 vccd1 vccd1 _6271_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8853__A2 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5222_ input12/X _8271_/A _5222_/B1 _5191_/X _5221_/X vssd1 vssd1 vccd1 vccd1 _6566_/B
+ sky130_fd_sc_hd__o221a_4
X_8010_ _8416_/A _7954_/X _8009_/Y _7826_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _8010_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6864__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4875__B1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8066__B1 _8469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5153_ _5148_/Y _6128_/B _5151_/Y _5152_/Y vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__a31o_1
XANTENNA__8605__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5419__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7813__B1 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5084_ _5139_/A _5080_/A _5140_/A _4870_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5150_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8912_ _8912_/A vssd1 vssd1 vccd1 vccd1 _8950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8843_ _8842_/Y _8845_/B _8846_/A vssd1 vssd1 vccd1 vccd1 _8844_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4971__B _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7041__A1 _7341_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8774_ _8424_/A _8711_/X _8407_/A _8803_/B _8820_/B vssd1 vssd1 vccd1 vccd1 _8774_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _6128_/B _6847_/A _5136_/A _5985_/X vssd1 vssd1 vccd1 vccd1 _5986_/X sky130_fd_sc_hd__o211a_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7725_ _7756_/A _7725_/B vssd1 vssd1 vccd1 vccd1 _7725_/Y sky130_fd_sc_hd__nor2_1
X_4937_ _4937_/A vssd1 vssd1 vccd1 vccd1 _4938_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7656_ _7657_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7656_/Y sky130_fd_sc_hd__nand2_1
X_4868_ _4868_/A vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__buf_8
XFILLER_0_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8541__A1 _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7344__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8541__B2 _8187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6607_ _5094_/A _6913_/B _5310_/Y _6912_/B vssd1 vssd1 vccd1 vccd1 _6607_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_117_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6552__B1 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7587_ _7583_/X _7584_/Y _7585_/X _7586_/X vssd1 vssd1 vccd1 vccd1 _7587_/X sky130_fd_sc_hd__a31o_2
XFILLER_0_144_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4799_ _4799_/A _4799_/B vssd1 vssd1 vccd1 vccd1 _4800_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6538_ _6538_/A vssd1 vssd1 vccd1 vccd1 _6585_/A sky130_fd_sc_hd__inv_2
XFILLER_0_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5107__A1 _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5107__B2 _6507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6469_ _6837_/A _6469_/B vssd1 vssd1 vccd1 vccd1 _6469_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8208_ _8150_/A _8198_/B _7707_/C vssd1 vssd1 vccd1 vccd1 _8208_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8139_ _8140_/A _8146_/B vssd1 vssd1 vccd1 vccd1 _8139_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6419__A _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5323__A _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6607__A1 _5094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7804__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6607__B2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7280__A1 _6358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4881__B _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5043__B1 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8780__A1 _8412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7583__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5594__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5993__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7335__A2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8532__A1 _8165_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8532__B2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8296__B1 _7837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8835__A2 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5649__A2 _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7432__B _7432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5821__A2 _6770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8220__B1 _8219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5827_/A _6017_/A _7299_/A _5803_/A vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_76_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5034__B1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8771__A1 _7983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7574__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5585__A1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5771_ _5787_/A1 _4934_/A input50/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5585__B2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7510_ _7510_/A _7510_/B vssd1 vssd1 vccd1 vccd1 _7511_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4722_ _4722_/A hold34/A vssd1 vssd1 vccd1 vccd1 _4762_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8490_ _8490_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7441_ _7681_/A _7441_/B vssd1 vssd1 vccd1 vccd1 _7441_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_154_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4653_ _8958_/Q vssd1 vssd1 vccd1 vccd1 _8194_/A sky130_fd_sc_hd__buf_8
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7731__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput40 mports_i[135] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__8975__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5888__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 mports_i[145] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7372_ _7372_/A _7372_/B vssd1 vssd1 vccd1 vccd1 _7700_/B sky130_fd_sc_hd__nand2_8
Xinput62 mports_i[155] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4584_ _4578_/Y _8261_/A _4583_/Y vssd1 vssd1 vccd1 vccd1 _4584_/Y sky130_fd_sc_hd__a21oi_1
Xinput73 mports_i[165] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput84 mports_i[175] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__buf_2
Xinput95 mports_i[185] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__buf_2
X_6323_ _4518_/A _6342_/A _6321_/Y _5096_/A _6322_/X vssd1 vssd1 vccd1 vccd1 _6323_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6298__C1 _7725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7623__A _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6254_ input6/X vssd1 vssd1 vccd1 vccd1 _6254_/Y sky130_fd_sc_hd__inv_2
X_5205_ _5208_/A1 _4927_/A _5208_/B1 _4931_/A _5204_/X vssd1 vssd1 vccd1 vccd1 _5211_/A
+ sky130_fd_sc_hd__o221a_4
X_6185_ _6185_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _6185_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5143__A _6514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5136_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__7262__A1 _6326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6065__A2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4982__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5067_ _5108_/A _6505_/B _6170_/A _5063_/X _5066_/X vssd1 vssd1 vccd1 vccd1 _5067_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5812__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8173__B hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7014__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7014__B2 _4408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8826_ _8826_/A vssd1 vssd1 vccd1 vccd1 _8826_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8762__A1 _7945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8757_ _7932_/Y _8833_/B _8725_/A _8756_/X vssd1 vssd1 vccd1 vccd1 _8757_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_109_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5969_ _5993_/C vssd1 vssd1 vccd1 vccd1 _7630_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6773__B1 _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7970__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7708_ _6241_/X _7347_/A _7242_/A _7349_/A _7715_/S vssd1 vssd1 vccd1 vccd1 _7708_/X
+ sky130_fd_sc_hd__a221o_1
X_8688_ _8203_/X _8580_/A _8206_/X _8583_/A vssd1 vssd1 vccd1 vccd1 _8688_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8514__A1 _8117_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8514__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7639_ _7639_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7640_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5318__A _5356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5536__A2_N _5535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5500__A1 _5505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5500__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6149__A _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5053__A _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7789__C1 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5988__A _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6056__A2 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4892__A _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8364__A _8364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5016__B1 _5004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8753__A1 _8381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5567__A1 _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7308__A2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7427__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6819__A1 _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6295__A2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7492__A1 _5548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__A _6059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5898__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7244__A1 _6248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7990_ _7990_/A vssd1 vssd1 vccd1 vccd1 _7990_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7795__A2 _7802_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6941_ _6941_/A _6941_/B vssd1 vssd1 vccd1 vccd1 _6941_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6872_ _6801_/A _6867_/A _6450_/A vssd1 vssd1 vccd1 vccd1 _6872_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8744__A1 _7867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8611_ _8698_/B _7878_/Y _8590_/X vssd1 vssd1 vccd1 vccd1 _8611_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5823_ _5825_/A1 _4934_/A input51/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5823_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5558__A1 _5505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5558__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8542_ _8190_/X _8299_/A _8803_/A _8304_/A vssd1 vssd1 vccd1 vccd1 _8543_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5754_ _5754_/A vssd1 vssd1 vccd1 vccd1 _5754_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6522__A _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4705_ _4714_/A _4705_/B vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__nand2_1
X_8473_ _8068_/Y _8567_/B _8467_/X _8472_/X vssd1 vssd1 vccd1 vccd1 _8473_/X sky130_fd_sc_hd__o22a_1
X_5685_ _5685_/A vssd1 vssd1 vccd1 vccd1 _5685_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7424_ _7424_/A _7476_/B vssd1 vssd1 vccd1 vccd1 _7424_/X sky130_fd_sc_hd__and2_1
XFILLER_0_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4636_ hold31/A hold30/A vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4977__A _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4533__A2 _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7355_ _7354_/X _5106_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7355_/X sky130_fd_sc_hd__mux2_1
XANTENNA__8449__A _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4567_ _4567_/A _7876_/A vssd1 vssd1 vccd1 vccd1 _4567_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6306_ _5845_/B _6277_/A _6278_/Y _5096_/A vssd1 vssd1 vccd1 vccd1 _6306_/X sky130_fd_sc_hd__a22o_1
X_7286_ _7286_/A vssd1 vssd1 vccd1 vccd1 _7286_/X sky130_fd_sc_hd__buf_1
X_4498_ _4498_/A _4509_/A vssd1 vssd1 vccd1 vccd1 _4499_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6286__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6237_ _6402_/A _6948_/A _6236_/X vssd1 vssd1 vccd1 vccd1 _6237_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__6691__C1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6168_ _6304_/A _7678_/B _5672_/A _6167_/Y _5715_/B vssd1 vssd1 vccd1 vccd1 _6168_/Y
+ sky130_fd_sc_hd__o221ai_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6038__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7235__A1 _6941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5119_ _5119_/A vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5246__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6099_ _6180_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6099_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5601__A _5601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7786__A2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5797__A1 _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5320__B _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8735__A1 _7825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7538__A2 _7512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8735__B2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8809_ _8808_/X _8547_/Y _8824_/S vssd1 vssd1 vccd1 vccd1 _8809_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7943__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5721__A1 _5738_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4887__A _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8359__A _8359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8671__B1 _8117_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput230 sports_i[0] vssd1 vssd1 vccd1 vccd1 _7779_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput241 sports_i[10] vssd1 vssd1 vccd1 vccd1 _7922_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__8806__B _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput252 sports_i[11] vssd1 vssd1 vccd1 vccd1 _7935_/A sky130_fd_sc_hd__buf_1
XANTENNA__7226__A1 _7683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput263 sports_i[12] vssd1 vssd1 vccd1 vccd1 _7948_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput274 sports_i[17] vssd1 vssd1 vccd1 vccd1 _8015_/A sky130_fd_sc_hd__buf_1
XANTENNA__5511__A _5511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput285 sports_i[27] vssd1 vssd1 vccd1 vccd1 _8175_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput296 sports_i[37] vssd1 vssd1 vccd1 vccd1 _7813_/B2 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5788__A1 _5788_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5788__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5230__B _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5657__S _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6342__A _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5470_ _5470_/A vssd1 vssd1 vccd1 vccd1 _5470_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4421_ _8160_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _5145_/A sky130_fd_sc_hd__nand2_8
Xoutput704 _6685_/X vssd1 vssd1 vccd1 vccd1 sports_o[77] sky130_fd_sc_hd__buf_12
XANTENNA__5712__A1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput715 _6778_/X vssd1 vssd1 vccd1 vccd1 sports_o[87] sky130_fd_sc_hd__buf_12
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput726 _6904_/X vssd1 vssd1 vccd1 vccd1 sports_o[97] sky130_fd_sc_hd__buf_12
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7140_ _5659_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7140_/X sky130_fd_sc_hd__a21o_1
X_4352_ hold41/A vssd1 vssd1 vccd1 vccd1 _4674_/C sky130_fd_sc_hd__inv_2
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5405__B _6646_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7465__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7071_ _7071_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7071_/X sky130_fd_sc_hd__and2_1
XANTENNA__5476__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6022_ _5274_/A _6089_/A1 _5275_/X input60/X vssd1 vssd1 vccd1 vccd1 _6022_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__8716__B _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7620__B _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5228__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7973_ _7777_/X _7972_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _7973_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__5779__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5779__B2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6924_ _6924_/A _7673_/B vssd1 vssd1 vccd1 vccd1 _6924_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6855_ _6002_/Y _6913_/B _6851_/Y _6853_/Y _6854_/Y vssd1 vssd1 vccd1 vccd1 _6856_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_147_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8451__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7348__A _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5806_ _5274_/X _5881_/A1 _5275_/X input52/X vssd1 vssd1 vccd1 vccd1 _5806_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6786_ _6968_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6786_/X sky130_fd_sc_hd__or2_2
XFILLER_0_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7940__A2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8525_ _8555_/A vssd1 vssd1 vccd1 vccd1 _8525_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5951__A1 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5737_ _5737_/A _6133_/B vssd1 vssd1 vccd1 vccd1 _5737_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8456_ _8455_/Y _8427_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8457_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5668_ _8140_/A _5690_/A _5667_/Y vssd1 vssd1 vccd1 vccd1 _5668_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7407_ _7701_/A _5239_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7409_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4619_ _8846_/A _8846_/B _8845_/B vssd1 vssd1 vccd1 vccd1 _4619_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__5703__A1 _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8387_ _8384_/X _8299_/X _8304_/X _8386_/X vssd1 vssd1 vccd1 vccd1 _8388_/A sky130_fd_sc_hd__a22o_1
X_5599_ _5596_/Y _4885_/A _5597_/Y _4890_/A _5598_/Y vssd1 vssd1 vccd1 vccd1 _5666_/C
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7338_ _7338_/A vssd1 vssd1 vccd1 vccd1 _7338_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6259__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7456__A1 _7105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7456__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7269_ _7269_/A vssd1 vssd1 vccd1 vccd1 _7269_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_110_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6719__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8184__A2 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7931__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8788__S _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5942__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7705__B _7705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7695__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7695__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5506__A _5506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5170__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8644__B1 _8009_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7998__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7960__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output514_A _6988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ _4975_/A _4868_/A _4976_/A _4870_/A _4969_/X vssd1 vssd1 vccd1 vccd1 _6461_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_116_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8271__B _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8175__A2 _6102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6640_ _6629_/Y _6511_/A _6630_/Y _6639_/X vssd1 vssd1 vccd1 vccd1 _6640_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5933__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6571_ _6567_/A _6510_/A _7380_/A _6512_/X vssd1 vssd1 vccd1 vccd1 _6571_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8310_ _8480_/B _8310_/B vssd1 vssd1 vccd1 vccd1 _8311_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_41_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5522_ _6024_/A _5745_/A vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__nor2_1
XANTENNA__7135__B1 _7134_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8241_ _8239_/Y _7954_/A _8240_/Y _7826_/A _7872_/A vssd1 vssd1 vccd1 vccd1 _8241_/X
+ sky130_fd_sc_hd__a221o_1
X_5453_ _5453_/A vssd1 vssd1 vccd1 vccd1 _5454_/B sky130_fd_sc_hd__inv_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput501 _7921_/X vssd1 vssd1 vccd1 vccd1 mports_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput512 _6984_/X vssd1 vssd1 vccd1 vccd1 sports_o[109] sky130_fd_sc_hd__buf_12
X_4404_ _4404_/A _8968_/Q vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__nand2_1
Xoutput523 _7346_/Y vssd1 vssd1 vccd1 vccd1 sports_o[119] sky130_fd_sc_hd__buf_12
XANTENNA__6894__C1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8172_ _8181_/A _8172_/B vssd1 vssd1 vccd1 vccd1 _8173_/A sky130_fd_sc_hd__nand2_1
Xoutput534 _7446_/X vssd1 vssd1 vccd1 vccd1 sports_o[129] sky130_fd_sc_hd__buf_12
XANTENNA__5161__A2 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput545 _7530_/X vssd1 vssd1 vccd1 vccd1 sports_o[139] sky130_fd_sc_hd__buf_12
X_5384_ _6024_/A vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput556 _7617_/Y vssd1 vssd1 vccd1 vccd1 sports_o[149] sky130_fd_sc_hd__buf_12
X_7123_ _5544_/X _7026_/X _7121_/X _7122_/X vssd1 vssd1 vccd1 vccd1 _7123_/X sky130_fd_sc_hd__o22a_1
Xoutput567 _7706_/Y vssd1 vssd1 vccd1 vccd1 sports_o[159] sky130_fd_sc_hd__buf_12
XANTENNA__7438__B2 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4335_ _4335_/A _7847_/A vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__nand2_1
Xoutput578 _7751_/Y vssd1 vssd1 vccd1 vccd1 sports_o[169] sky130_fd_sc_hd__buf_12
Xoutput589 _5203_/Y vssd1 vssd1 vccd1 vccd1 sports_o[179] sky130_fd_sc_hd__buf_12
X_7054_ _7272_/A _5150_/A _7138_/A vssd1 vssd1 vccd1 vccd1 _7054_/Y sky130_fd_sc_hd__o21ai_1
X_6005_ _6000_/X _8578_/B _6876_/A _6004_/X vssd1 vssd1 vccd1 vccd1 _6006_/A sky130_fd_sc_hd__a31o_2
XANTENNA__8954__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _7948_/Y _7769_/X _7949_/Y _6500_/X _7955_/Y vssd1 vssd1 vccd1 vccd1 _7956_/Y
+ sky130_fd_sc_hd__a221oi_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6628_/B _6905_/X _6906_/X vssd1 vssd1 vccd1 vccd1 _6907_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_38_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7887_ _6965_/A _7883_/Y _8163_/A _7884_/Y vssd1 vssd1 vccd1 vccd1 _7887_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6838_ _6807_/B _6837_/A _6724_/A _6837_/Y vssd1 vssd1 vccd1 vccd1 _6838_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7913__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6769_ _6760_/Y _6450_/X _6761_/Y _6762_/Y _6768_/X vssd1 vssd1 vccd1 vccd1 _6769_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8508_ _8567_/B _8107_/Y _8497_/S vssd1 vssd1 vccd1 vccd1 _8508_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8401__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8439_ _8439_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8439_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7017__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5152__A2 _5105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6101__A1 _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6101__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6652__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7062__C1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7601__A1 _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4966__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8157__A2 _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7904__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5915__A1 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6620__A _6620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8013__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8617__B1 _7903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7451__A _7451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8093__A1 _8093_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8093__B2 _7835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4794__B _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8977__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 mports_i[103] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5851__B1 _5846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7810_ _6500_/A _7813_/B2 _7813_/A2 _7769_/A vssd1 vssd1 vccd1 vccd1 _7810_/X sky130_fd_sc_hd__a22o_1
X_8790_ _8464_/A _8803_/B _8469_/A _8711_/X _8788_/S vssd1 vssd1 vccd1 vccd1 _8790_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5603__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8713__C _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7741_ _7740_/X _6358_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7742_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__buf_8
XANTENNA__6514__B _6514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8148__A2 _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6159__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4315__A _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7672_ _7672_/A _7723_/B vssd1 vssd1 vccd1 vccd1 _7672_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6159__B2 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4884_ _5129_/A vssd1 vssd1 vccd1 vccd1 _4885_/A sky130_fd_sc_hd__inv_6
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6623_ _7441_/B _6925_/B vssd1 vssd1 vccd1 vccd1 _6623_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5906__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7108__A0 _7107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6554_ _6551_/Y _6925_/B _6581_/A _6882_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6554_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5505_ _5505_/A vssd1 vssd1 vccd1 vccd1 _5505_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7345__B _7345_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7659__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6485_ _6484_/X _5064_/B _7000_/S vssd1 vssd1 vccd1 vccd1 _6485_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5146__A _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8224_ _7975_/X _8215_/X _8220_/X _8223_/X vssd1 vssd1 vccd1 vccd1 _8224_/X sky130_fd_sc_hd__a22o_2
XANTENNA__6790__A1_N _6511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5436_ _5436_/A vssd1 vssd1 vccd1 vccd1 _5436_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6331__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6331__B2 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8155_ _7975_/X _8137_/X _8149_/X _8154_/Y vssd1 vssd1 vccd1 vccd1 _8155_/X sky130_fd_sc_hd__a22o_2
X_5367_ _5367_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5367_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4985__A _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput375 _8744_/X vssd1 vssd1 vccd1 vccd1 mports_o[108] sky130_fd_sc_hd__buf_12
XANTENNA__5580__S _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput386 _8780_/X vssd1 vssd1 vccd1 vccd1 mports_o[118] sky130_fd_sc_hd__buf_12
Xoutput397 _8814_/X vssd1 vssd1 vccd1 vccd1 mports_o[128] sky130_fd_sc_hd__buf_12
X_7106_ _6648_/B _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7106_/X sky130_fd_sc_hd__a21o_1
X_4318_ _4337_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__nand2_1
X_8086_ _8093_/A1 _4946_/A _8093_/B1 _5119_/A vssd1 vssd1 vccd1 vccd1 _8086_/Y sky130_fd_sc_hd__o22ai_2
X_5298_ _5333_/B vssd1 vssd1 vccd1 vccd1 _7083_/A sky130_fd_sc_hd__inv_2
XANTENNA__7292__C1 _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7037_ _8919_/A _7037_/B vssd1 vssd1 vccd1 vccd1 _7037_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7831__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4645__A1 _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4645__B2 _4937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8387__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7044__C1 _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8192__A _8192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6398__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _7944_/A1 _5146_/A _7944_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _7939_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7898__A1 _7905_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6440__A _6440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4879__B _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4895__A _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6873__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7271__A _7271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8075__A1 _8080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6625__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5061__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7889__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7889__B2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8838__B1 _8249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8302__A2 hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ _6287_/A1 _4930_/X input7/X _4933_/A _6269_/X vssd1 vssd1 vccd1 vccd1 _7720_/B
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6313__A1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5221_ input91/X _8271_/B input28/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4324__B1 _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6864__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4875__A1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4875__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8066__A1 _8464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8066__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5152_ _6128_/B _5105_/A _5136_/A vssd1 vssd1 vccd1 vccd1 _5152_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6077__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7813__A1 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5083_ input87/X _8310_/B input25/X _4874_/X vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5824__B1 _5810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8911_ _4525_/B _8188_/S _8913_/A vssd1 vssd1 vccd1 vccd1 _8912_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8842_ _8845_/A _8842_/B vssd1 vssd1 vccd1 vccd1 _8842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8774__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8773_ _8771_/X _8725_/X _8772_/X _8442_/Y _8759_/Y vssd1 vssd1 vccd1 vccd1 _8773_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5985_ _5976_/X _5715_/B _6356_/S _5984_/X vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_94_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7724_ _6310_/X _7723_/B _7723_/Y vssd1 vssd1 vccd1 vccd1 _7724_/Y sky130_fd_sc_hd__o21ai_1
X_4936_ _8368_/A vssd1 vssd1 vccd1 vccd1 _8706_/B sky130_fd_sc_hd__buf_8
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8526__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_10 _7179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7655_ _7378_/X _6095_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7657_/B sky130_fd_sc_hd__o21ai_1
X_4867_ _4953_/A vssd1 vssd1 vccd1 vccd1 _4868_/A sky130_fd_sc_hd__buf_8
XFILLER_0_7_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8541__A2 _8145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7356__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6606_ _5336_/Y _6475_/X _5303_/Y _6851_/B vssd1 vssd1 vccd1 vccd1 _6606_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6552__A1 _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7586_ _6801_/B _7389_/A _6815_/B _7361_/X vssd1 vssd1 vccd1 vccd1 _7586_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4798_ _4798_/A _7511_/B vssd1 vssd1 vccd1 vccd1 _4799_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6552__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4699__B _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537_ _8842_/B _6535_/Y _6536_/X vssd1 vssd1 vccd1 vccd1 _6538_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5107__A2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6468_ _5019_/A _6549_/A _5024_/B _6876_/C _6968_/A vssd1 vssd1 vccd1 vccd1 _6468_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7501__B1 _7499_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8207_ _8203_/X _7954_/X _8206_/X _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8207_/X
+ sky130_fd_sc_hd__a221o_1
X_5419_ input98/X _4871_/A input36/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6855__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6399_ _6202_/B _7754_/B _6398_/X vssd1 vssd1 vccd1 vccd1 _6399_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8057__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8138_ _8150_/B vssd1 vssd1 vccd1 vccd1 _8146_/B sky130_fd_sc_hd__inv_2
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6068__B1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6419__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7804__A1 _7803_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6607__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8069_ _7777_/X _8068_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _8069_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__7030__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6154__B _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5043__A1 _5064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6240__B1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5043__B2 _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8780__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5594__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6791__A1 _6786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5993__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8532__A2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6170__A _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5503__C1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5514__A _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8048__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6329__B _6375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8599__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output427_A _8242_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5806__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7559__B1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8756__C1 _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8220__A1 _8217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8220__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5034__A1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6064__B _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5034__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5722_/A _5111_/A _5723_/A _4931_/A _5769_/X vssd1 vssd1 vccd1 vccd1 _5770_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _8239_/A _4721_/B vssd1 vssd1 vccd1 vccd1 _4722_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6080__A _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7440_ _7438_/X _7640_/B _5381_/X _7680_/B _7439_/Y vssd1 vssd1 vccd1 vccd1 _7440_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4652_ _5116_/A vssd1 vssd1 vccd1 vccd1 _6941_/A sky130_fd_sc_hd__inv_4
XFILLER_0_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput30 mports_i[126] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5408__B _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput41 mports_i[136] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7371_ _7701_/A _5159_/A _6264_/X vssd1 vssd1 vccd1 vccd1 _7376_/B sky130_fd_sc_hd__o21ai_1
Xinput52 mports_i[146] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4583_ _4818_/B _4909_/A vssd1 vssd1 vccd1 vccd1 _4583_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4312__B _4312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput63 mports_i[156] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput74 mports_i[166] vssd1 vssd1 vccd1 vccd1 _4810_/B sky130_fd_sc_hd__buf_6
X_6322_ _6593_/A _6322_/B vssd1 vssd1 vccd1 vccd1 _6322_/X sky130_fd_sc_hd__or2_1
XANTENNA__8287__A1 _7807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput85 mports_i[176] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_2
Xinput96 mports_i[186] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6253_ _6253_/A vssd1 vssd1 vccd1 vccd1 _6253_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5424__A _5425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5204_ input90/X _4934_/A input27/X _4937_/A vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8944__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6184_ _6941_/B _6626_/B vssd1 vssd1 vccd1 vccd1 _6184_/Y sky130_fd_sc_hd__nand2_1
X_5135_ _6233_/B _6499_/A _5128_/Y _6497_/B _6202_/B vssd1 vssd1 vccd1 vccd1 _5135_/Y
+ sky130_fd_sc_hd__o221ai_1
XANTENNA__7798__B1 _7803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7262__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ _5066_/A _5136_/A vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__and2_1
XANTENNA__8454__B _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7014__A2 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8825_ _8824_/X _8200_/X _8829_/S vssd1 vssd1 vccd1 vccd1 _8826_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_67_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6222__B1 _6221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5968_ _5965_/Y _4885_/A _5966_/Y _4890_/A _5967_/Y vssd1 vssd1 vccd1 vccd1 _5993_/C
+ sky130_fd_sc_hd__o221a_2
X_8756_ _7929_/Y _8711_/A _8396_/X _8770_/B _8824_/S vssd1 vssd1 vccd1 vccd1 _8756_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7970__B1 _7969_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4919_ input1/X _8516_/B _4888_/A _4913_/X _4918_/X vssd1 vssd1 vccd1 vccd1 _4919_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7707_ _8716_/A _7707_/B _7707_/C _7707_/D vssd1 vssd1 vccd1 vccd1 _7707_/X sky130_fd_sc_hd__or4_1
X_8687_ _8684_/X _8590_/X _8685_/Y _8686_/X vssd1 vssd1 vccd1 vccd1 _8687_/X sky130_fd_sc_hd__a31o_1
X_5899_ _5899_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _7607_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_152_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8514__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7638_ _7638_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _7640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_118_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _8976_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7722__B1 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5318__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7569_ _7167_/A _7349_/A _6779_/Y _7680_/B _7568_/Y vssd1 vssd1 vccd1 vccd1 _7569_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8278__A1 _7784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6289__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5500__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6149__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7789__B1 _7788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7253__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8450__A1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8202__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6213__B1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5016__B2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8753__A2 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5509__A _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output377_A _7934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5943__S _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__B _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output711_A _6735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8555__A _8555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__A1 _5272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6940_ _6940_/A vssd1 vssd1 vccd1 vccd1 _6940_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6075__A _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6871_ _6871_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6871_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8744__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5822_ _5031_/X _5772_/X _5820_/Y _5821_/X vssd1 vssd1 vccd1 vccd1 _5822_/X sky130_fd_sc_hd__a22o_2
X_8610_ _7869_/Y _8581_/X _7871_/Y _8583_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8610_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8290__A _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5558__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7952__B1 _7958_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8541_ _4894_/A _8145_/Y _4891_/X _8187_/X _8540_/Y vssd1 vssd1 vccd1 vccd1 _8803_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5753_ _6711_/S _5751_/X _5752_/X vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4704_ _4693_/A _4693_/B _4713_/A vssd1 vssd1 vccd1 vccd1 _4705_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8472_ _8471_/Y _8578_/B hold36/A _4727_/C _8496_/S vssd1 vssd1 vccd1 vccd1 _8472_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5684_ _5619_/X _5735_/B _6593_/A vssd1 vssd1 vccd1 vccd1 _5684_/X sky130_fd_sc_hd__mux2_1
X_7423_ _5308_/X _7680_/B _7421_/X _7348_/A _7422_/X vssd1 vssd1 vccd1 vccd1 _7423_/X
+ sky130_fd_sc_hd__a221o_1
X_4635_ _4635_/A _4635_/B vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6527__A1_N _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7354_ _5150_/A _7640_/B _7349_/Y _6514_/B vssd1 vssd1 vccd1 vccd1 _7354_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__inv_2
XFILLER_0_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4977__B _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6305_ _6303_/Y _7629_/B _5171_/B _6304_/Y vssd1 vssd1 vccd1 vccd1 _6305_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7285_ _7284_/X _7746_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__mux2_4
X_4497_ _7384_/A vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__inv_2
X_6236_ _6233_/Y _6202_/B _6234_/Y _6235_/Y vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5494__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6691__B1 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6167_ _6166_/B _6123_/Y _6166_/Y vssd1 vssd1 vccd1 vccd1 _6167_/Y sky130_fd_sc_hd__o21ai_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8432__A1 _8782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5237_/A vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__clkinv_4
X_6098_ _6141_/A1 _5102_/A _6141_/B1 _5191_/A _6097_/X vssd1 vssd1 vccd1 vccd1 _6180_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5246__A1 _6566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5246__B2 _5248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5049_ _5046_/Y _8455_/B _5047_/Y _4891_/X _5048_/Y vssd1 vssd1 vccd1 vccd1 _5050_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8735__A2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8808_ _8551_/A _8738_/Y _8712_/A _8549_/X vssd1 vssd1 vccd1 vccd1 _8808_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_137_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7943__B1 _7942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5954__C1 _5953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8739_ _8755_/A _7856_/A _7851_/A _8738_/Y _8782_/A vssd1 vssd1 vccd1 vccd1 _8739_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7544__A _7544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5182__B1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5721__A2 _5827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8359__B _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8120__B1 _8111_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5064__A _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8671__A1 _8510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8671__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6682__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput220 mports_i[92] vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__buf_2
XANTENNA__8375__A _8375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput231 sports_i[100] vssd1 vssd1 vccd1 vccd1 _4658_/A sky130_fd_sc_hd__clkbuf_8
Xinput242 sports_i[110] vssd1 vssd1 vccd1 vccd1 _7905_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput253 sports_i[120] vssd1 vssd1 vccd1 vccd1 _8028_/A sky130_fd_sc_hd__clkbuf_2
Xinput264 sports_i[130] vssd1 vssd1 vccd1 vccd1 _8192_/A sky130_fd_sc_hd__clkbuf_4
Xinput275 sports_i[18] vssd1 vssd1 vccd1 vccd1 _8030_/A sky130_fd_sc_hd__buf_1
Xinput286 sports_i[28] vssd1 vssd1 vccd1 vccd1 _8189_/C sky130_fd_sc_hd__clkbuf_4
Xinput297 sports_i[38] vssd1 vssd1 vccd1 vccd1 _7818_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5788__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6985__A1 _6349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6985__B2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4996__A0 _4993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8726__A2 _8317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6342__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5239__A _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7162__A1 _6758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7162__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4420_ _4420_/A _4443_/A vssd1 vssd1 vccd1 vccd1 _4420_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_151_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput705 _6692_/X vssd1 vssd1 vccd1 vccd1 sports_o[78] sky130_fd_sc_hd__buf_12
Xoutput716 _6791_/X vssd1 vssd1 vccd1 vccd1 sports_o[88] sky130_fd_sc_hd__buf_12
Xoutput727 _6918_/Y vssd1 vssd1 vccd1 vccd1 sports_o[98] sky130_fd_sc_hd__buf_12
XFILLER_0_111_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4351_ _4800_/B hold26/A vssd1 vssd1 vccd1 vccd1 _4351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8662__A1 _8081_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7070_ _5218_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7070_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7465__A2 _5464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5476__A1 _7524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6021_ _6021_/A vssd1 vssd1 vccd1 vccd1 _6021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6673__B1 _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5476__B2 _6727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5228__A1 _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5228__B2 _6566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7972_ _7962_/Y _7874_/X _7963_/Y _7875_/X _7971_/Y vssd1 vssd1 vccd1 vccd1 _7972_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5779__A2 _5744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6976__B2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6923_ _6968_/A _6923_/B vssd1 vssd1 vccd1 vccd1 _6923_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6854_ _6854_/A _6854_/B vssd1 vssd1 vccd1 vccd1 _6854_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5805_ _5805_/A vssd1 vssd1 vccd1 vccd1 _5805_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_91_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6785_ _5827_/A _6841_/A _6779_/Y _6854_/A _6784_/Y vssd1 vssd1 vccd1 vccd1 _6786_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5149__A _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8524_ _8523_/Y _8499_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8555_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5736_ _6547_/A _5781_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5737_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8455_ _8455_/A _8455_/B vssd1 vssd1 vccd1 vccd1 _8455_/Y sky130_fd_sc_hd__nand2_1
X_5667_ _5667_/A vssd1 vssd1 vccd1 vccd1 _5667_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7364__A _7364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5164__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4618_ _4618_/A _4658_/A vssd1 vssd1 vccd1 vccd1 _8845_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7406_ _5248_/A _7696_/B _6597_/B _7361_/X _7405_/Y vssd1 vssd1 vccd1 vccd1 _7406_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8386_ _4894_/A _8351_/A _4891_/X _8404_/A _8385_/X vssd1 vssd1 vccd1 vccd1 _8386_/X
+ sky130_fd_sc_hd__o221a_2
X_5598_ _5274_/A _5637_/A1 _5275_/A input44/X vssd1 vssd1 vccd1 vccd1 _5598_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_142_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7083__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7337_ _7336_/X _5028_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7338_/A sky130_fd_sc_hd__mux2_1
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__inv_2
XANTENNA__4500__B _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7268_ _6337_/X _7138_/A _7267_/X vssd1 vssd1 vccd1 vccd1 _7269_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__8653__A1 _8439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7456__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5467__A1 _5543_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5467__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6664__B1 _6657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6219_ _5741_/B _6185_/A _6218_/Y _5125_/X vssd1 vssd1 vccd1 vccd1 _6219_/X sky130_fd_sc_hd__a22o_1
X_7199_ _7198_/X _5923_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7200_/A sky130_fd_sc_hd__mux2_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6967__A1 _6277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6967__B2 _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7392__A1 _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7144__A1 _7524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7144__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5155__B1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7695__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4410__B _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8644__A1 _8416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8644__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5458__A1 _7459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5522__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output507_A _6960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4969__B1 _4977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6072__B _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6570_ _6568_/X _6628_/B _6569_/Y vssd1 vssd1 vccd1 vccd1 _7380_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__5933__A2 _6007_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5521_ _5518_/Y _4885_/A _5519_/Y _4890_/A _5520_/Y vssd1 vssd1 vccd1 vccd1 _5745_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7135__A1 _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6800__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8240_ _8240_/A vssd1 vssd1 vccd1 vccd1 _8240_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5452_ _6644_/A _5451_/X _6793_/S vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8883__A1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6343__C1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5697__A1 _5697_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput502 _7018_/X vssd1 vssd1 vccd1 vccd1 sports_o[0] sky130_fd_sc_hd__buf_12
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5697__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput513 _7074_/X vssd1 vssd1 vccd1 vccd1 sports_o[10] sky130_fd_sc_hd__buf_12
X_4403_ _8239_/A _6024_/A _4412_/C vssd1 vssd1 vccd1 vccd1 _4404_/A sky130_fd_sc_hd__nand3_1
XANTENNA__6894__B1 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8171_ _8181_/A _8171_/B vssd1 vssd1 vccd1 vccd1 _8171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput524 _7078_/X vssd1 vssd1 vccd1 vccd1 sports_o[11] sky130_fd_sc_hd__buf_12
X_5383_ _5383_/A vssd1 vssd1 vccd1 vccd1 _6633_/A sky130_fd_sc_hd__inv_2
XANTENNA__4320__B _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput535 _7082_/X vssd1 vssd1 vccd1 vccd1 sports_o[12] sky130_fd_sc_hd__buf_12
Xoutput546 _7087_/X vssd1 vssd1 vccd1 vccd1 sports_o[13] sky130_fd_sc_hd__buf_12
Xoutput557 _7093_/X vssd1 vssd1 vccd1 vccd1 sports_o[14] sky130_fd_sc_hd__buf_12
X_7122_ _6679_/B _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7122_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8635__A1 _8375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput568 _7098_/X vssd1 vssd1 vccd1 vccd1 sports_o[15] sky130_fd_sc_hd__buf_12
XANTENNA__7438__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4334_ _4334_/A _4334_/B vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__nand2_1
Xoutput579 _7104_/X vssd1 vssd1 vccd1 vccd1 sports_o[16] sky130_fd_sc_hd__buf_12
XFILLER_0_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5449__A1 _5497_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5449__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7053_ _7053_/A vssd1 vssd1 vccd1 vccd1 _7053_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6528__A _6528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6004_ _5845_/B _6002_/Y _5997_/Y _6003_/X vssd1 vssd1 vccd1 vccd1 _6004_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5151__B _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6962__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6949__A1 _7705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7955_ _7958_/A1 _5780_/X _7958_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7955_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_49_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5621__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7359__A _7359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5621__B2 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6906_ _6906_/A _6906_/B vssd1 vssd1 vccd1 vccd1 _6906_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7886_ _7881_/Y _6059_/B _7882_/Y _5359_/B _7885_/X vssd1 vssd1 vccd1 vccd1 _7886_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6837_ _6837_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6837_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_147_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6768_ _5770_/X _6510_/A _6767_/Y _6512_/X vssd1 vssd1 vccd1 vccd1 _6768_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8507_ _8104_/Y _8299_/X _8506_/Y _8304_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8507_/X
+ sky130_fd_sc_hd__a221o_1
X_5719_ _5685_/A _4931_/A _5686_/A _5111_/A _5718_/X vssd1 vssd1 vccd1 vccd1 _5741_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7126__A1 _5500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6699_ _6699_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6699_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7126__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7094__A _7094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5137__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8438_ _8438_/A vssd1 vssd1 vccd1 vccd1 _8438_/X sky130_fd_sc_hd__buf_1
XFILLER_0_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5688__B2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6885__B1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8369_ _8369_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8369_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7822__A _7829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7429__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8626__A1 _8372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6101__A2 _4909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7062__B1 _5161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7601__A2 _5899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5612__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6173__A _7696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7365__A1 _5161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6168__A2 _7678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8562__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7365__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6901__A _7660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7117__A1 _5498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6620__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8314__B1 _8313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4421__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output457_A _7863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8617__A1 _7901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8617__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7451__B _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8093__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5851__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 mports_i[104] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8250__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5603__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7740_ _6355_/X _7754_/A _7739_/X vssd1 vssd1 vccd1 vccd1 _7740_/X sky130_fd_sc_hd__o21a_1
X_4952_ _4952_/A vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__buf_1
XANTENNA__8969__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4883_ input1/X vssd1 vssd1 vccd1 vccd1 _4883_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6159__A2 _6174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7671_ _6913_/A _7542_/A _7694_/A _6119_/Y _7670_/Y vssd1 vssd1 vccd1 vccd1 _7672_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_129_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6622_ _6622_/A vssd1 vssd1 vccd1 vccd1 _7441_/B sky130_fd_sc_hd__inv_2
XANTENNA__6811__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6553_ _6553_/A vssd1 vssd1 vccd1 vccd1 _6581_/A sky130_fd_sc_hd__inv_2
XANTENNA__7108__A1 _5460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8305__B1 _8303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7118__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5504_ _6669_/B vssd1 vssd1 vccd1 vccd1 _7115_/A sky130_fd_sc_hd__inv_2
X_6484_ _6899_/B _6480_/X _6483_/X vssd1 vssd1 vccd1 vccd1 _6484_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7659__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5146__B _6514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5435_ _5435_/A vssd1 vssd1 vccd1 vccd1 _5435_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_113_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8223_ _7777_/A _8222_/X _7792_/A vssd1 vssd1 vccd1 vccd1 _8223_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_42_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5366_ _5337_/A _5111_/A _5338_/A _4931_/A _5365_/X vssd1 vssd1 vccd1 vccd1 _5367_/A
+ sky130_fd_sc_hd__o221a_4
X_8154_ _8153_/X _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _8154_/Y sky130_fd_sc_hd__a21oi_1
Xoutput376 _8748_/X vssd1 vssd1 vccd1 vccd1 mports_o[109] sky130_fd_sc_hd__buf_12
XFILLER_0_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput387 _8783_/X vssd1 vssd1 vccd1 vccd1 mports_o[119] sky130_fd_sc_hd__buf_12
X_7105_ _7105_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7105_/X sky130_fd_sc_hd__and2_1
X_4317_ _7847_/A _4658_/A vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__nand2_1
Xoutput398 _8818_/X vssd1 vssd1 vccd1 vccd1 mports_o[129] sky130_fd_sc_hd__buf_12
X_8085_ _8085_/A vssd1 vssd1 vccd1 vccd1 _8085_/Y sky130_fd_sc_hd__inv_2
X_5297_ _5294_/Y _4886_/A _5295_/Y _4891_/A _5296_/Y vssd1 vssd1 vccd1 vccd1 _7432_/B
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5162__A _7304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7036_ _7036_/A vssd1 vssd1 vccd1 vccd1 _7036_/X sky130_fd_sc_hd__buf_1
XANTENNA__7831__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4645__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8241__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8192__B _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6398__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7595__B2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7089__A _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7938_ _7935_/Y _7013_/A _7936_/Y _5117_/A _7937_/Y vssd1 vssd1 vccd1 vccd1 _8376_/A
+ sky130_fd_sc_hd__a221oi_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7869_ _7864_/Y _6965_/A _7865_/Y _8163_/A _7868_/Y vssd1 vssd1 vccd1 vccd1 _7869_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7817__A _7829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7536__B _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6440__B _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6570__A2 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5337__A _5337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5530__B1 _5511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8075__A2 _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__A1 _6089_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7586__A1 _6801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7586__B2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__B1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6010__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6561__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8838__A1 _8247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8838__B2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4572__B2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8944__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5220_ _5217_/X _6233_/B _6170_/A _5219_/Y vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4324__A1 _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4875__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5151_ _6544_/A _6234_/B vssd1 vssd1 vccd1 vccd1 _5151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_138_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8066__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6077__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6077__B2 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5082_ _5131_/A2 _8480_/B _5131_/B2 _4870_/X _5081_/X vssd1 vssd1 vccd1 vccd1 _6499_/A
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__7813__A2 _7813_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5824__A1 _5809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5824__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8910_ _8910_/A vssd1 vssd1 vccd1 vccd1 _8949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8841_ _4593_/Y _4828_/Y _4619_/Y vssd1 vssd1 vccd1 vccd1 _8855_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6525__B _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4326__A _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8772_ _8782_/A _8772_/B vssd1 vssd1 vccd1 vccd1 _8772_/X sky130_fd_sc_hd__or2_1
X_5984_ _6084_/B _6841_/B _7623_/B _5096_/A vssd1 vssd1 vccd1 vccd1 _5984_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7723_ _7723_/A _7723_/B vssd1 vssd1 vccd1 vccd1 _7723_/Y sky130_fd_sc_hd__nand2_1
X_4935_ _4935_/A vssd1 vssd1 vccd1 vccd1 _8368_/A sky130_fd_sc_hd__buf_12
XFILLER_0_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8526__B1 _8130_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7637__A _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 _7179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7654_ _7648_/X _7651_/X _7652_/X _7653_/X vssd1 vssd1 vccd1 vccd1 _7654_/X sky130_fd_sc_hd__a31o_2
X_4866_ _4866_/A vssd1 vssd1 vccd1 vccd1 _8944_/D sky130_fd_sc_hd__inv_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6605_ _5362_/A _6429_/S _6603_/X _6604_/X vssd1 vssd1 vccd1 vccd1 _6605_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7356__B _7356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4797_ _4821_/A vssd1 vssd1 vccd1 vccd1 _7511_/B sky130_fd_sc_hd__inv_2
XANTENNA__6552__A2 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7585_ _7542_/A _5879_/A _7326_/A vssd1 vssd1 vccd1 vccd1 _7585_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_132_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5157__A _5359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8829__A1 _8215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6536_ _8194_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _6536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6467_ _6517_/B vssd1 vssd1 vccd1 vccd1 _6467_/X sky130_fd_sc_hd__buf_8
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7501__B2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7372__A _7372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8206_ _8210_/A1 _6544_/B _8210_/B1 _4518_/A _8205_/X vssd1 vssd1 vccd1 vccd1 _8206_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5512__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5418_ _5440_/A _4868_/A _5441_/A _5089_/A _5417_/X vssd1 vssd1 vccd1 vccd1 _5465_/A
+ sky130_fd_sc_hd__o221a_4
X_6398_ _7753_/A _6234_/B _6397_/X _5128_/A _6386_/S vssd1 vssd1 vccd1 vccd1 _6398_/X
+ sky130_fd_sc_hd__a221o_1
X_5349_ input96/X _5192_/X input33/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8057__A2 _8451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8137_ _8148_/A1 _6626_/B _8142_/A _6941_/A _8136_/X vssd1 vssd1 vccd1 vccd1 _8137_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6068__A1 _6136_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6068__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7804__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8068_ _8058_/Y _7874_/X _8059_/Y _7875_/X _8067_/Y vssd1 vssd1 vccd1 vccd1 _8068_/Y
+ sky130_fd_sc_hd__a221oi_4
X_7019_ _7059_/A vssd1 vssd1 vccd1 vccd1 _7019_/X sky130_fd_sc_hd__buf_8
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5043__A2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6240__A1 _6247_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6240__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6791__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5766__S _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5993__C _5993_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7266__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8967__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8296__A2 _7803_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5514__B _7120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8048__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5806__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6626__A _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7221__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7559__A1 _6758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6345__B _6375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5034__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8508__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7548__A1_N _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4720_/A _7272_/B vssd1 vssd1 vccd1 vccd1 _4721_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5990__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4651_ hold44/A _8198_/A vssd1 vssd1 vccd1 vccd1 _5116_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6080__B _6897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7731__B2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 mports_i[117] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput31 mports_i[127] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
X_4582_ _8284_/A vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__clkinv_4
X_7370_ _7510_/B vssd1 vssd1 vccd1 vccd1 _7701_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__5742__B1 _5739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 mports_i[137] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 mports_i[147] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput64 mports_i[157] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_2
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput75 mports_i[167] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_2
X_6321_ _6321_/A _8189_/A vssd1 vssd1 vccd1 vccd1 _6321_/Y sky130_fd_sc_hd__nand2_1
Xinput86 mports_i[177] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_2
XFILLER_0_141_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8288__A _8288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 mports_i[187] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6298__A1 _7729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6252_ _6253_/A _8480_/B input6/X _4870_/X _6251_/X vssd1 vssd1 vccd1 vccd1 _6252_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__6298__B2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7495__B1 _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5203_ _6266_/A _6536_/B _5159_/Y _5202_/X vssd1 vssd1 vccd1 vccd1 _5203_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6183_ _6183_/A1 _4929_/A input3/X _4932_/A _6182_/X vssd1 vssd1 vccd1 vccd1 _6941_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7247__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5134_ _6261_/A vssd1 vssd1 vccd1 vccd1 _6202_/B sky130_fd_sc_hd__buf_4
XANTENNA__7798__A1 _4566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7798__B2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5065_ _6359_/S vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__inv_4
XANTENNA__6536__A _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5440__A _5440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8824_ _8823_/X _8211_/A _8824_/S vssd1 vssd1 vccd1 vccd1 _8824_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6222__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6222__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8755_ _8755_/A _8755_/B _8755_/C vssd1 vssd1 vccd1 vccd1 _8770_/B sky130_fd_sc_hd__and3_2
X_5967_ _5274_/A _6031_/A1 _5275_/A input58/X vssd1 vssd1 vccd1 vccd1 _5967_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5586__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7970__A1 _8404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6773__A2 _6770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7970__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7706_ _7704_/Y _7332_/A _7705_/Y vssd1 vssd1 vccd1 vccd1 _7706_/Y sky130_fd_sc_hd__a21oi_2
X_4918_ input80/X _8716_/B input17/X _4917_/X vssd1 vssd1 vccd1 vccd1 _4918_/X sky130_fd_sc_hd__o22a_1
X_8686_ _8821_/A _8686_/B vssd1 vssd1 vccd1 vccd1 _8686_/X sky130_fd_sc_hd__and2_1
XFILLER_0_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _5924_/A vssd1 vssd1 vccd1 vccd1 _5898_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_117_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7637_ _7694_/A _7637_/B vssd1 vssd1 vccd1 vccd1 _7637_/X sky130_fd_sc_hd__or2_1
X_4849_ _8953_/D vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__inv_2
XANTENNA__7722__A1 _7349_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5733__B1 _5723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7568_ _7686_/A _7568_/B vssd1 vssd1 vccd1 vccd1 _7568_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6519_ _6506_/A _5105_/A _6449_/A vssd1 vssd1 vccd1 vccd1 _6519_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7499_ _5584_/B _7753_/B _7497_/Y _7498_/Y vssd1 vssd1 vccd1 vccd1 _7499_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6289__A1 _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5615__A _7304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7789__A1 _7786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7789__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7041__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4472__B1 _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8202__A2 _8209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6213__A1 _6229_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5016__A2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6213__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7961__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4775__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5509__B _5549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4413__B _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7713__A1 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5724__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7216__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5488__C1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8555__B _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output704_A _6685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5260__A _7413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6452__A1 _4966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8729__B1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6870_ _7604_/B _6869_/X _6870_/S vssd1 vssd1 vccd1 vccd1 _6871_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6204__A1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5821_ _6202_/B _6770_/A _5136_/X vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__o21a_1
XANTENNA__8290__B _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7952__A1 _7958_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7187__A _7187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8540_ _8540_/A _8755_/B vssd1 vssd1 vccd1 vccd1 _8540_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4766__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5963__B1 _5937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5752_ _6166_/B _5752_/B vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ _4733_/B vssd1 vssd1 vccd1 vccd1 _4725_/A sky130_fd_sc_hd__inv_2
XFILLER_0_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8471_ _8471_/A vssd1 vssd1 vccd1 vccd1 _8471_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7704__A1 _6207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5683_ _8189_/A _7542_/B _5682_/Y vssd1 vssd1 vccd1 vccd1 _5735_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__8901__B1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7422_ _7422_/A _7660_/B vssd1 vssd1 vccd1 vccd1 _7422_/X sky130_fd_sc_hd__and2_1
XFILLER_0_60_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4634_ _4634_/A _8967_/D vssd1 vssd1 vccd1 vccd1 _4635_/B sky130_fd_sc_hd__or2_1
XFILLER_0_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4565_ _8181_/A _7707_/C vssd1 vssd1 vccd1 vccd1 _7311_/A sky130_fd_sc_hd__nor2_8
X_7353_ _7351_/X _7332_/A _7352_/Y vssd1 vssd1 vccd1 vccd1 _7353_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5435__A _5435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6304_ _6304_/A _6965_/B vssd1 vssd1 vccd1 vccd1 _6304_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__8665__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7284_ _6364_/X _7138_/X _7282_/X _7283_/X vssd1 vssd1 vccd1 vccd1 _7284_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4496_ _8240_/A _4436_/A _4495_/Y _4460_/B vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6140__B1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6235_ _6128_/B _6207_/A _5136_/X vssd1 vssd1 vccd1 vccd1 _6235_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__8680__A2 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7650__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5494__A2 _5464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6691__A1 _5558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/A _6166_/B vssd1 vssd1 vccd1 vccd1 _6166_/Y sky130_fd_sc_hd__nand2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5117_/A vssd1 vssd1 vccd1 vccd1 _8857_/B sky130_fd_sc_hd__buf_12
X_6097_ _6140_/A1 _5192_/A input63/X _5193_/A vssd1 vssd1 vccd1 vccd1 _6097_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5246__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5048_ _4893_/A input84/X _4896_/A input21/X vssd1 vssd1 vccd1 vccd1 _5048_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8196__A1 _8189_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8196__B2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8807_ _8829_/S _8805_/X _8806_/Y vssd1 vssd1 vccd1 vccd1 _8807_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_83_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6713__B _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6999_ _6395_/A _6994_/B _6397_/X _6989_/B vssd1 vssd1 vccd1 vccd1 _6999_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7943__A1 _8351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7943__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8738_ _8738_/A vssd1 vssd1 vccd1 vccd1 _8738_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5954__B1 _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5329__B _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8669_ _8698_/B _8107_/Y _8590_/X vssd1 vssd1 vccd1 vccd1 _8669_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7544__B _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5182__A1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5182__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8120__B2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5064__B _5064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8671__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6682__A1 _5498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5999__B _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6682__B2 _5544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput210 mports_i[83] vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__8375__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput221 mports_i[93] vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__buf_2
Xinput232 sports_i[101] vssd1 vssd1 vccd1 vccd1 _8252_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput243 sports_i[111] vssd1 vssd1 vccd1 vccd1 _7918_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput254 sports_i[121] vssd1 vssd1 vccd1 vccd1 _8054_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__6176__A _6212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput265 sports_i[131] vssd1 vssd1 vccd1 vccd1 _8209_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5080__A _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput276 sports_i[19] vssd1 vssd1 vccd1 vccd1 _8045_/A sky130_fd_sc_hd__buf_1
Xinput287 sports_i[29] vssd1 vssd1 vccd1 vccd1 _8210_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__7631__B1 _7385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput298 sports_i[39] vssd1 vssd1 vccd1 vccd1 _7859_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__6985__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4408__B _4408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4996__A1 _7332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8187__A1 _8189_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7934__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6623__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6342__C _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7162__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6370__B1 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput706 _6703_/X vssd1 vssd1 vccd1 vccd1 sports_o[79] sky130_fd_sc_hd__buf_12
Xoutput717 _6806_/X vssd1 vssd1 vccd1 vccd1 sports_o[89] sky130_fd_sc_hd__buf_12
X_4350_ _8512_/S _4810_/B vssd1 vssd1 vccd1 vccd1 _4350_/Y sky130_fd_sc_hd__nand2_1
Xoutput728 _6930_/X vssd1 vssd1 vccd1 vccd1 sports_o[99] sky130_fd_sc_hd__buf_12
XFILLER_0_50_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7470__A _7470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5476__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6020_ _6020_/A vssd1 vssd1 vccd1 vccd1 _6020_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7870__B1 _7877_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5702__B _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5228__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7971_ _7971_/A1 _7876_/X _7971_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7971_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__4318__B _4318_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6976__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6922_ _6115_/A _6841_/A _6119_/Y _6854_/A _6921_/X vssd1 vssd1 vccd1 vccd1 _6923_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7629__B _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6853_ _6432_/X _6852_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6853_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6728__A2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5804_ _5804_/A vssd1 vssd1 vccd1 vccd1 _5804_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6025__S _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6784_ _6784_/A _6784_/B vssd1 vssd1 vccd1 vccd1 _6784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8523_ _8523_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8523_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5735_ _6875_/B _5735_/B vssd1 vssd1 vccd1 vccd1 _5735_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8454_ _8454_/A _8555_/B vssd1 vssd1 vccd1 vccd1 _8454_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5666_ _8160_/A _6231_/C _5666_/C vssd1 vssd1 vccd1 vccd1 _5667_/A sky130_fd_sc_hd__or3_1
XFILLER_0_5_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5164__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7405_ _6594_/Y _7680_/B _7403_/X _7404_/Y vssd1 vssd1 vccd1 vccd1 _7405_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_0_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4617_ _4617_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6361__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8385_ _8300_/B _8352_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8385_/X sky130_fd_sc_hd__o21a_1
X_5597_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5597_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7336_ _5000_/X _7754_/A _7335_/X vssd1 vssd1 vccd1 vccd1 _7336_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_102_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4548_ hold1/X vssd1 vssd1 vccd1 vccd1 _4837_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8102__B2 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6113__B1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7267_ _6333_/Y _7088_/A _7266_/X _7059_/A _7089_/A vssd1 vssd1 vccd1 vccd1 _7267_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8476__A _8476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8653__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4479_ _4518_/A vssd1 vssd1 vccd1 vccd1 _6500_/A sky130_fd_sc_hd__inv_12
XANTENNA__5467__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6664__A1 _5464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6218_ _6628_/B _6216_/X _6217_/Y vssd1 vssd1 vccd1 vccd1 _6218_/Y sky130_fd_sc_hd__a21oi_1
X_7198_ _6868_/A _7023_/X _7197_/X vssd1 vssd1 vccd1 vccd1 _7198_/X sky130_fd_sc_hd__o21a_1
X_6149_ _6937_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6149_/Y sky130_fd_sc_hd__nand2_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6416__A1 _4876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6416__B2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6967__A2 _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6724__A _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6443__B _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6719__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7916__B2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7144__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5155__A1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5155__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5075__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8644__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5803__A _5803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6655__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7080__A1 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4969__A1 _4978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4969__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6634__A _6634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7907__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5684__S _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5520_ _5274_/A _5764_/A1 _5275_/A input48/X vssd1 vssd1 vccd1 vccd1 _5520_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8332__A1 _8346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7135__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5451_ _5465_/A _5077_/A _6017_/A _6671_/B vssd1 vssd1 vccd1 vccd1 _5451_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6343__B1 _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4601__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5697__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput503 _6936_/X vssd1 vssd1 vccd1 vccd1 sports_o[100] sky130_fd_sc_hd__buf_12
X_4402_ _4402_/A vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__buf_12
XANTENNA__6894__A1 _6107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8170_ _7768_/X _8165_/Y _8169_/Y _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8170_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput514 _6988_/X vssd1 vssd1 vccd1 vccd1 sports_o[110] sky130_fd_sc_hd__buf_12
X_5382_ _6875_/B _5308_/B _5381_/X vssd1 vssd1 vccd1 vccd1 _5383_/A sky130_fd_sc_hd__o21ai_1
Xoutput525 _7353_/Y vssd1 vssd1 vccd1 vccd1 sports_o[120] sky130_fd_sc_hd__buf_12
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput536 _7455_/X vssd1 vssd1 vccd1 vccd1 sports_o[130] sky130_fd_sc_hd__buf_12
XFILLER_0_50_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7121_ _7121_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7121_/X sky130_fd_sc_hd__and2_1
Xoutput547 _7540_/Y vssd1 vssd1 vccd1 vccd1 sports_o[140] sky130_fd_sc_hd__buf_12
X_4333_ _4333_/A _6231_/C vssd1 vssd1 vccd1 vccd1 _4334_/B sky130_fd_sc_hd__nand2_1
Xoutput558 _7627_/Y vssd1 vssd1 vccd1 vccd1 sports_o[150] sky130_fd_sc_hd__buf_12
Xoutput569 _7711_/X vssd1 vssd1 vccd1 vccd1 sports_o[160] sky130_fd_sc_hd__buf_12
XANTENNA__6809__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5449__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7052_ _7051_/X _7352_/B _7097_/S vssd1 vssd1 vccd1 vccd1 _7053_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4657__B1 _4566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6003_ _5999_/Y _8919_/A _5013_/Y vssd1 vssd1 vccd1 vccd1 _6003_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8399__A1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6949__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7954_ _7954_/A vssd1 vssd1 vccd1 vccd1 _7954_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5621__A2 _5552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6905_ _6058_/A _6059_/B _8924_/B _6095_/A vssd1 vssd1 vccd1 vccd1 _6905_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_49_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7885_ _7761_/A _7883_/Y _8857_/B _7884_/Y vssd1 vssd1 vccd1 vccd1 _7885_/X sky130_fd_sc_hd__a22o_1
X_6836_ _5899_/A _6908_/B _6833_/Y _6835_/Y vssd1 vssd1 vccd1 vccd1 _6836_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8571__A1 _8252_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6767_ _6767_/A vssd1 vssd1 vccd1 vccd1 _6767_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7375__A _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8506_ _8506_/A vssd1 vssd1 vccd1 vccd1 _8506_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5718_ _5718_/A1 _4934_/A input47/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5718_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_72_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6698_ _5535_/X _6876_/C _6694_/Y _6696_/Y _6697_/Y vssd1 vssd1 vccd1 vccd1 _6699_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7126__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5137__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8437_ _8432_/X _8436_/Y _8572_/S vssd1 vssd1 vccd1 vccd1 _8438_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6334__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5649_ _5159_/B _5644_/A _5648_/Y _5125_/X vssd1 vssd1 vccd1 vccd1 _5649_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5688__A2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6885__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8368_ _8368_/A vssd1 vssd1 vccd1 vccd1 _8441_/B sky130_fd_sc_hd__inv_2
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7319_ _7319_/A vssd1 vssd1 vccd1 vccd1 _7319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8626__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8299_ _8299_/A vssd1 vssd1 vccd1 vccd1 _8299_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__7314__S _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7062__A1 _6526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7062__B2 _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6173__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8011__B1 _8011_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8562__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7365__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6901__B _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8314__A1 _8309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7117__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8314__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6325__B1 _6314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4421__B _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8617__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5300__A1 _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5851__A2 _5824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 mports_i[105] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8250__B1 _8249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5603__A2 _5640_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4951_ _4926_/X _4942_/X _6224_/S vssd1 vssd1 vccd1 vccd1 _4952_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_87_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7670_ _7767_/A _6122_/Y _7669_/X vssd1 vssd1 vccd1 vccd1 _7670_/Y sky130_fd_sc_hd__o21ai_1
X_4882_ _4974_/A vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__buf_6
XFILLER_0_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8553__B2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6621_ _6621_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6621_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6811__B _6811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6552_ _6551_/A _8151_/B _5197_/X _5196_/A vssd1 vssd1 vccd1 vccd1 _6553_/A sky130_fd_sc_hd__a22o_1
XANTENNA__8305__A1 _7825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8305__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5503_ _5845_/B _6671_/B _5502_/X _6133_/B _6386_/S vssd1 vssd1 vccd1 vccd1 _5503_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6316__B1 _4674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6483_ _6854_/A _6482_/Y _5059_/A _6549_/A vssd1 vssd1 vccd1 vccd1 _6483_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4331__B _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8222_ _4312_/B _5197_/X _8222_/B1 _5230_/B _8221_/X vssd1 vssd1 vccd1 vccd1 _8222_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_30_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5434_ _6646_/B vssd1 vssd1 vccd1 vccd1 _7105_/A sky130_fd_sc_hd__inv_2
XFILLER_0_70_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8153_ hold12/A _8150_/Y _8151_/Y _8152_/X vssd1 vssd1 vccd1 vccd1 _8153_/X sky130_fd_sc_hd__a31o_4
X_5365_ input96/X _4934_/A input33/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput366 _7782_/X vssd1 vssd1 vccd1 vccd1 mports_o[0] sky130_fd_sc_hd__buf_12
X_7104_ _7104_/A vssd1 vssd1 vccd1 vccd1 _7104_/X sky130_fd_sc_hd__buf_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput377 _7934_/X vssd1 vssd1 vccd1 vccd1 mports_o[10] sky130_fd_sc_hd__buf_12
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput388 _7947_/X vssd1 vssd1 vccd1 vccd1 mports_o[11] sky130_fd_sc_hd__buf_12
X_4316_ _4316_/A _6231_/C vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__nand2_1
Xoutput399 _7961_/X vssd1 vssd1 vccd1 vccd1 mports_o[12] sky130_fd_sc_hd__buf_12
X_8084_ _8084_/A vssd1 vssd1 vccd1 vccd1 _8084_/Y sky130_fd_sc_hd__inv_2
X_5296_ _5274_/X input95/X _4896_/A input32/X vssd1 vssd1 vccd1 vccd1 _5296_/Y sky130_fd_sc_hd__a22oi_1
X_7035_ _7034_/X _5028_/X _7097_/S vssd1 vssd1 vccd1 vccd1 _7036_/A sky130_fd_sc_hd__mux2_4
XANTENNA__7292__B2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8241__B1 _8240_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7044__B2 _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8792__A1 _8491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7937_ _7944_/A1 _4947_/B _7944_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _7937_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_78_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7868_ _7877_/A1 _5146_/A _7877_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _7868_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__8544__A1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5358__A1 _5272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7817__B _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6819_ _6906_/A _5895_/X _6818_/Y vssd1 vssd1 vccd1 vccd1 _6820_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7752__C1 _7306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7799_ _5185_/A _7803_/B1 _4566_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _7799_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6721__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4522__A _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6307__B1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5530__A1 _5510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5530__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6449__A _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7807__B1 _7814_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7035__A1 _5028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8232__B1 _8235_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5800__B _6181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6184__A _6941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7586__A2 _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6794__B1 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5349__A1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6546__B1 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6010__A2 _5923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8838__A2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6849__A1 _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4324__A2 _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5521__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5150_ _5150_/A vssd1 vssd1 vccd1 vccd1 _6544_/A sky130_fd_sc_hd__inv_2
XFILLER_0_138_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6077__A2 _6136_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7274__A1 _4793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5081_ input86/X _8310_/B input24/X _4874_/X vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5824__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8840_ _8244_/X _8806_/B _8838_/X _8839_/X vssd1 vssd1 vccd1 vccd1 _8840_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4607__A _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5037__B1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8774__A1 _8424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8774__B2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5588__A1 _5575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8771_ _7983_/Y _8711_/A _8788_/S _8770_/X vssd1 vssd1 vccd1 vccd1 _8771_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5588__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ _6875_/B _5914_/A _5982_/Y vssd1 vssd1 vccd1 vccd1 _7623_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4326__B _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6785__B1 _6779_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7722_ _7349_/Y _6965_/B _7640_/B _6278_/B vssd1 vssd1 vccd1 vccd1 _7723_/A sky130_fd_sc_hd__o22a_1
X_4934_ _4934_/A vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8526__A1 _8550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8526__B2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7653_ _6107_/A _7389_/A _6110_/A _7361_/X vssd1 vssd1 vccd1 vccd1 _7653_/X sky130_fd_sc_hd__a22o_1
X_4865_ hold2/X _4865_/B vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 _7596_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6033__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6604_ _5356_/B _6801_/A _6924_/A _5247_/X _6450_/A vssd1 vssd1 vccd1 vccd1 _6604_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4342__A hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7584_ _7584_/A _7680_/B vssd1 vssd1 vccd1 vccd1 _7584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4796_ hold29/X _8584_/B vssd1 vssd1 vccd1 vccd1 _4821_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6535_ _6535_/A vssd1 vssd1 vccd1 vccd1 _6535_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_132_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6466_ _6466_/A vssd1 vssd1 vccd1 vccd1 _6466_/X sky130_fd_sc_hd__buf_1
XANTENNA__8468__B _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7501__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7372__B _7372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8205_ _6017_/A _8209_/A2 _8204_/X vssd1 vssd1 vccd1 vccd1 _8205_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5512__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5417_ input99/X _4871_/A input37/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5417_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_113_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6397_ input79/X _8579_/C _6400_/A1 _8713_/C _6396_/X vssd1 vssd1 vccd1 vccd1 _6397_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_2_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8136_ _8151_/A _4947_/B _8150_/B _5123_/A vssd1 vssd1 vccd1 vccd1 _8136_/X sky130_fd_sc_hd__o22a_1
X_5348_ _5348_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _5348_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6068__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8462__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8067_ _8067_/A1 _7876_/X _8067_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _8067_/Y sky130_fd_sc_hd__o22ai_2
X_5279_ input30/X _4896_/A input93/X _4893_/A _5278_/X vssd1 vssd1 vccd1 vccd1 _5280_/A
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5276__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7018_ _7018_/A vssd1 vssd1 vccd1 vccd1 _7018_/X sky130_fd_sc_hd__buf_1
XANTENNA__7017__A1 _4942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8214__B1 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6208__S _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5028__B1 _5004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6776__B1 _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8969_ _8978_/CLK _8969_/D fanout732/X vssd1 vssd1 vccd1 vccd1 _8969_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6240__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6732__A _6732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7547__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7740__A2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5751__A1 _7167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5503__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6700__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__B2 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7500__A2_N _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8394__A _8394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5267__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5806__A2 _5881_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6626__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8756__A1 _7929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7559__A2 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8508__A1 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6519__B1 _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5990__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _8958_/Q vssd1 vssd1 vccd1 vccd1 _8198_/A sky130_fd_sc_hd__inv_2
XFILLER_0_126_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7731__A2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 mports_i[108] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_2
XFILLER_0_142_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput21 mports_i[118] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5742__A1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput32 mports_i[128] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4581_ _8336_/S hold21/A vssd1 vssd1 vccd1 vccd1 _8284_/A sky130_fd_sc_hd__nor2_1
Xinput43 mports_i[138] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput54 mports_i[148] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6320_ _7266_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6321_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput65 mports_i[158] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_2
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput76 mports_i[168] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_4
Xinput87 mports_i[178] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__buf_2
Xinput98 mports_i[188] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6298__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7192__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7495__A1 _6697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6251_ _6262_/A1 _8310_/B input69/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6251_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8692__B1 _8219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5202_ _5176_/Y _6128_/B _5189_/Y _5190_/Y _5201_/X vssd1 vssd1 vccd1 vccd1 _5202_/X
+ sky130_fd_sc_hd__a41o_1
X_6182_ _6182_/A1 _4935_/A input65/X _4939_/A vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5133_ _6356_/S vssd1 vssd1 vccd1 vccd1 _6261_/A sky130_fd_sc_hd__inv_2
XANTENNA__5258__B1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7798__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5064_ _6212_/A _5064_/B vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__or2_1
XFILLER_0_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8747__A1 _7886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8823_ _8203_/X _8738_/A _8206_/X _8712_/A vssd1 vssd1 vccd1 vccd1 _8823_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7973__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6222__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7648__A _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8754_ _8379_/X _8806_/B _8752_/X _8753_/Y vssd1 vssd1 vccd1 vccd1 _8754_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8953__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5966_ _5966_/A vssd1 vssd1 vccd1 vccd1 _5966_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7970__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7705_ _7756_/A _7705_/B vssd1 vssd1 vccd1 vccd1 _7705_/Y sky130_fd_sc_hd__nor2_1
X_4917_ _4917_/A vssd1 vssd1 vccd1 vccd1 _4917_/X sky130_fd_sc_hd__buf_8
XANTENNA__5981__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8685_ _8820_/A _8685_/B vssd1 vssd1 vccd1 vccd1 _8685_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5897_ _5936_/A _4932_/A _5937_/A _4929_/A _5896_/X vssd1 vssd1 vccd1 vccd1 _5924_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7636_ _7590_/A _7628_/Y _8759_/A _6059_/Y _7635_/X vssd1 vssd1 vccd1 vccd1 _7636_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_117_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4848_ _4848_/A vssd1 vssd1 vccd1 vccd1 _8934_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7722__A2 _6965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5733__A1 _5722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7567_ _5774_/A _7619_/B _7563_/X _7565_/X _7566_/Y vssd1 vssd1 vccd1 vccd1 _7567_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__5733__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4779_ _4786_/A _4788_/A _4788_/B vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__nand3_2
XANTENNA__7383__A _7383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6518_ _6854_/A _5088_/X _6544_/A _6549_/A vssd1 vssd1 vccd1 vccd1 _6518_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_132_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8198__B _8198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7498_ _7498_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7498_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6289__A2 _7720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6449_ _6449_/A vssd1 vssd1 vccd1 vccd1 _6450_/A sky130_fd_sc_hd__buf_8
XFILLER_0_101_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7238__A1 _6207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8119_ _8119_/A1 _7876_/X _8119_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _8119_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__6727__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7322__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7789__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4472__A1 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4472__B2 _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6213__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5421__B1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7961__A2 _8369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6181__B _6181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5078__A _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7713__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5724__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7477__A1 _5498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8674__B1 _8130_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7477__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5488__B1 _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7229__A1 _6212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5260__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6452__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8729__A1 _7803_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5820_ _5820_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _5820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7952__A2 _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5751_ _7167_/A _8160_/A _6456_/B _5750_/Y vssd1 vssd1 vccd1 vccd1 _5751_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5963__A1 _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5963__B2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4702_ _4751_/A _4823_/B _4751_/B vssd1 vssd1 vccd1 vccd1 _4733_/B sky130_fd_sc_hd__nand3_2
X_8470_ _8468_/Y _8469_/Y hold36/A vssd1 vssd1 vccd1 vccd1 _8471_/A sky130_fd_sc_hd__mux2_1
X_5682_ _6727_/B _5682_/B vssd1 vssd1 vccd1 vccd1 _5682_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7704__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8901__A1 _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7421_ _7083_/A _7630_/B _5301_/X _7638_/B vssd1 vssd1 vccd1 vccd1 _7421_/X sky130_fd_sc_hd__a22o_1
X_4633_ _4633_/A _4634_/A _4633_/C vssd1 vssd1 vccd1 vccd1 _4635_/A sky130_fd_sc_hd__nand3_1
XANTENNA__8299__A _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7352_ _7756_/A _7352_/B vssd1 vssd1 vccd1 vccd1 _7352_/Y sky130_fd_sc_hd__nor2_1
X_4564_ _4597_/A vssd1 vssd1 vccd1 vccd1 _5106_/A sky130_fd_sc_hd__inv_2
XFILLER_0_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6303_ _6965_/B vssd1 vssd1 vccd1 vccd1 _6303_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8665__B1 _8091_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7283_ _6367_/B _7288_/B vssd1 vssd1 vccd1 vccd1 _7283_/X sky130_fd_sc_hd__and2b_1
X_4495_ _5079_/A _6342_/A vssd1 vssd1 vccd1 vccd1 _4495_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5479__B1 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6234_ _6234_/A _6234_/B vssd1 vssd1 vccd1 vccd1 _6234_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6140__A1 _6140_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6140__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6691__A2 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6165_ _8140_/A _6161_/Y _6164_/Y vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__o21ai_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6547__A _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8026__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7142__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5116_/A vssd1 vssd1 vccd1 vccd1 _5117_/A sky130_fd_sc_hd__buf_12
XFILLER_0_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6266__B _7372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6096_ _8194_/A _6094_/X _6095_/X vssd1 vssd1 vccd1 vccd1 _6926_/B sky130_fd_sc_hd__a21o_1
X_5047_ _5047_/A vssd1 vssd1 vccd1 vccd1 _5047_/Y sky130_fd_sc_hd__inv_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5651__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7378__A _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8196__A2 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8806_ _8806_/A _8806_/B vssd1 vssd1 vccd1 vccd1 _8806_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6998_ _6998_/A vssd1 vssd1 vccd1 vccd1 _6998_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5403__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7943__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5949_ _8189_/A _5980_/B _5948_/X vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__5954__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8737_ _7821_/Y _8806_/B _8735_/X _8736_/Y vssd1 vssd1 vccd1 vccd1 _8737_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7156__A0 _7155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8668_ _8503_/A _8581_/A _8104_/Y _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8668_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5706__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7619_ _7619_/A _7619_/B vssd1 vssd1 vccd1 vccd1 _7619_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8599_ _8293_/X _8577_/X _8597_/X _8598_/Y vssd1 vssd1 vccd1 vccd1 _8599_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5182__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8105__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8120__A2 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6131__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7560__B _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6682__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput200 mports_i[74] vssd1 vssd1 vccd1 vccd1 _5402_/A sky130_fd_sc_hd__buf_2
Xinput211 mports_i[84] vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__7052__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput222 mports_i[94] vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__clkbuf_2
Xinput233 sports_i[102] vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5890__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput244 sports_i[112] vssd1 vssd1 vccd1 vccd1 _7931_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput255 sports_i[122] vssd1 vssd1 vccd1 vccd1 _8067_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__6176__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput266 sports_i[132] vssd1 vssd1 vccd1 vccd1 _8222_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput277 sports_i[1] vssd1 vssd1 vccd1 vccd1 _7790_/A2 sky130_fd_sc_hd__buf_2
Xinput288 sports_i[2] vssd1 vssd1 vccd1 vccd1 _7802_/A2 sky130_fd_sc_hd__buf_2
Xinput299 sports_i[3] vssd1 vssd1 vccd1 vccd1 _7813_/A2 sky130_fd_sc_hd__buf_2
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8187__A2 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7934__A2 _8345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5945__A1 _6007_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4424__B _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5945__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6342__D hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4440__A _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6370__A1 _6349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput707 _7058_/X vssd1 vssd1 vccd1 vccd1 sports_o[7] sky130_fd_sc_hd__buf_12
Xoutput718 _7065_/X vssd1 vssd1 vccd1 vccd1 sports_o[8] sky130_fd_sc_hd__buf_12
XANTENNA__8647__B1 _8427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput729 _7069_/X vssd1 vssd1 vccd1 vccd1 sports_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7470__B _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7870__A1 _7877_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6673__A2 _5498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7870__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5271__A _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7970_ _8404_/A _7954_/X _7969_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7970_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6921_ _6124_/X _7629_/B _8163_/A _6920_/X vssd1 vssd1 vccd1 vccd1 _6921_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4615__A _7835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6189__A1 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6852_ _6852_/A _6852_/B vssd1 vssd1 vccd1 vccd1 _6852_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7386__B1 _7385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7925__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5803_ _5803_/A vssd1 vssd1 vccd1 vccd1 _7568_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6783_ _6432_/X _6782_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6784_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8522_ _8514_/X _8349_/A _8518_/Y _8521_/Y vssd1 vssd1 vccd1 vccd1 _8522_/X sky130_fd_sc_hd__a31o_2
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5734_ _7551_/A _7299_/A _6281_/S _6758_/B vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8453_ _8453_/A _8759_/B vssd1 vssd1 vccd1 vccd1 _8453_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7645__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5665_ _6079_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _5690_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8350__A2 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7404_ _7542_/A _6578_/B _7334_/A vssd1 vssd1 vccd1 vccd1 _7404_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6041__S _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4616_ _4615_/X _4499_/B _4499_/A _7510_/A vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4350__A _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6361__A1 _6368_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5164__A2 _5208_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8384_ _4870_/X _7969_/Y _4874_/X _7942_/Y _8383_/X vssd1 vssd1 vccd1 vccd1 _8384_/X
+ sky130_fd_sc_hd__o221a_2
X_5596_ _5596_/A vssd1 vssd1 vccd1 vccd1 _5596_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6361__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7335_ _5019_/A _7753_/B _7032_/A _7349_/A _7715_/S vssd1 vssd1 vccd1 vccd1 _7335_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8638__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4547_ _4602_/A _4602_/B _4603_/B vssd1 vssd1 vccd1 vccd1 _4595_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__8102__A2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6113__A1 _6140_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7266_ _7266_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _7266_/X sky130_fd_sc_hd__and2_1
XANTENNA__6113__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4478_ _7769_/A _4478_/B vssd1 vssd1 vccd1 vccd1 _4478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8476__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7380__B _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6664__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7861__A1 _7840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6217_ _6628_/B _6217_/B vssd1 vssd1 vccd1 vccd1 _6217_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6277__A _6277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7861__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7197_ _6002_/A _7004_/X _7620_/A _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7197_/X
+ sky130_fd_sc_hd__a221o_2
X_6148_ _6183_/A1 _4953_/X input3/X _4870_/A _6147_/X vssd1 vssd1 vccd1 vccd1 _6937_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6416__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7613__A1 _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6079_ _6079_/A _6909_/A vssd1 vssd1 vccd1 vccd1 _6122_/A sky130_fd_sc_hd__nor2_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6216__S _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7916__A2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5927__A1 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7555__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7047__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5356__A _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5155__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5075__B _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6104__A1 _6104_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6104__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6655__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7080__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4969__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6634__B _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7907__A2 _7906_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7746__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8341__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5266__A _5266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8332__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5450_ _5435_/A _5089_/A _5436_/A _4868_/A _5449_/X vssd1 vssd1 vccd1 vccd1 _6671_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6343__A1 _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6343__B2 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4401_ _8160_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _4402_/A sky130_fd_sc_hd__nor2_1
Xoutput504 _6943_/X vssd1 vssd1 vccd1 vccd1 sports_o[101] sky130_fd_sc_hd__buf_12
XANTENNA__6894__A2 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8577__A _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5381_ _6634_/A _8188_/S _5400_/A _5682_/B _6481_/B vssd1 vssd1 vccd1 vccd1 _5381_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput515 _6993_/X vssd1 vssd1 vccd1 vccd1 sports_o[111] sky130_fd_sc_hd__buf_12
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput526 _7357_/Y vssd1 vssd1 vccd1 vccd1 sports_o[121] sky130_fd_sc_hd__buf_12
X_7120_ _7120_/A vssd1 vssd1 vccd1 vccd1 _7121_/A sky130_fd_sc_hd__inv_2
Xoutput537 _7464_/X vssd1 vssd1 vccd1 vccd1 sports_o[131] sky130_fd_sc_hd__buf_12
XANTENNA__8096__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4332_ _4332_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__nand2_1
Xoutput548 _7549_/X vssd1 vssd1 vccd1 vccd1 sports_o[141] sky130_fd_sc_hd__buf_12
Xoutput559 _7636_/Y vssd1 vssd1 vccd1 vccd1 sports_o[151] sky130_fd_sc_hd__buf_12
XANTENNA__6809__B _6809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7051_ _6507_/B _7026_/X _7049_/Y _7050_/X vssd1 vssd1 vccd1 vccd1 _7051_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4657__A1 _4481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6002_ _6002_/A vssd1 vssd1 vccd1 vccd1 _6002_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4657__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5854__B1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4329__B _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7953_ _7948_/Y _6024_/A _7949_/Y _6513_/A _7952_/Y vssd1 vssd1 vccd1 vccd1 _8358_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5082__A1 _5131_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6544__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5082__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4345__A hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6904_ _6094_/X _6429_/S _6903_/X vssd1 vssd1 vccd1 vccd1 _6904_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7884_ _7884_/A vssd1 vssd1 vccd1 vccd1 _7884_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8020__B2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6835_ _6835_/A _6940_/A vssd1 vssd1 vccd1 vccd1 _6835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8571__A2 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6560__A _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6582__A1 _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6766_ _6926_/A _5720_/X _6765_/Y vssd1 vssd1 vccd1 vccd1 _6767_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5717_ _5159_/B _6743_/A _5125_/X _5656_/Y _5716_/X vssd1 vssd1 vccd1 vccd1 _5717_/X
+ sky130_fd_sc_hd__a221o_1
X_8505_ _8504_/X _8457_/A _8755_/B vssd1 vssd1 vccd1 vccd1 _8506_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_33_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6697_ _6841_/A _6697_/B vssd1 vssd1 vccd1 vccd1 _6697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_127_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5137__A2 _6507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8436_ _8555_/B _8434_/X _8435_/Y vssd1 vssd1 vccd1 vccd1 _8436_/Y sky130_fd_sc_hd__o21ai_2
X_5648_ _5643_/X _6628_/B _5647_/Y vssd1 vssd1 vccd1 vccd1 _5648_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8367_ _8363_/X _8366_/X _8496_/S vssd1 vssd1 vccd1 vccd1 _8367_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5579_ _6079_/A _6695_/B vssd1 vssd1 vccd1 vccd1 _5610_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7318_ _7314_/X _4942_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7319_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8087__B2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8298_ _8564_/B _8297_/X _8349_/A vssd1 vssd1 vccd1 vccd1 _8298_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6904__B1_N _6903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7249_ _7248_/X _6263_/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7250_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7062__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6270__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8011__A1 _8011_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8011__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6022__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8562__A2 _8235_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7566__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5376__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7770__B1 _4481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4702__B _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8314__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6325__A1 _6315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6325__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7522__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8078__B2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7825__A1 _7827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7825__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5836__B1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5300__A2 _7432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7038__C1 _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 mports_i[106] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_0_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8250__A1 _8247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8250__B2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4950_ _6359_/S vssd1 vssd1 vccd1 vccd1 _6224_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4881_ _6284_/A _5762_/A vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_74_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8553__A2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6620_ _6620_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6620_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6564__A1 _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6551_ _6551_/A vssd1 vssd1 vccd1 vccd1 _6551_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8305__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5502_ _5501_/X _5451_/X _6481_/B vssd1 vssd1 vccd1 vccd1 _5502_/X sky130_fd_sc_hd__mux2_1
X_6482_ _6481_/B _5062_/D _6481_/Y vssd1 vssd1 vccd1 vccd1 _6482_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7513__B1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8221_ _7874_/A _8221_/A2 _8174_/A _4478_/B vssd1 vssd1 vccd1 vccd1 _8221_/X sky130_fd_sc_hd__a22o_1
X_5433_ _5031_/X _6630_/A _5429_/X _5432_/X vssd1 vssd1 vccd1 vccd1 _5433_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8978__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8069__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8152_ _8148_/A1 _6868_/B _8143_/B _8174_/A vssd1 vssd1 vccd1 vccd1 _8152_/X sky130_fd_sc_hd__a2bb2o_1
X_5364_ _8842_/B _5362_/Y _5363_/X vssd1 vssd1 vccd1 vccd1 _5364_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput367 _8702_/X vssd1 vssd1 vccd1 vccd1 mports_o[100] sky130_fd_sc_hd__buf_12
X_7103_ _7101_/X _6630_/A _7175_/S vssd1 vssd1 vccd1 vccd1 _7104_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7816__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput378 _8751_/X vssd1 vssd1 vccd1 vccd1 mports_o[110] sky130_fd_sc_hd__buf_12
XANTENNA__6619__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4315_ _8185_/B vssd1 vssd1 vccd1 vccd1 _6231_/C sky130_fd_sc_hd__inv_6
X_8083_ _7975_/X _8476_/A _8079_/X _8082_/X vssd1 vssd1 vccd1 vccd1 _8083_/X sky130_fd_sc_hd__a22o_4
X_5295_ _5295_/A vssd1 vssd1 vccd1 vccd1 _5295_/Y sky130_fd_sc_hd__inv_2
Xoutput389 _8786_/X vssd1 vssd1 vccd1 vccd1 mports_o[120] sky130_fd_sc_hd__buf_12
X_7034_ _5000_/X _7026_/X _7032_/X _7033_/X vssd1 vssd1 vccd1 vccd1 _7034_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7292__A2 _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8241__A1 _8239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7044__A2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6252__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8792__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7936_ _7936_/A vssd1 vssd1 vccd1 vccd1 _7936_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8529__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7867_ _7864_/Y _7761_/A _7865_/Y _8857_/B _7866_/Y vssd1 vssd1 vccd1 vccd1 _7867_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_19_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7201__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6818_ _6818_/A _6906_/A vssd1 vssd1 vccd1 vccd1 _6818_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_136_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7752__B1 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7798_ _4566_/A _5299_/B _7803_/B1 _5171_/B _7797_/X vssd1 vssd1 vccd1 vccd1 _7798_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_135_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4522__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6749_ _7551_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6749_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7504__B1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8701__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8419_ _8418_/Y _8361_/Y _8755_/B vssd1 vssd1 vccd1 vccd1 _8419_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5634__A _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5530__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7807__A1 _7814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5353__B _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7807__B2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5818__B1 _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8232__A1 _8235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8232__B2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6184__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6243__B1 _6247_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7991__B1 _7998_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6794__B2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6912__B _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7296__A _7296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5809__A _5809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6546__A1 _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6546__B2 _6526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7743__B _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6849__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7745__A2_N _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7235__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5521__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5080_ _5080_/A vssd1 vssd1 vccd1 vccd1 _8480_/B sky130_fd_sc_hd__buf_8
XFILLER_0_138_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7274__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8574__B _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5037__A1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5037__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8774__A2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8590__A _8590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5588__A2 _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5982_ _5982_/A _6875_/B vssd1 vssd1 vccd1 vccd1 _5982_/Y sky130_fd_sc_hd__nand2_1
X_8770_ _8447_/X _8770_/B vssd1 vssd1 vccd1 vccd1 _8770_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6785__A1 _5827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7982__B1 _7985_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6785__B2 _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4933_ _4933_/A vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__buf_12
X_7721_ _7719_/Y _7332_/A _7720_/Y vssd1 vssd1 vccd1 vccd1 _7721_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8526__A2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4864_ _8934_/A _8934_/B _4864_/C vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__nand3_1
XANTENNA__4623__A _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6537__A1 _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7652_ _7542_/A _6891_/A _7326_/A vssd1 vssd1 vccd1 vccd1 _7652_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 _5206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6603_ _6601_/X _6933_/A _6968_/A _6602_/X vssd1 vssd1 vccd1 vccd1 _6603_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7583_ _7177_/A _7668_/B _5905_/Y _7629_/B _7753_/B vssd1 vssd1 vccd1 vccd1 _7583_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4795_ _4607_/A _4793_/Y _4794_/Y _4792_/B vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6534_ _6534_/A _6534_/B vssd1 vssd1 vccd1 vccd1 _6534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6465_ _6464_/X _7332_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6466_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_42_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5454__A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5416_ _5385_/A _8491_/B _5386_/A _4933_/A _5415_/X vssd1 vssd1 vccd1 vccd1 _6630_/A
+ sky130_fd_sc_hd__o221a_4
X_8204_ _7852_/A _8198_/B _8189_/B vssd1 vssd1 vccd1 vccd1 _8204_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6396_ _8444_/A _6401_/A1 _8257_/C input16/X vssd1 vssd1 vccd1 vccd1 _6396_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5512__A2 _5543_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8135_ _7975_/X _8523_/A _8131_/X _8134_/X vssd1 vssd1 vccd1 vccd1 _8135_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5347_ _6233_/B _7422_/A _5334_/Y _5346_/Y vssd1 vssd1 vccd1 vccd1 _5348_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__8462__A1 _8055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8066_ _8464_/A _7954_/X _8469_/A _7826_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _8066_/X
+ sky130_fd_sc_hd__a221o_1
X_5278_ _8444_/A input34/X _8257_/C _5326_/B1 vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5276__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7017_ _7012_/X _4942_/X _7097_/S vssd1 vssd1 vccd1 vccd1 _7018_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_98_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8214__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8214__B2 _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5028__B2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8968_ _8978_/CLK _8968_/D input229/X vssd1 vssd1 vccd1 vccd1 _8968_/Q sky130_fd_sc_hd__dfrtp_4
X_7919_ _7909_/Y _7874_/A _7910_/Y _8174_/A _7918_/Y vssd1 vssd1 vccd1 vccd1 _8335_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8899_ _8899_/A _8899_/B _8899_/C vssd1 vssd1 vccd1 vccd1 _8899_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_93_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5348__B _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5751__A2 _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6700__A1 _5558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__A2 _6671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6700__B2 _5562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6179__B _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8394__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5267__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5267__B2 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4708__A _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8205__A1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8614__S _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6923__A _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7964__B1 _7971_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8508__A2 _8107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5990__A2 _6061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7754__A _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput11 mports_i[109] vssd1 vssd1 vccd1 vccd1 _4823_/B sky130_fd_sc_hd__clkbuf_8
Xinput22 mports_i[119] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4580_ hold21/A _8904_/A vssd1 vssd1 vccd1 vccd1 _8261_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_142_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 mports_i[129] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_2
Xinput44 mports_i[139] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput55 mports_i[149] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 mports_i[159] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput77 mports_i[169] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5274__A _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput88 mports_i[179] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput99 mports_i[189] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__buf_2
X_6250_ _6250_/A vssd1 vssd1 vccd1 vccd1 _6250_/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8692__A1 _8217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7495__A2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8692__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5201_ _6181_/B _7368_/B _6563_/A _6211_/B _6359_/S vssd1 vssd1 vccd1 vccd1 _5201_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6181_ _7681_/B _6181_/B vssd1 vssd1 vccd1 vccd1 _6181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_110_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5132_ input24/X _8579_/C input86/X _8713_/C _5131_/X vssd1 vssd1 vccd1 vccd1 _5132_/Y
+ sky130_fd_sc_hd__a221oi_2
XANTENNA__7247__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5258__A1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6817__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5258__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5063_ _6284_/A _5059_/A _5058_/X _5062_/X vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4337__B _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8524__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8822_ _8819_/X _8725_/X _8820_/Y _8821_/X vssd1 vssd1 vccd1 vccd1 _8822_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_149_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7955__B1 _7958_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8753_ _8381_/Y _8820_/B _8829_/S vssd1 vssd1 vccd1 vccd1 _8753_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5965_ _5965_/A vssd1 vssd1 vccd1 vccd1 _5965_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5430__A1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5430__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7704_ _6207_/A _7723_/B _7703_/X vssd1 vssd1 vccd1 vccd1 _7704_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4916_ _5193_/A vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5896_ _5962_/A1 _4935_/A input55/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__o22a_1
X_8684_ _8187_/X _8581_/A _8190_/X _8583_/A _8621_/S vssd1 vssd1 vccd1 vccd1 _8684_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7635_ _7700_/B _7628_/Y _7633_/X _7723_/B _7634_/X vssd1 vssd1 vccd1 vccd1 _7635_/X
+ sky130_fd_sc_hd__a221o_1
X_4847_ _4847_/A vssd1 vssd1 vccd1 vccd1 _8934_/A sky130_fd_sc_hd__inv_4
XFILLER_0_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8380__B1 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5883__S _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5194__B1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5733__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4778_ _4806_/B _4810_/B vssd1 vssd1 vccd1 vccd1 _4788_/B sky130_fd_sc_hd__nand2_1
X_7566_ _7590_/A _7566_/B vssd1 vssd1 vccd1 vccd1 _7566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6930__A1 _6923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7383__B _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4941__B1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6517_ _6517_/A _6517_/B vssd1 vssd1 vccd1 vccd1 _6517_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4800__B _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8132__B1 _8132_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7497_ _7497_/A _7497_/B vssd1 vssd1 vccd1 vccd1 _7497_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6448_ _6448_/A vssd1 vssd1 vccd1 vccd1 _6449_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5497__A1 _5497_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5497__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7891__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6379_ _6379_/A vssd1 vssd1 vccd1 vccd1 _6379_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5912__A _6841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8118_ _8510_/A _7954_/X _8117_/Y _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8118_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7238__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6727__B _6727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5631__B _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8049_ _8054_/A1 _5145_/A _8054_/B1 _5616_/A vssd1 vssd1 vccd1 vccd1 _8049_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_98_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8942__B hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8199__B1 _8845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4472__A2 _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8434__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6743__A _6743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7558__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7410__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5421__A1 _5465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5359__A _5359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5421__B2 _6648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5972__A2 _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7174__A1 _6788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5724__A2 _5792_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4710__B _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5094__A _5094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7477__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8674__A1 _8550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8674__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5488__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6685__B1 _5530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7229__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output425_A _8224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4999__B1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8729__A2 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6653__A _6653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7937__B1 _7944_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7468__B _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _5750_/A vssd1 vssd1 vccd1 vccd1 _5750_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5963__A2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4701_ _4701_/A _8973_/Q vssd1 vssd1 vccd1 vccd1 _4751_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5681_ _5738_/C vssd1 vssd1 vccd1 vccd1 _7542_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8901__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4632_ hold10/A _8977_/D _4837_/A _4863_/B vssd1 vssd1 vccd1 vccd1 _4633_/C sky130_fd_sc_hd__o2bb2a_1
X_7420_ _7416_/X _7418_/Y _7419_/X vssd1 vssd1 vccd1 vccd1 _7420_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_71_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4901__A _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4563_ hold12/A _4563_/B vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__nor2_2
X_7351_ _7350_/X _5042_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7351_/X sky130_fd_sc_hd__mux2_1
XANTENNA__8114__B1 _8119_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6302_ _6299_/Y _8455_/B _6300_/Y _4891_/X _6301_/Y vssd1 vssd1 vccd1 vccd1 _6965_/B
+ sky130_fd_sc_hd__o221a_2
X_7282_ _7743_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7282_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_111_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8665__A1 _8511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8665__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4494_ _4810_/B _5091_/A _4800_/B _4871_/A _4493_/X vssd1 vssd1 vccd1 vccd1 _6342_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5479__A1 _5764_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5479__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6233_ _6233_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _6233_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7873__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6140__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6828__A _6828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6164_ _6965_/A _6221_/A _8140_/A vssd1 vssd1 vccd1 vccd1 _6164_/Y sky130_fd_sc_hd__o21ai_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5139_/A _8491_/B _5140_/A _4933_/A _5114_/X vssd1 vssd1 vccd1 vccd1 _7356_/B
+ sky130_fd_sc_hd__o221a_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6095_/A _7316_/A vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__and2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5046_ _5046_/A vssd1 vssd1 vccd1 vccd1 _5046_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5651__A1 _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5651__B2 _5679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7928__B1 _7931_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8805_ _8538_/X _8788_/S _8803_/Y _8804_/Y vssd1 vssd1 vccd1 vccd1 _8805_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5403__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6997_ _6996_/X _7750_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6998_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8736_ _7837_/X _8820_/B _8829_/S vssd1 vssd1 vccd1 vccd1 _8736_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5948_ _6281_/S _5948_/B vssd1 vssd1 vccd1 vccd1 _5948_/X sky130_fd_sc_hd__or2_1
XANTENNA__5954__A2 _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8667_ _8490_/A _8577_/X _8665_/X _8666_/X vssd1 vssd1 vccd1 vccd1 _8667_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7156__A1 _5741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5879_ _5879_/A _6084_/B vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__and2_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7394__A _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5907__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5167__B1 _5130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7618_ _7378_/X _5923_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7618_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_145_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5706__A2 _5655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8598_ _8297_/X _8685_/B _8686_/B vssd1 vssd1 vccd1 vccd1 _8598_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7549_ _7545_/X _7547_/Y _7548_/X vssd1 vssd1 vccd1 vccd1 _7549_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8105__B1 _8104_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8656__A1 _8451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5642__A _5679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput201 mports_i[75] vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6457__B _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput212 mports_i[85] vssd1 vssd1 vccd1 vccd1 _5519_/A sky130_fd_sc_hd__buf_2
XANTENNA__5890__A1 _5824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput223 mports_i[95] vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__buf_2
XANTENNA__5890__B2 _5853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput234 sports_i[103] vssd1 vssd1 vccd1 vccd1 _7791_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput245 sports_i[113] vssd1 vssd1 vccd1 vccd1 _7944_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput256 sports_i[123] vssd1 vssd1 vccd1 vccd1 _8080_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput267 sports_i[133] vssd1 vssd1 vccd1 vccd1 _8235_/B1 sky130_fd_sc_hd__buf_4
Xinput278 sports_i[20] vssd1 vssd1 vccd1 vccd1 _8058_/A sky130_fd_sc_hd__buf_1
XANTENNA__7631__A2 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput289 sports_i[30] vssd1 vssd1 vccd1 vccd1 _8221_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7288__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7395__A1 _5218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5089__A _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7395__B2 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5945__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5817__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4721__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7698__A2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6370__A2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput708 _6710_/X vssd1 vssd1 vccd1 vccd1 sports_o[80] sky130_fd_sc_hd__buf_12
XFILLER_0_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8647__B2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput719 _6822_/X vssd1 vssd1 vccd1 vccd1 sports_o[90] sky130_fd_sc_hd__buf_12
XFILLER_0_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6648__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7870__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5881__A1 _5881_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5881__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7987__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6920_ _6432_/X _6919_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6920_/X sky130_fd_sc_hd__o21a_1
X_6851_ _6851_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6851_/Y sky130_fd_sc_hd__nand2_1
X_5802_ _5031_/X _5770_/X _5801_/X vssd1 vssd1 vccd1 vccd1 _5802_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6782_ _6852_/A _7171_/A vssd1 vssd1 vccd1 vccd1 _6782_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8521_ _8535_/A _8759_/B _8349_/A vssd1 vssd1 vccd1 vccd1 _8521_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5733_ _5722_/A _4868_/A _5723_/A _5089_/A _5732_/X vssd1 vssd1 vccd1 vccd1 _6758_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8452_ _8451_/Y _8433_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8453_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7689__A2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5664_ _5661_/Y _4885_/A _5662_/Y _4890_/A _5663_/Y vssd1 vssd1 vccd1 vccd1 _7532_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_60_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7403_ _6576_/B _7532_/A _7767_/A _5292_/Y _7348_/A vssd1 vssd1 vccd1 vccd1 _7403_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_143_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4615_ _7835_/A _4841_/B vssd1 vssd1 vccd1 vccd1 _4615_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8383_ _7916_/Y hold36/A _8482_/B vssd1 vssd1 vccd1 vccd1 _8383_/X sky130_fd_sc_hd__a21o_1
X_5595_ _5609_/B vssd1 vssd1 vccd1 vccd1 _5595_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4350__B _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6361__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8638__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4546_ _4546_/A _4551_/B vssd1 vssd1 vccd1 vccd1 _4602_/A sky130_fd_sc_hd__nand2_1
X_7334_ _7334_/A vssd1 vssd1 vccd1 vccd1 _7754_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6113__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7265_ _7265_/A vssd1 vssd1 vccd1 vccd1 _7265_/X sky130_fd_sc_hd__buf_1
XANTENNA__6558__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4477_ _6440_/B vssd1 vssd1 vccd1 vccd1 _7769_/A sky130_fd_sc_hd__clkinv_16
X_6216_ _6215_/Y _6184_/Y _8842_/B vssd1 vssd1 vccd1 vccd1 _6216_/X sky130_fd_sc_hd__mux2_1
X_7196_ _7196_/A vssd1 vssd1 vccd1 vccd1 _7196_/X sky130_fd_sc_hd__buf_1
XANTENNA__7861__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6147_ _6182_/A1 _5090_/A input65/X _4874_/A vssd1 vssd1 vccd1 vccd1 _6147_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6992__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6078_ _6075_/Y _4886_/A _6076_/Y _4891_/A _6077_/Y vssd1 vssd1 vccd1 vccd1 _6909_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5624__A1 _5596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5624__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7389__A _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _5026_/X _5028_/X _6224_/S vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__mux2_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8023__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8719_ _8297_/X _8820_/B _8829_/S vssd1 vssd1 vccd1 vccd1 _8719_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__7836__B _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4541__A _4557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5356__B _5356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7852__A _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8629__A1 _8379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6104__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5312__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7299__A _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5379__B1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8622__S _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8947__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6343__A2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4400_ _4454_/B vssd1 vssd1 vccd1 vccd1 _4420_/A sky130_fd_sc_hd__inv_2
XFILLER_0_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5551__B1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5380_ _5337_/A _5080_/A _5338_/A _4870_/X _5379_/X vssd1 vssd1 vccd1 vccd1 _5400_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput505 _6950_/X vssd1 vssd1 vccd1 vccd1 sports_o[102] sky130_fd_sc_hd__buf_12
XFILLER_0_112_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput516 _6998_/X vssd1 vssd1 vccd1 vccd1 sports_o[112] sky130_fd_sc_hd__buf_12
XFILLER_0_23_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput527 _7377_/X vssd1 vssd1 vccd1 vccd1 sports_o[122] sky130_fd_sc_hd__buf_12
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4331_ _4337_/A _4331_/B vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__nand2_1
XANTENNA__8096__A2 _8490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput538 _7472_/X vssd1 vssd1 vccd1 vccd1 sports_o[132] sky130_fd_sc_hd__buf_12
Xoutput549 _7557_/X vssd1 vssd1 vccd1 vccd1 sports_o[142] sky130_fd_sc_hd__buf_12
X_7050_ _6497_/B _7288_/B vssd1 vssd1 vccd1 vccd1 _7050_/X sky130_fd_sc_hd__and2b_1
X_6001_ _6001_/A _6547_/A vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5854__A1 _5827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5854__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7952_ _7958_/A1 _5145_/A _7958_/B1 _5616_/A vssd1 vssd1 vccd1 vccd1 _7952_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5082__A2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6903_ _6899_/Y _6467_/X _6900_/Y _6901_/Y _6902_/Y vssd1 vssd1 vccd1 vccd1 _6903_/X
+ sky130_fd_sc_hd__a41o_2
X_7883_ _7883_/A vssd1 vssd1 vccd1 vccd1 _7883_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4345__B hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8556__B1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6841__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6834_ _6434_/B _4824_/B _8759_/A vssd1 vssd1 vccd1 vccd1 _6940_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__8020__A2 _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6031__A1 _6031_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6031__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7656__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6765_ _6765_/A _6926_/A vssd1 vssd1 vccd1 vccd1 _6765_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8504_ _8503_/Y _8483_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8504_/X sky130_fd_sc_hd__mux2_1
X_5716_ _6261_/A _6732_/A _5708_/X _5715_/X _5136_/X vssd1 vssd1 vccd1 vccd1 _5716_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5790__B1 _5810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6696_ _6432_/X _6695_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6696_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5176__B _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6987__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8435_ _8435_/A _8441_/B vssd1 vssd1 vccd1 vccd1 _8435_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5647_ _6628_/B _5647_/B vssd1 vssd1 vccd1 vccd1 _5647_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6334__A2 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7672__A _7672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7879__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5542__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8366_ _4913_/X _8765_/B _4917_/X _7932_/Y _8365_/X vssd1 vssd1 vccd1 vccd1 _8366_/X
+ sky130_fd_sc_hd__o221a_2
X_5578_ _5575_/Y _4886_/A _5576_/Y _4891_/A _5577_/Y vssd1 vssd1 vccd1 vccd1 _6695_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7317_ _7507_/A _7372_/A vssd1 vssd1 vccd1 vccd1 _7741_/S sky130_fd_sc_hd__nand2_8
XANTENNA__5904__B _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ _5780_/A _6342_/A vssd1 vssd1 vccd1 vccd1 _4529_/Y sky130_fd_sc_hd__nor2_1
X_8297_ _8295_/Y _8364_/A _8296_/X vssd1 vssd1 vccd1 vccd1 _8297_/X sky130_fd_sc_hd__a21o_2
XANTENNA__5192__A _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6098__A1 _6141_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6098__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7248_ _6261_/B _7138_/X _7246_/X _7247_/X vssd1 vssd1 vccd1 vccd1 _7248_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout732 input229/X vssd1 vssd1 vccd1 vccd1 fanout732/X sky130_fd_sc_hd__buf_6
X_7179_ _6801_/B _7138_/X _7177_/X _7178_/X vssd1 vssd1 vccd1 vccd1 _7179_/X sky130_fd_sc_hd__o22a_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4536__A _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6270__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7847__A _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8011__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6022__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6470__B _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7770__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5367__A _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7770__B2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6325__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7522__A1 _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5533__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8078__A2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6089__A1 _6089_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6089__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7825__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5836__A1 _5871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5836__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6926__A _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6645__B _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 mports_i[107] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_87_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4880_ _5096_/A vssd1 vssd1 vccd1 vccd1 _5762_/A sky130_fd_sc_hd__inv_6
XFILLER_0_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7210__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6550_ _6550_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6550_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5772__B1 _5788_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5501_ _6679_/B _7299_/A _6017_/A _5500_/X vssd1 vssd1 vccd1 vccd1 _5501_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6481_ _6481_/A _6481_/B vssd1 vssd1 vccd1 vccd1 _6481_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7513__A1 _5659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8220_ _8217_/X _7954_/A _8219_/X _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8220_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5432_ _6202_/B _6635_/A _5136_/X vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_30_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8069__A2 _8068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5363_ _8194_/A _5363_/B vssd1 vssd1 vccd1 vccd1 _5363_/X sky130_fd_sc_hd__or2_1
X_8151_ _8151_/A _8151_/B vssd1 vssd1 vccd1 vccd1 _8151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7277__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7102_ _7295_/S vssd1 vssd1 vccd1 vccd1 _7175_/S sky130_fd_sc_hd__buf_6
XFILLER_0_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput368 _8705_/X vssd1 vssd1 vccd1 vccd1 mports_o[101] sky130_fd_sc_hd__buf_12
X_4314_ hold37/X vssd1 vssd1 vccd1 vccd1 _8185_/B sky130_fd_sc_hd__buf_8
X_5294_ _5294_/A vssd1 vssd1 vccd1 vccd1 _5294_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7816__A2 _7807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8082_ _7777_/A _8081_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _8082_/X sky130_fd_sc_hd__o21ba_1
Xoutput379 _8754_/X vssd1 vssd1 vccd1 vccd1 mports_o[111] sky130_fd_sc_hd__buf_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7033_ _5019_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7033_/X sky130_fd_sc_hd__a21o_1
XANTENNA__8947__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8777__B1 _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6252__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7935_ _7935_/A vssd1 vssd1 vccd1 vccd1 _7935_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8529__B1 _8148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8262__S _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7866_ _7877_/A1 _4947_/B _7877_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _7866_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__6004__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6817_ _6817_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6817_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6290__B _6375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7752__A1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7797_ _6965_/A _7802_/A2 _8163_/A _4326_/B vssd1 vssd1 vccd1 vccd1 _7797_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6555__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5187__A _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6748_ _6506_/A _5765_/X _6449_/A vssd1 vssd1 vccd1 vccd1 _6748_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8498__A _8498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6307__A2 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6679_ _6841_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _6679_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7504__A1 _5552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8701__B1 _8240_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8418_ _8418_/A vssd1 vssd1 vccd1 vccd1 _8418_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5634__B _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8349_ _8349_/A _8349_/B vssd1 vssd1 vccd1 vccd1 _8349_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7807__A2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5818__A1 _5011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8437__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8232__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6243__A1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6243__B2 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7991__A1 _7998_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7577__A _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6546__A2 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5097__A _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output455_A _8522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8347__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6482__A1 _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6375__B _6375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4493__B1 _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8223__A2 _8222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5037__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5981_ _8189_/A _6042_/B _5980_/X vssd1 vssd1 vccd1 vccd1 _5982_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7982__A1 _7985_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6785__A2 _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7982__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7720_ _7756_/A _7720_/B vssd1 vssd1 vccd1 vccd1 _7720_/Y sky130_fd_sc_hd__nor2_1
X_4932_ _4932_/A vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__buf_8
XANTENNA__4904__A _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7651_ _7651_/A _7651_/B vssd1 vssd1 vccd1 vccd1 _7651_/X sky130_fd_sc_hd__or2_1
X_4863_ _4866_/A _4863_/B _4863_/C vssd1 vssd1 vccd1 vccd1 _4864_/C sky130_fd_sc_hd__and3_1
XFILLER_0_7_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6602_ _7422_/A _6913_/B _5264_/Y _6912_/B vssd1 vssd1 vccd1 vccd1 _6602_/X sky130_fd_sc_hd__a22o_1
XANTENNA_14 _7454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8810__S _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7582_ _6804_/Y _7619_/B _7578_/X _7580_/Y _7581_/Y vssd1 vssd1 vccd1 vccd1 _7582_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4794_ hold29/X _5192_/A vssd1 vssd1 vccd1 vccd1 _4794_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_103_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6533_ _5159_/A _6908_/B _6569_/B _6512_/X vssd1 vssd1 vccd1 vccd1 _6534_/B sky130_fd_sc_hd__a22oi_1
XFILLER_0_82_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5735__A _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6464_ _6463_/X _4992_/X _7000_/S vssd1 vssd1 vccd1 vccd1 _6464_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8203_ _8210_/A1 _6456_/B _8210_/B1 _6495_/B _8202_/X vssd1 vssd1 vccd1 vccd1 _8203_/X
+ sky130_fd_sc_hd__o221a_2
X_5415_ input97/X _8368_/A input35/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5415_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6395_ _6395_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _7753_/A sky130_fd_sc_hd__and2_1
XFILLER_0_3_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8134_ _7777_/A _8133_/Y _7792_/A vssd1 vssd1 vccd1 vccd1 _8134_/X sky130_fd_sc_hd__o21ba_1
X_5346_ _6616_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8765__B _8765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8462__A2 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6566__A _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8065_ _8058_/Y _7769_/A _8059_/Y _6500_/A _8064_/Y vssd1 vssd1 vccd1 vccd1 _8469_/A
+ sky130_fd_sc_hd__a221oi_4
X_5277_ _5272_/Y _4885_/A _5273_/Y _4890_/A _5276_/Y vssd1 vssd1 vccd1 vccd1 _5333_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5276__A2 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7016_ _7295_/S vssd1 vssd1 vccd1 vccd1 _7097_/S sky130_fd_sc_hd__buf_8
XFILLER_0_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5028__A2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8967_ _8967_/CLK _8967_/D input229/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__7973__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6776__A2 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7918_ _7918_/A1 _7876_/A _7918_/B1 _7835_/A vssd1 vssd1 vccd1 vccd1 _7918_/Y sky130_fd_sc_hd__o22ai_2
X_8898_ _8898_/A _8898_/B vssd1 vssd1 vccd1 vccd1 _8974_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7849_ _7847_/Y _7848_/Y _8185_/B vssd1 vssd1 vccd1 vccd1 _7849_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_136_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5751__A3 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5645__A _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7489__B1 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6700__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5267__A2 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4475__B1 _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4708__B hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8205__A2 _8209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7964__A1 _7971_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7964__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6519__A2 _5105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7716__A1 _6263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 mports_i[10] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput23 mports_i[11] vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__clkbuf_4
Xinput34 mports_i[12] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_2
Xinput45 mports_i[13] vssd1 vssd1 vccd1 vccd1 _5272_/A sky130_fd_sc_hd__buf_2
XFILLER_0_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput56 mports_i[14] vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput67 mports_i[15] vssd1 vssd1 vccd1 vccd1 _5337_/A sky130_fd_sc_hd__clkbuf_4
Xinput78 mports_i[16] vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput89 mports_i[17] vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8692__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5200_ _5200_/A vssd1 vssd1 vccd1 vccd1 _6563_/A sky130_fd_sc_hd__inv_2
XFILLER_0_110_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6180_ _6180_/A vssd1 vssd1 vccd1 vccd1 _7681_/B sky130_fd_sc_hd__inv_2
XFILLER_0_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5131_ _8444_/A _5131_/A2 _8257_/C _5131_/B2 vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5258__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5062_ _8709_/A _8189_/A _8189_/B _5062_/D vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__or4_4
XANTENNA__7652__B1 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4618__B _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8821_ _8821_/A _8829_/S vssd1 vssd1 vccd1 vccd1 _8821_/X sky130_fd_sc_hd__and2_1
XANTENNA__7404__B1 _7334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7955__A1 _7958_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7955__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8752_ _8384_/X _8711_/X _8386_/X _8803_/B _8820_/B vssd1 vssd1 vccd1 vccd1 _8752_/X
+ sky130_fd_sc_hd__a221o_1
X_5964_ _6839_/B vssd1 vssd1 vccd1 vccd1 _7611_/A sky130_fd_sc_hd__inv_2
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5430__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7703_ _6234_/A _7753_/B _6944_/Y _7349_/A _7749_/S vssd1 vssd1 vccd1 vccd1 _7703_/X
+ sky130_fd_sc_hd__a221o_1
X_4915_ _8271_/B vssd1 vssd1 vccd1 vccd1 _8716_/B sky130_fd_sc_hd__buf_8
X_8683_ _8556_/X _8686_/B _8681_/X _8682_/Y vssd1 vssd1 vccd1 vccd1 _8683_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5895_ _5853_/X _7316_/A _8924_/B _5885_/X vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7634_ _6867_/A _7681_/A _7361_/X _6882_/A vssd1 vssd1 vccd1 vccd1 _7634_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4846_ _4848_/A _4847_/A hold4/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8380__A1 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8380__B2 _7945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5194__A1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6391__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5194__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7565_ _7700_/B _7566_/B _6771_/A _7754_/A vssd1 vssd1 vccd1 vccd1 _7565_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4777_ _4777_/A _4777_/B vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7156__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5465__A _5465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6930__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4941__A1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6516_ _6516_/A _6899_/B vssd1 vssd1 vccd1 vccd1 _6517_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8668__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4941__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8132__A1 _8132_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7496_ _5581_/Y _7668_/B _7495_/X _7266_/B vssd1 vssd1 vccd1 vccd1 _7497_/A sky130_fd_sc_hd__a22o_1
XANTENNA__8132__B2 _7835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6447_ _6517_/B vssd1 vssd1 vccd1 vccd1 _6958_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6143__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8683__A2 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5497__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7891__B1 _7890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6378_ _6388_/A1 _8480_/B input15/X _4870_/X _6377_/X vssd1 vssd1 vccd1 vccd1 _6379_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5912__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8117_ _8110_/Y _7769_/X _8111_/Y _6500_/X _8116_/Y vssd1 vssd1 vccd1 vccd1 _8117_/Y
+ sky130_fd_sc_hd__a221oi_4
X_5329_ _5329_/A _8842_/B vssd1 vssd1 vccd1 vccd1 _5329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8048_ _8045_/Y _7013_/A _8046_/Y _5117_/A _8047_/Y vssd1 vssd1 vccd1 vccd1 _8451_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__8199__A1 _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7946__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6743__B _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5421__A2 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5359__B _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5972__A3 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7174__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6921__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5094__B _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6134__B1 _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8686__A _8821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7590__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5488__A2 _6653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6685__B2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4719__A _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6437__A1 _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7634__B1 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4999__A1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4999__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output418_A _8122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7937__A1 _7944_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7937__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8360__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _8239_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5680_ _5125_/X _5657_/X _5678_/X _6402_/A _5679_/X vssd1 vssd1 vccd1 vccd1 _5680_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8362__A1 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4631_ _4844_/B vssd1 vssd1 vccd1 vccd1 _4634_/A sky130_fd_sc_hd__inv_2
XANTENNA__8901__A3 _4662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7350_ _6499_/A _7640_/B _7349_/Y _6497_/B vssd1 vssd1 vccd1 vccd1 _7350_/X sky130_fd_sc_hd__o22a_1
X_4562_ _7876_/A vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__inv_8
XFILLER_0_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8114__A1 _8119_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8114__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6301_ _8713_/C _6309_/A1 _8579_/C input71/X vssd1 vssd1 vccd1 vccd1 _6301_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_25_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8665__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7281_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7281_/X sky130_fd_sc_hd__buf_1
X_4493_ _4823_/B _5089_/A _4818_/B _4953_/A vssd1 vssd1 vccd1 vccd1 _4493_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_111_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5479__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6232_ _6304_/A _6944_/A _6231_/X vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__7873__B1 _7871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6828__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6163_ input65/X _8579_/C _6182_/A1 _4893_/A _6162_/X vssd1 vssd1 vccd1 vccd1 _6221_/A
+ sky130_fd_sc_hd__a221oi_4
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7005__A _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5114_ input87/X _8368_/A input25/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__o22a_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6047_/A _5111_/A _6048_/A _4931_/A _6093_/X vssd1 vssd1 vccd1 vccd1 _6094_/X
+ sky130_fd_sc_hd__o221a_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5100__A1 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5045_ _5046_/A _4953_/X _5047_/A _4870_/A _5044_/X vssd1 vssd1 vccd1 vccd1 _5059_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5100__B2 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5651__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6563__B _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7928__A1 _7931_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7928__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8804_ _8117_/Y _8711_/X _8788_/S vssd1 vssd1 vccd1 vccd1 _8804_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6996_ _6995_/Y _6385_/A _7000_/S vssd1 vssd1 vccd1 vccd1 _6996_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5403__A2 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8735_ _7825_/X _8711_/X _7832_/Y _8803_/B _8820_/B vssd1 vssd1 vccd1 vccd1 _8735_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5947_ _6002_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _5980_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8666_ _8698_/B _8516_/A _8590_/X vssd1 vssd1 vccd1 vccd1 _8666_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5878_ _5999_/B _7177_/A _5877_/X _5174_/A vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5167__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5907__B _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7617_ _7590_/A _7609_/Y _7610_/Y _7616_/X vssd1 vssd1 vccd1 vccd1 _7617_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__6364__B1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5167__B2 _5222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4829_ _4828_/Y _4619_/Y hold7/X vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8597_ _7800_/X _8583_/X _8303_/X _8581_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8597_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6903__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7548_ _7701_/A _7547_/A _7359_/A _6746_/Y vssd1 vssd1 vccd1 vccd1 _7548_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__8105__A1 _8503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8105__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7479_ _7479_/A vssd1 vssd1 vccd1 vccd1 _7479_/X sky130_fd_sc_hd__buf_1
XFILLER_0_114_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5923__A _5923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5642__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput202 mports_i[76] vssd1 vssd1 vccd1 vccd1 _5435_/A sky130_fd_sc_hd__buf_2
Xinput213 mports_i[86] vssd1 vssd1 vccd1 vccd1 _5723_/A sky130_fd_sc_hd__buf_2
XANTENNA__7616__B1 _7614_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput224 mports_i[96] vssd1 vssd1 vccd1 vccd1 _6021_/A sky130_fd_sc_hd__buf_2
XANTENNA__5890__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput235 sports_i[104] vssd1 vssd1 vccd1 vccd1 _7803_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput246 sports_i[114] vssd1 vssd1 vccd1 vccd1 _7958_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput257 sports_i[124] vssd1 vssd1 vccd1 vccd1 _8093_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7092__A1 _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput268 sports_i[134] vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__clkbuf_2
Xinput279 sports_i[21] vssd1 vssd1 vccd1 vccd1 _8071_/A sky130_fd_sc_hd__buf_1
XANTENNA__7631__A3 _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7919__B2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8041__B1 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8592__A1 _7763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7395__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8344__A1 _7932_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5817__B _5829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6355__B1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput709 _6716_/X vssd1 vssd1 vccd1 vccd1 sports_o[81] sky130_fd_sc_hd__buf_12
XFILLER_0_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5833__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6648__B _6648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5330__A1 _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5881__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__8280__B1 _7800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6850_ _6843_/Y _6450_/X _6846_/Y _6848_/Y _6849_/X vssd1 vssd1 vccd1 vccd1 _6850_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_77_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7386__A2 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5801_ _6170_/A _5786_/X _5136_/X _5798_/Y _5800_/Y vssd1 vssd1 vccd1 vccd1 _5801_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6781_ _5832_/B _6780_/A _6780_/Y _6724_/A vssd1 vssd1 vccd1 vccd1 _6784_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8520_ _8519_/Y _8490_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8535_/A sky130_fd_sc_hd__mux2_1
X_5732_ _5792_/A1 _4871_/A input49/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5732_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4912__A _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8451_ _8451_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8451_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5663_ _5274_/X _5697_/A1 _5275_/X input46/X vssd1 vssd1 vccd1 vccd1 _5663_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6346__B1 _6342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7402_ _6587_/Y _7619_/B _7397_/X _7400_/Y _7401_/Y vssd1 vssd1 vccd1 vccd1 _7402_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4614_ _7311_/A vssd1 vssd1 vccd1 vccd1 _7835_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8382_ _8564_/B _8381_/Y _8349_/A vssd1 vssd1 vccd1 vccd1 _8382_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5594_ _5591_/Y _4886_/A _5592_/Y _4891_/A _5593_/Y vssd1 vssd1 vccd1 vccd1 _5609_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_142_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7333_ _7328_/Y _7332_/A _7332_/Y vssd1 vssd1 vccd1 vccd1 _7333_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8638__A2 _8772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4545_ _4554_/A _8150_/A vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6839__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7846__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7264_ _7263_/Y _7729_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7265_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4476_ _4476_/A _7852_/A _4476_/C vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__and3_1
XANTENNA__6558__B _6558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6215_ _7705_/B _6626_/B vssd1 vssd1 vccd1 vccd1 _6215_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5321__A1 _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7195_ _7194_/X _5924_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7196_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6146_ _6135_/X _6402_/A _6145_/X vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__a21o_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _5274_/X _6136_/A1 _5275_/X input62/X vssd1 vssd1 vccd1 vccd1 _6077_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__5085__B1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5624__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6821__A1 _5885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5028_ _5003_/A _4933_/X _5004_/A _4930_/X _5027_/X vssd1 vssd1 vccd1 vccd1 _5028_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8023__B1 _8423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout733_A input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7377__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5388__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6979_ _6979_/A vssd1 vssd1 vccd1 vccd1 _6979_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5918__A _5918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8718_ _7771_/X _8711_/X _8303_/X _8803_/B _8820_/B vssd1 vssd1 vccd1 vccd1 _8718_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8326__A1 _7867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8649_ _8648_/X _8433_/A _8690_/S vssd1 vssd1 vccd1 vccd1 _8650_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4541__B _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6888__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7852__B _7858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8629__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6749__A _7551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5372__B _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8801__A2 _8107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7299__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8565__A1 _8226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5379__A1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5379__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8317__A1 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6328__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6879__A1 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5000__B1 _5004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7540__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5551__A1 _5635_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6659__A _7459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5551__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput506 _6954_/X vssd1 vssd1 vccd1 vccd1 sports_o[103] sky130_fd_sc_hd__buf_12
Xoutput517 _7002_/X vssd1 vssd1 vccd1 vccd1 sports_o[113] sky130_fd_sc_hd__buf_12
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4330_ _7847_/A _4611_/B vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__nand2_1
Xoutput528 _7392_/Y vssd1 vssd1 vccd1 vccd1 sports_o[123] sky130_fd_sc_hd__buf_12
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput539 _7479_/X vssd1 vssd1 vccd1 vccd1 sports_o[133] sky130_fd_sc_hd__buf_12
XFILLER_0_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5282__B _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6000_ _5997_/Y _5999_/Y _5185_/A vssd1 vssd1 vccd1 vccd1 _6000_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5854__A2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7056__A1 _5105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5502__S _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5067__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6803__A1 _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7951_ _7948_/Y _7013_/A _7949_/Y _5117_/A _7950_/Y vssd1 vssd1 vccd1 vccd1 _8369_/A
+ sky130_fd_sc_hd__a221oi_4
X_6902_ _6112_/B _6801_/A _6528_/A _6110_/A _6450_/A vssd1 vssd1 vccd1 vccd1 _6902_/Y
+ sky130_fd_sc_hd__o221ai_4
X_7882_ _7882_/A vssd1 vssd1 vccd1 vccd1 _7882_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8556__A1 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8556__B2 _8200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6833_ _6941_/A _6835_/A _6832_/Y vssd1 vssd1 vccd1 vccd1 _6833_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6841__B _6841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6031__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5738__A _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6764_ _6764_/A vssd1 vssd1 vccd1 vccd1 _6765_/A sky130_fd_sc_hd__inv_2
XANTENNA__8308__A1 _7786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8503_ _8503_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8503_/Y sky130_fd_sc_hd__nand2_1
X_5715_ _5715_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5715_/X sky130_fd_sc_hd__and2_1
XANTENNA__5790__A1 _5809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6695_ _6852_/A _6695_/B vssd1 vssd1 vccd1 vccd1 _6695_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5790__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8434_ _8433_/Y _8400_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8434_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5646_ _8842_/B _7507_/B _5645_/Y vssd1 vssd1 vccd1 vccd1 _5647_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7672__B _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8365_ _7906_/Y _8336_/S _8364_/Y vssd1 vssd1 vccd1 vccd1 _8365_/X sky130_fd_sc_hd__a21o_1
X_5577_ _5274_/X _5587_/A1 _5275_/X input41/X vssd1 vssd1 vccd1 vccd1 _5577_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__6569__A _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7164__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7316_ _7316_/A hold20/A vssd1 vssd1 vccd1 vccd1 _7372_/A sky130_fd_sc_hd__nand2_8
XANTENNA__7819__B1 _8845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4528_ _4528_/A _4528_/B vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8296_ _8584_/A _7803_/Y _7837_/X _8261_/A vssd1 vssd1 vccd1 vccd1 _8296_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6098__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7295__A1 _7756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7247_ _6252_/X _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7247_/X sky130_fd_sc_hd__a21o_1
X_4459_ _4459_/A vssd1 vssd1 vccd1 vccd1 _4460_/B sky130_fd_sc_hd__inv_2
Xfanout733 input229/X vssd1 vssd1 vccd1 vccd1 fanout733/X sky130_fd_sc_hd__buf_6
X_7178_ _5879_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7178_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7047__A1 _7345_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8244__B1 _8252_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6129_ _5108_/A _7673_/B _5136_/A _6112_/X _6128_/Y vssd1 vssd1 vccd1 vccd1 _6129_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8795__A1 _8476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6270__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7847__B _7858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6751__B _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6022__A2 _6089_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7770__A2 _4318_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5367__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7522__A2 _5655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5533__A1 _5500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5533__B2 _6697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6730__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6089__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5836__A2 _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7038__B2 _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8235__B1 _8235_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7249__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7210__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6153__S _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5221__B1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5772__A1 _5788_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5772__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7773__A _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5500_ _5505_/A _4953_/X _5506_/A _4870_/A _5499_/X vssd1 vssd1 vccd1 vccd1 _5500_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4980__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6480_ _5050_/Y _6475_/A _5051_/X _6694_/B vssd1 vssd1 vccd1 vccd1 _6480_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7513__A2 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5431_ _5385_/A _8271_/A _5386_/A _5191_/X _5430_/X vssd1 vssd1 vccd1 vccd1 _6635_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6389__A _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5524__A1 _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8150_ _8150_/A _8150_/B vssd1 vssd1 vccd1 vccd1 _8150_/Y sky130_fd_sc_hd__nand2_1
X_5362_ _5362_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5362_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7277__A1 _6349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7101_ _6635_/A _7026_/X _7099_/X _7100_/X vssd1 vssd1 vccd1 vccd1 _7101_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4313_ _8185_/A _4313_/B vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__nand2_1
Xoutput369 _8720_/X vssd1 vssd1 vccd1 vccd1 mports_o[102] sky130_fd_sc_hd__buf_12
X_8081_ _8071_/Y _7874_/X _8072_/Y _7875_/X _8080_/Y vssd1 vssd1 vccd1 vccd1 _8081_/Y
+ sky130_fd_sc_hd__a221oi_4
X_5293_ _5280_/A _6470_/B _5292_/Y vssd1 vssd1 vccd1 vccd1 _6591_/B sky130_fd_sc_hd__a21bo_1
X_7032_ _7032_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7032_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8226__B1 _8235_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5232__S _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8777__A1 _8009_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7013__A _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6252__A2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7948__A _7948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7934_ _7760_/X _8345_/A _7930_/X _7933_/X vssd1 vssd1 vccd1 vccd1 _7934_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6852__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8529__A1 _8145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5460__B1 _5402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8529__B2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7865_ _7865_/A vssd1 vssd1 vccd1 vccd1 _7865_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7201__A1 _6028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6816_ _6828_/A vssd1 vssd1 vccd1 vccd1 _6817_/A sky130_fd_sc_hd__inv_2
XANTENNA__7201__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7796_ _4566_/A _6059_/B _7803_/B1 _5359_/B _7795_/X vssd1 vssd1 vccd1 vccd1 _7796_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6747_ _7544_/A _7536_/B _7707_/B _5765_/X vssd1 vssd1 vccd1 vccd1 _6747_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5763__A1 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5763__B2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7683__A _7683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6678_ _6432_/X _6677_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6678_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__8701__A1 _8239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7504__A2 _7686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8701__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8417_ _8416_/Y _8394_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8418_/A sky130_fd_sc_hd__mux2_1
X_5629_ _8150_/A _7526_/B _7509_/A vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6299__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5407__S _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8348_ _8348_/A vssd1 vssd1 vccd1 vccd1 _8349_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8279_ _8279_/A vssd1 vssd1 vccd1 vccd1 _8279_/X sky130_fd_sc_hd__buf_1
XANTENNA__5931__A _5931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5279__B1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8217__B1 _8222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8768__A1 _7972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6243__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7440__B2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__B1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6481__B _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8940__A1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6951__B1 _7242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6703__B1 _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6002__A _6002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7259__A1 _7725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6937__A _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6482__A2 _5062_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8208__B1 _7707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4493__A1 _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4493__B2 _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5980_ _6017_/A _5980_/B vssd1 vssd1 vccd1 vccd1 _5980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5442__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7982__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4931_ _4931_/A vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__buf_8
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5288__A _5288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7650_ _7767_/A _7650_/B vssd1 vssd1 vccd1 vccd1 _7651_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7195__A0 _7194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4862_ _4848_/A _4847_/A hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7734__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6601_ _7083_/A _6475_/X _5285_/X _6851_/B vssd1 vssd1 vccd1 vccd1 _6601_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7581_ _7590_/A _7581_/B vssd1 vssd1 vccd1 vccd1 _7581_/Y sky130_fd_sc_hd__nor2_1
X_4793_ _4793_/A vssd1 vssd1 vccd1 vccd1 _4793_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6942__B1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6532_ _7356_/B _6059_/B _8924_/B _5159_/A vssd1 vssd1 vccd1 vccd1 _6569_/B sky130_fd_sc_hd__a22o_1
XANTENNA__4920__A _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6463_ _6455_/Y _6876_/C _6459_/X _6899_/B _6462_/Y vssd1 vssd1 vccd1 vccd1 _6463_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8695__B1 _8590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8202_ _8140_/A _8209_/A2 _8201_/X vssd1 vssd1 vccd1 vccd1 _8202_/X sky130_fd_sc_hd__a21o_1
X_5414_ _5031_/X _5367_/A _5412_/Y _5413_/X vssd1 vssd1 vccd1 vccd1 _5414_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6394_ _6401_/A1 _8480_/B input16/X _4870_/X _6393_/X vssd1 vssd1 vccd1 vccd1 _6395_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8133_ _8123_/Y _7874_/A _8124_/Y _8174_/A _8132_/Y vssd1 vssd1 vccd1 vccd1 _8133_/Y
+ sky130_fd_sc_hd__a221oi_4
X_5345_ _5345_/A vssd1 vssd1 vccd1 vccd1 _6616_/A sky130_fd_sc_hd__inv_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6847__A _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8064_ _8067_/A1 _5780_/A _8067_/B1 _5079_/A vssd1 vssd1 vccd1 vccd1 _8064_/Y sky130_fd_sc_hd__o22ai_4
X_5276_ _5274_/X input94/X _5275_/X input31/X vssd1 vssd1 vccd1 vccd1 _5276_/Y sky130_fd_sc_hd__a22oi_2
XANTENNA__6566__B _6566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7015_ _7015_/A vssd1 vssd1 vccd1 vccd1 _7295_/S sky130_fd_sc_hd__buf_6
XANTENNA__7670__A1 _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8966_ _8967_/CLK _8966_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__5433__B1 _5429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7973__A2 _7972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7917_ _8352_/A _7768_/X _7916_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7917_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5984__A1 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5984__B2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8897_ _4824_/B _8896_/Y _4810_/A vssd1 vssd1 vccd1 vccd1 _8898_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5198__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7186__A0 _7185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7848_ _8160_/A _7859_/B vssd1 vssd1 vccd1 vccd1 _7848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5736__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7779_ _7778_/Y _8174_/A _4331_/B _7779_/B1 _7874_/A vssd1 vssd1 vccd1 vccd1 _7779_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5926__A _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5645__B _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7489__A1 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5661__A _5661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7661__B2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8610__B1 _7871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7964__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5975__A1 _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output398_A _8818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 mports_i[110] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 mports_i[120] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput35 mports_i[130] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput46 mports_i[140] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
Xinput57 mports_i[150] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_1
Xinput68 mports_i[160] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_2
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput79 mports_i[170] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5130_ _5130_/A vssd1 vssd1 vccd1 vccd1 _8257_/C sky130_fd_sc_hd__buf_8
XFILLER_0_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6455__A2 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7652__A1 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5061_ _8189_/A _7037_/B _5060_/X vssd1 vssd1 vccd1 vccd1 _5062_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__4466__A1 _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7404__A1 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8601__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8820_ _8820_/A _8820_/B vssd1 vssd1 vccd1 vccd1 _8820_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4915__A _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7955__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5963_ _5936_/A _5191_/X _5937_/A _8271_/A _5962_/X vssd1 vssd1 vccd1 vccd1 _6847_/A
+ sky130_fd_sc_hd__o221a_4
X_8751_ _8372_/X _8806_/B _8749_/X _8750_/X vssd1 vssd1 vccd1 vccd1 _8751_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4634__B _8967_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4914_ _5192_/A vssd1 vssd1 vccd1 vccd1 _8271_/B sky130_fd_sc_hd__buf_8
X_7702_ _6218_/Y _7359_/A _7698_/X _7700_/Y _7701_/Y vssd1 vssd1 vccd1 vccd1 _7702_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8682_ _8547_/A _8685_/B _8686_/B vssd1 vssd1 vccd1 vccd1 _8682_/Y sky130_fd_sc_hd__a21oi_1
X_5894_ _5159_/B _5853_/X _5883_/X _5136_/X _5893_/X vssd1 vssd1 vccd1 vccd1 _5894_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5718__A1 _5718_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4845_ _4845_/A _4845_/B _4845_/C vssd1 vssd1 vccd1 vccd1 _4847_/A sky130_fd_sc_hd__nand3_4
X_7633_ _6029_/B _7660_/B _7629_/Y _7631_/X _7632_/Y vssd1 vssd1 vccd1 vccd1 _7633_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__5718__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8380__A2 _7972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4650__A _8958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7564_ _7510_/B _5770_/X _7398_/A vssd1 vssd1 vccd1 vccd1 _7566_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__6391__A1 _6400_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5194__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4776_ _4776_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _4777_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6391__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6515_ _7055_/A _8755_/C _8163_/A _6514_/Y vssd1 vssd1 vccd1 vccd1 _6516_/A sky130_fd_sc_hd__a31o_1
XANTENNA__8668__B1 _8104_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4941__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7495_ _6697_/B _5682_/B _8709_/A vssd1 vssd1 vccd1 vccd1 _7495_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_130_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8132__A2 _7876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6446_ _6946_/S vssd1 vssd1 vccd1 vccd1 _6517_/B sky130_fd_sc_hd__inv_2
XANTENNA__6143__A1 _6094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6143__B2 _6908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7680__B _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7891__A1 _7888_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6377_ _6387_/A1 _8310_/B input77/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6377_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7891__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8116_ _8119_/A1 _5780_/X _8119_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _8116_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5328_ _5328_/A _5361_/A vssd1 vssd1 vccd1 vccd1 _5363_/B sky130_fd_sc_hd__nand2_1
X_8047_ _8054_/A1 _4947_/B _8054_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _8047_/Y sky130_fd_sc_hd__o22ai_2
X_5259_ input34/X _4953_/X _5326_/B1 _5089_/X _5258_/X vssd1 vssd1 vccd1 vccd1 _7413_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__8199__A2 _8209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7946__A2 _7945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5957__A1 _5965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8949_ _8979_/CLK _8949_/D fanout732/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5957__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7159__B1 _7158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4560__A _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6382__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6921__A3 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8659__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6134__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8686__B _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6487__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7095__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6437__A2 _4960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4999__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7937__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8152__A1_N _8148_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8362__A2 _7901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5566__A _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4630_ _4760_/A _4837_/A _8893_/A vssd1 vssd1 vccd1 vccd1 _4844_/B sky130_fd_sc_hd__and3_1
XANTENNA__4470__A _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6373__A1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4561_ _8181_/A hold12/A vssd1 vssd1 vccd1 vccd1 _7876_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_142_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8114__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6300_ input8/X vssd1 vssd1 vccd1 vccd1 _6300_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7280_ _7279_/X _6358_/X _7295_/S vssd1 vssd1 vccd1 vccd1 _7281_/A sky130_fd_sc_hd__mux2_2
X_4492_ _8481_/S _4727_/C vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6231_ _7767_/A _7829_/A _6231_/C _6944_/A vssd1 vssd1 vccd1 vccd1 _6231_/X sky130_fd_sc_hd__or4_1
XANTENNA__7873__A1 _7869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7873__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6162_ _8444_/A _6183_/A1 _8257_/C input3/X vssd1 vssd1 vccd1 vccd1 _6162_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_21_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5113_ _5070_/A _8491_/B _5071_/A _4933_/A _5112_/X vssd1 vssd1 vccd1 vccd1 _7345_/B
+ sky130_fd_sc_hd__o221a_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7625__B2 _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6093_ _6104_/A1 _4934_/A input61/X _4938_/A vssd1 vssd1 vccd1 vccd1 _6093_/X sky130_fd_sc_hd__o22a_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ input84/X _5090_/A input21/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__o22a_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7928__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8803_ _8803_/A _8803_/B vssd1 vssd1 vccd1 vccd1 _8803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8050__B2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5939__B2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6995_ _6379_/Y _6899_/B _6994_/X vssd1 vssd1 vccd1 vccd1 _6995_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6600__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8734_ _7807_/X _8725_/X _8731_/Y _8733_/X vssd1 vssd1 vccd1 vccd1 _8734_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6860__A _6868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5946_ _5931_/A _4868_/A _5932_/A _4870_/A _5945_/X vssd1 vssd1 vccd1 vccd1 _6002_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_137_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8665_ _8511_/A _8581_/X _8091_/Y _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8665_/X
+ sky130_fd_sc_hd__a221o_1
X_5877_ _7592_/A _5814_/X _6711_/S vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6071__S _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4828_ _8845_/A hold18/X vssd1 vssd1 vccd1 vccd1 _4828_/Y sky130_fd_sc_hd__nand2_1
X_7616_ _7700_/B _7609_/Y _7614_/Y _7754_/A _7615_/X vssd1 vssd1 vccd1 vccd1 _7616_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5167__A2 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6364__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8596_ _8596_/A vssd1 vssd1 vccd1 vccd1 _8596_/X sky130_fd_sc_hd__buf_1
XANTENNA__7561__B1 _7385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4759_ _4759_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4760_/B sky130_fd_sc_hd__nand2_1
X_7547_ _7547_/A _7691_/B vssd1 vssd1 vccd1 vccd1 _7547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8105__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7478_ _7477_/X _5496_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7479_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5923__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6429_ _6422_/X _4942_/X _6429_/S vssd1 vssd1 vccd1 vccd1 _6430_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput203 mports_i[77] vssd1 vssd1 vccd1 vccd1 _5511_/A sky130_fd_sc_hd__buf_2
XANTENNA__7616__A1 _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput214 mports_i[87] vssd1 vssd1 vccd1 vccd1 _5788_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__8813__B1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7616__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput225 mports_i[97] vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__buf_2
Xinput236 sports_i[105] vssd1 vssd1 vccd1 vccd1 _7814_/A1 sky130_fd_sc_hd__buf_4
Xinput247 sports_i[115] vssd1 vssd1 vccd1 vccd1 _7971_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput258 sports_i[125] vssd1 vssd1 vccd1 vccd1 _8106_/A1 sky130_fd_sc_hd__buf_4
Xinput269 sports_i[135] vssd1 vssd1 vccd1 vccd1 _8252_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7919__A2 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8041__A1 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8592__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6770__A _6770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5386__A _5386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8344__A2 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7077__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6355__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7855__A1 _7840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5833__B _7171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7855__B2 _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8804__B1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8280__A1 _7798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8280__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8032__A1 _5359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7776__A _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7386__A3 _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5800_ _6762_/A _6181_/B vssd1 vssd1 vccd1 vccd1 _5800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6780_ _6780_/A _6780_/B vssd1 vssd1 vccd1 vccd1 _6780_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6594__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7791__B1 _7791_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5731_ _5011_/Y _5721_/X _6755_/A _5997_/B _5730_/Y vssd1 vssd1 vccd1 vccd1 _5731_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5662_ _5662_/A vssd1 vssd1 vccd1 vccd1 _5662_/Y sky130_fd_sc_hd__inv_2
X_8450_ _8349_/A _8442_/Y _8443_/X _8449_/Y vssd1 vssd1 vccd1 vccd1 _8450_/X sky130_fd_sc_hd__o22a_2
XANTENNA__6346__A1 _4793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4613_ _4613_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__nand2_1
X_7401_ _7590_/A _7401_/B vssd1 vssd1 vccd1 vccd1 _7401_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8381_ _8364_/Y _8337_/Y _8380_/X vssd1 vssd1 vccd1 vccd1 _8381_/Y sky130_fd_sc_hd__o21ai_2
X_5593_ _4893_/A _5635_/A1 _4896_/A input42/X vssd1 vssd1 vccd1 vccd1 _5593_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7332_ _7332_/A _7332_/B vssd1 vssd1 vccd1 vccd1 _7332_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8099__A1 _8106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4544_ _4563_/B vssd1 vssd1 vccd1 vccd1 _8150_/A sky130_fd_sc_hd__buf_8
XANTENNA__8099__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8400__A _8400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6839__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7263_ _7263_/A vssd1 vssd1 vccd1 vccd1 _7263_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7846__A1 _8315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6649__A2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4475_ _4474_/Y _4326_/B _8189_/B vssd1 vssd1 vccd1 vccd1 _4476_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7016__A _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6214_ _6227_/A _8491_/B input4/X _4933_/A _6213_/X vssd1 vssd1 vccd1 vccd1 _7705_/B
+ sky130_fd_sc_hd__o221a_4
X_7194_ _6847_/A _7138_/X _7192_/X _7193_/X vssd1 vssd1 vccd1 vccd1 _7194_/X sky130_fd_sc_hd__o22a_2
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6145_ _5159_/B _6908_/A _6144_/X _5125_/X vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__a22o_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A vssd1 vssd1 vccd1 vccd1 _6076_/Y sky130_fd_sc_hd__inv_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5085__A1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5085__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5027_ input83/X _8706_/B input20/X _4940_/X vssd1 vssd1 vccd1 vccd1 _5027_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6821__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8559__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8023__A1 _8427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8023__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7686__A _7686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8970__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6590__A _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5388__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6978_ _6977_/X _7733_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6979_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5918__B _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8717_ _8824_/S vssd1 vssd1 vccd1 vccd1 _8820_/B sky130_fd_sc_hd__buf_4
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5929_ _5866_/A _8271_/A _5867_/A _5191_/X _5928_/X vssd1 vssd1 vccd1 vccd1 _6827_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8326__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6337__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8648_ _8647_/X _8782_/B _8689_/S vssd1 vssd1 vccd1 vccd1 _8648_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6337__B2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6888__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8579_ _8696_/A _8755_/C _8579_/C vssd1 vssd1 vccd1 vccd1 _8580_/A sky130_fd_sc_hd__and3_1
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8310__A _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6749__B _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7837__B2 _7707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5848__B1 _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5312__A2 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8456__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6273__B1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6812__A2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8014__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8565__A2 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5379__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4587__B1 _4557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5828__B _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6328__A1 _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4339__B1 _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6879__A2 _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5000__B2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5551__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6659__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput507 _6960_/X vssd1 vssd1 vccd1 vccd1 sports_o[104] sky130_fd_sc_hd__buf_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput518 _7319_/X vssd1 vssd1 vccd1 vccd1 sports_o[114] sky130_fd_sc_hd__buf_12
XFILLER_0_105_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput529 _7402_/X vssd1 vssd1 vccd1 vccd1 sports_o[124] sky130_fd_sc_hd__buf_12
XANTENNA__5839__B1 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7270__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7056__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5067__A1 _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7950_ _7958_/A1 _4946_/A _7958_/B1 _5119_/A vssd1 vssd1 vccd1 vccd1 _7950_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6901_ _7660_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6901_/Y sky130_fd_sc_hd__nand2_1
X_7881_ _7881_/A vssd1 vssd1 vccd1 vccd1 _7881_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8556__A2 _8157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4923__A _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6832_ _6827_/A _6801_/A _6824_/X _6826_/X _6831_/Y vssd1 vssd1 vccd1 vccd1 _6832_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_147_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7764__B1 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5738__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6763_ _5744_/X _7316_/A _8194_/A _5770_/X vssd1 vssd1 vccd1 vccd1 _6764_/A sky130_fd_sc_hd__a22o_1
XANTENNA__8308__A2 hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8502_ _8502_/A vssd1 vssd1 vccd1 vccd1 _8502_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6319__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5714_ _5909_/B _7148_/A _5713_/Y _5174_/A vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__a22o_1
XANTENNA__6319__B2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6694_ _6694_/A _6694_/B vssd1 vssd1 vccd1 vccd1 _6694_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5790__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8433_ _8433_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5527__C1 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5645_ _5645_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _5645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5576_ _5576_/A vssd1 vssd1 vccd1 vccd1 _5576_/Y sky130_fd_sc_hd__inv_2
X_8364_ _8364_/A vssd1 vssd1 vccd1 vccd1 _8364_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4527_ _4527_/A vssd1 vssd1 vccd1 vccd1 _4528_/B sky130_fd_sc_hd__inv_2
X_7315_ _7398_/A _7683_/B vssd1 vssd1 vccd1 vccd1 _7507_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8295_ _8295_/A _8336_/S vssd1 vssd1 vccd1 vccd1 _8295_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_130_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4458_ _4458_/A _4458_/B vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__nand2_1
X_7246_ _7246_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7246_/X sky130_fd_sc_hd__and2_1
X_7177_ _7177_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7177_/X sky130_fd_sc_hd__and2_1
X_4389_ _4389_/A vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__inv_2
X_6128_ _6128_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _6128_/Y sky130_fd_sc_hd__nand2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8244__A1 _8251_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8244__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__B1 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7452__C1 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6059_ _6059_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _6059_/Y sky130_fd_sc_hd__nand2_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7355__S _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5533__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6730__A1 _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6730__B2 _6732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5297__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6495__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7038__A2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8235__A1 _8235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8235__B2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8538__A2 _8364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4743__A _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7210__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output595_A _5376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4462__B hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5221__A1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5221__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5772__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7773__B _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5430_ input97/X _5192_/X input35/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5430_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5361_ _5361_/A vssd1 vssd1 vccd1 vccd1 _6626_/B sky130_fd_sc_hd__buf_8
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7100_ _6634_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7100_/X sky130_fd_sc_hd__a21o_1
X_4312_ _4337_/A _4312_/B vssd1 vssd1 vccd1 vccd1 _4313_/B sky130_fd_sc_hd__nand2_1
XANTENNA__7277__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8474__A1 _8491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8080_ _8080_/A1 _7876_/X _8080_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _8080_/Y sky130_fd_sc_hd__o22ai_2
X_5292_ _5292_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7031_ _7031_/A vssd1 vssd1 vccd1 vccd1 _7031_/X sky130_fd_sc_hd__buf_1
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7029__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8226__A1 _8235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8226__B2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8824__S _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7985__B1 _7985_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7933_ _7777_/X _7932_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _7933_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6852__B _6852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5460__A1 _5401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8529__A2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5460__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4653__A _8958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7864_ _7864_/A vssd1 vssd1 vccd1 vccd1 _7864_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_147_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6815_ _6924_/A _6815_/B vssd1 vssd1 vccd1 vccd1 _6815_/X sky130_fd_sc_hd__or2_1
XANTENNA__7201__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7795_ _7761_/A _7802_/A2 _8857_/B _4326_/B vssd1 vssd1 vccd1 vccd1 _7795_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8956__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6746_ _6746_/A vssd1 vssd1 vccd1 vccd1 _6746_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_135_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5763__A2 _7551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6960__A1 _6263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7683__B _7683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6677_ _6852_/A _7120_/A vssd1 vssd1 vccd1 vccd1 _6677_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7175__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8701__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8416_ _8416_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8416_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5628_ _5628_/A _7311_/A vssd1 vssd1 vccd1 vccd1 _7509_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_103_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6712__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8347_ _8345_/Y _8346_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8348_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5559_ _5558_/X _8181_/A _7311_/A _5544_/X vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__a22o_1
XANTENNA__7268__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8278_ _8277_/Y _7784_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8279_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5279__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5279__B2 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7229_ _6212_/B _7026_/X _7228_/X vssd1 vssd1 vccd1 vccd1 _7229_/X sky130_fd_sc_hd__o21a_1
XANTENNA__7204__A _7204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8217__A1 _4312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8217__B2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6779__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7858__B _7858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7440__A2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6762__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5451__A1 _5465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__B2 _6671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5659__A _5659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4563__A hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6400__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7874__A _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6951__A1 _6241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6951__B2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4962__B1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7900__B1 _7905_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6703__B2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6937__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6429__S _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8208__A1 _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4493__A2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output510_A _6975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output608_A _5706_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5442__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4930_ _8523_/B vssd1 vssd1 vccd1 vccd1 _4930_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4473__A _7818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5288__B _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7195__A1 _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4861_ hold5/X _4861_/B vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6600_ _6596_/X _6450_/X _6597_/X _6598_/Y _6599_/X vssd1 vssd1 vccd1 vccd1 _6600_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4792_ _4792_/A _4792_/B vssd1 vssd1 vccd1 vccd1 _4799_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7580_ _7581_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7580_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6942__A1 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6531_ _6525_/Y _6958_/B _6527_/X _6530_/X vssd1 vssd1 vccd1 vccd1 _6534_/A sky130_fd_sc_hd__a31o_1
XANTENNA__4920__B _7309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8695__A1 _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6462_ _6462_/A _6462_/B vssd1 vssd1 vccd1 vccd1 _6462_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_112_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8201_ _6081_/S _8198_/B _6231_/C vssd1 vssd1 vccd1 vccd1 _8201_/X sky130_fd_sc_hd__a21o_1
X_5413_ _6202_/B _6622_/A _5136_/X vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__o21a_1
X_6393_ _6400_/A1 _8310_/B input79/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8962__SET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8132_ _8132_/A1 _7876_/A _8132_/B1 _7835_/A vssd1 vssd1 vccd1 vccd1 _8132_/Y sky130_fd_sc_hd__o22ai_2
X_5344_ _6837_/A _5342_/X _5343_/X vssd1 vssd1 vccd1 vccd1 _5345_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5275_ _5275_/A vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__4648__A _8958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8063_ _8058_/Y _6965_/A _8059_/Y _8163_/A _8062_/Y vssd1 vssd1 vccd1 vccd1 _8464_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7014_ _7761_/A _8574_/B _7398_/A _4408_/B vssd1 vssd1 vccd1 vccd1 _7015_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_128_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7958__B1 _7958_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7678__B _7678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8965_ _8967_/CLK _8965_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__5433__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7916_ _7909_/Y _7769_/A _7910_/Y _6500_/A _7915_/Y vssd1 vssd1 vccd1 vccd1 _7916_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5984__A2 _6841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8896_ _4810_/B _4940_/X _4662_/C _8574_/B vssd1 vssd1 vccd1 vccd1 _8896_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7186__A1 _5885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7847_ _7847_/A _7858_/B vssd1 vssd1 vccd1 vccd1 _7847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7694__A _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7778_ _7874_/A _7778_/B vssd1 vssd1 vccd1 vccd1 _7778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6729_ _6729_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6729_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4830__B _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7489__A2 _5500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6249__S _6359_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4558__A _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput690 _6521_/X vssd1 vssd1 vccd1 vccd1 sports_o[64] sky130_fd_sc_hd__buf_12
XANTENNA__7661__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4475__A2 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8610__A1 _7869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8610__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5389__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4740__B _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 mports_i[111] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_2
Xinput25 mports_i[121] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput36 mports_i[131] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6013__A _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput47 mports_i[141] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_2
Xinput58 mports_i[151] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_1
XFILLER_0_134_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput69 mports_i[161] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_2
XANTENNA__6688__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7101__A1 _6635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4468__A _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5112__B1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5060_ _6281_/S _5060_/B vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__or2_1
XANTENNA__7652__A2 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6683__A _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7498__B _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8601__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7404__A2 _6578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5415__A1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5415__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8750_ _8833_/B _8366_/X _8725_/A vssd1 vssd1 vccd1 vccd1 _8750_/X sky130_fd_sc_hd__o21a_1
X_5962_ _5962_/A1 _5192_/X input55/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5962_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_59_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7701_ _7701_/A _7701_/B vssd1 vssd1 vccd1 vccd1 _7701_/Y sky130_fd_sc_hd__nor2_1
X_4913_ _4913_/A vssd1 vssd1 vccd1 vccd1 _4913_/X sky130_fd_sc_hd__buf_8
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8681_ _8552_/X _8581_/A _8549_/X _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8681_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7168__A1 _6770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5893_ _5893_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _5893_/X sky130_fd_sc_hd__and2_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4931__A _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5179__B1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7632_ _7694_/A _7632_/B vssd1 vssd1 vccd1 vccd1 _7632_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5718__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4844_ _8966_/D _4844_/B vssd1 vssd1 vccd1 vccd1 _4845_/C sky130_fd_sc_hd__nand2_1
XANTENNA__8403__A _8403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6915__A1 _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7563_ _7536_/A _7558_/Y _7559_/X _7562_/Y vssd1 vssd1 vccd1 vccd1 _7563_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6391__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8117__B1 _8111_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4775_ _8240_/A _8578_/A _4754_/Y _4773_/B vssd1 vssd1 vccd1 vccd1 _4776_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7019__A _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8668__A1 _8503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6514_ _6852_/A _6514_/B vssd1 vssd1 vccd1 vccd1 _6514_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8668__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7494_ _7510_/B _5645_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7494_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6445_ _6433_/X _6437_/Y _6439_/X _6443_/Y _6968_/A vssd1 vssd1 vccd1 vccd1 _6445_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__7340__A1 _5064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6143__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5762__A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5351__B1 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6376_ _6224_/S _7746_/B _6373_/X _6375_/Y vssd1 vssd1 vccd1 vccd1 _6376_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7891__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8115_ _8110_/Y _6965_/A _8111_/Y _8163_/A _8114_/Y vssd1 vssd1 vccd1 vccd1 _8510_/A
+ sky130_fd_sc_hd__a221oi_4
X_5327_ _8198_/A vssd1 vssd1 vccd1 vccd1 _8842_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__5103__B1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8840__A1 _8244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8046_ _8046_/A vssd1 vssd1 vccd1 vccd1 _8046_/Y sky130_fd_sc_hd__inv_2
X_5258_ input93/X _8709_/B input30/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6593__A _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5189_ _6560_/B _6133_/B vssd1 vssd1 vccd1 vccd1 _5189_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8053__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8971__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6603__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8948_ _8979_/CLK _8948_/D fanout732/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__5002__A _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7159__A1 _5765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8879_ _8886_/A _8894_/C _8899_/B vssd1 vssd1 vccd1 vccd1 _8879_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8356__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5937__A _5937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8659__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7599__A _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4560_ _4591_/B vssd1 vssd1 vccd1 vccd1 _4560_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_142_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4491_ _4727_/C hold36/A vssd1 vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__nand2_8
XANTENNA__7322__A1 _4966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6230_ _6227_/Y _8455_/B _6228_/Y _4891_/X _6229_/Y vssd1 vssd1 vccd1 vccd1 _6944_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7873__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6530__C1 _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5884__A1 _5902_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5884__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6965_/A _6931_/A vssd1 vssd1 vccd1 vccd1 _6161_/Y sky130_fd_sc_hd__nor2_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7086__A0 _7085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ input85/X _8368_/A input22/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5112_/X sky130_fd_sc_hd__o22a_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6092_/A vssd1 vssd1 vccd1 vccd1 _6092_/X sky130_fd_sc_hd__buf_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7625__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5636__A1 _5591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5064_/B _5230_/B _7536_/B _5109_/B _5042_/Y vssd1 vssd1 vccd1 vccd1 _6505_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6833__B1 _6832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7302__A _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8802_ _8499_/A _8806_/B _8800_/X _8801_/X vssd1 vssd1 vccd1 vccd1 _8802_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8050__A2 _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5939__A2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6994_ _6994_/A _6994_/B _6994_/C vssd1 vssd1 vccd1 vccd1 _6994_/X sky130_fd_sc_hd__or3_1
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6061__A1 _6061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6061__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8733_ _8733_/A _8833_/B vssd1 vssd1 vccd1 vccd1 _8733_/X sky130_fd_sc_hd__and2_1
X_5945_ _6007_/A1 _5090_/A input57/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5945_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_125_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8338__B1 _7916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4661__A _4661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8664_ _8664_/A vssd1 vssd1 vccd1 vccd1 _8664_/X sky130_fd_sc_hd__buf_1
XFILLER_0_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5347__A1_N _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5876_ _5870_/Y _5875_/Y _6081_/S vssd1 vssd1 vccd1 vccd1 _7592_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7615_ _6848_/A _7696_/B _6859_/A _7361_/X vssd1 vssd1 vccd1 vccd1 _7615_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4827_ _8857_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _4850_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6364__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8595_ _8594_/X _7784_/X _8686_/B vssd1 vssd1 vccd1 vccd1 _8596_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7546_ _7378_/X _5741_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7547_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4758_ _4758_/A _4823_/B vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7691__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7477_ _5498_/X _7696_/B _7475_/X _7326_/A _7476_/X vssd1 vssd1 vccd1 vccd1 _7477_/X
+ sky130_fd_sc_hd__a221o_1
X_4689_ _4734_/B _4689_/B vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6428_ _7001_/S vssd1 vssd1 vccd1 vccd1 _6429_/S sky130_fd_sc_hd__buf_6
XFILLER_0_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6521__C1 _6520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6359_ _6356_/X _6358_/X _6359_/S vssd1 vssd1 vccd1 vccd1 _6360_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput204 mports_i[78] vssd1 vssd1 vccd1 vccd1 _5506_/A sky130_fd_sc_hd__buf_2
XANTENNA__8813__A1 _8153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput215 mports_i[88] vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__clkbuf_4
Xinput226 mports_i[98] vssd1 vssd1 vccd1 vccd1 _6076_/A sky130_fd_sc_hd__buf_2
XANTENNA__5627__A1 _5601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5627__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput237 sports_i[106] vssd1 vssd1 vccd1 vccd1 _7827_/A sky130_fd_sc_hd__clkbuf_4
Xinput248 sports_i[116] vssd1 vssd1 vccd1 vccd1 _7985_/A1 sky130_fd_sc_hd__clkbuf_4
X_8029_ _8029_/A vssd1 vssd1 vccd1 vccd1 _8029_/Y sky130_fd_sc_hd__inv_2
Xinput259 sports_i[126] vssd1 vssd1 vccd1 vccd1 _8119_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6052__A1 _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6355__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7882__A _7882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7552__B2 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5563__B1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7855__A2 _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8804__A1 _8117_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5618__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5618__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8280__A2 _8429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output423_A _8213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8568__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6043__A1 _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7791__A1 _7791_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7791__B2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4481__A _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5730_ _6304_/A _6737_/A vssd1 vssd1 vccd1 vccd1 _5730_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5661_ _5661_/A vssd1 vssd1 vccd1 vccd1 _5661_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6346__A2 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8740__B1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7543__B2 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7400_ _7401_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7400_/Y sky130_fd_sc_hd__nand2_1
X_4612_ _4612_/A _4612_/B _4612_/C vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__nand3_1
X_8380_ _4913_/X _7972_/Y _4917_/X _7945_/Y vssd1 vssd1 vccd1 vccd1 _8380_/X sky130_fd_sc_hd__o22a_1
X_5592_ _5592_/A vssd1 vssd1 vccd1 vccd1 _5592_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7331_ _7756_/A vssd1 vssd1 vccd1 vccd1 _7332_/A sky130_fd_sc_hd__buf_8
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4543_ _8181_/A vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__inv_2
XANTENNA__8099__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8400__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5306__B1 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7262_ _6326_/X _7138_/A _7261_/X vssd1 vssd1 vccd1 vccd1 _7263_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__7846__A2 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4474_ _4474_/A _8166_/A vssd1 vssd1 vccd1 vccd1 _4474_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6213_ _6229_/A2 _8368_/A input66/X _4939_/A vssd1 vssd1 vccd1 vccd1 _6213_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7193_ _6841_/B _7019_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7193_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6144_ _6217_/B _6906_/B _6906_/A vssd1 vssd1 vccd1 vccd1 _6144_/X sky130_fd_sc_hd__mux2_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A vssd1 vssd1 vccd1 vccd1 _6075_/Y sky130_fd_sc_hd__inv_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5085__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6282__A1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6282__B2 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5026_ _6170_/A _5000_/X _5025_/X vssd1 vssd1 vccd1 vccd1 _5026_/X sky130_fd_sc_hd__a21bo_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8559__B1 _8219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8023__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6034__A1 _6059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _6976_/X _6337_/X _7000_/S vssd1 vssd1 vccd1 vccd1 _6977_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7782__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6082__S _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8716_ _8716_/A _8716_/B vssd1 vssd1 vccd1 vccd1 _8824_/S sky130_fd_sc_hd__nor2_8
XFILLER_0_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5928_ _5928_/A1 _5192_/X input54/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5793__B1 _5723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8647_ _8696_/A _8460_/A _8427_/A _8581_/A vssd1 vssd1 vccd1 vccd1 _8647_/X sky130_fd_sc_hd__a2bb2o_1
X_5859_ _5866_/A _4868_/A _5867_/A _4870_/A _5858_/X vssd1 vssd1 vccd1 vccd1 _5860_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6337__A2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5545__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8578_ _8578_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _8696_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7529_ _8759_/A _7529_/B vssd1 vssd1 vccd1 vccd1 _7529_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__8310__B _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7837__A2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5848__A1 _5772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5848__B2 _5824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6765__B _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4566__A _4566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6273__A1 _6286_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6273__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8014__A2 _8412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5233__C1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5397__A _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4587__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6981__C1 _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6328__A2 _7729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7525__B2 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5536__B1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5000__A2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5844__B _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput508 _6964_/X vssd1 vssd1 vccd1 vccd1 sports_o[105] sky130_fd_sc_hd__buf_12
XFILLER_0_151_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput519 _7323_/X vssd1 vssd1 vccd1 vccd1 sports_o[115] sky130_fd_sc_hd__buf_12
XFILLER_0_10_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5839__A1 _6811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5839__B2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__A _5860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8253__A2 _8252_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6900_ _7648_/B _6912_/B vssd1 vssd1 vccd1 vccd1 _6900_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8005__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7880_ _7760_/X _7867_/Y _7873_/X _7879_/X vssd1 vssd1 vccd1 vccd1 _7880_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_148_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6831_ _6831_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6831_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7764__A1 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7764__B2 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5775__B1 _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6762_ _6762_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6762_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5738__C _5738_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6972__C1 _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8501_ _8500_/X _8453_/A _8555_/B vssd1 vssd1 vccd1 vccd1 _8502_/A sky130_fd_sc_hd__mux2_1
X_5713_ _5713_/A vssd1 vssd1 vccd1 vccd1 _5713_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6319__A2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6693_ _5539_/X _5580_/X _6780_/A vssd1 vssd1 vccd1 vccd1 _6694_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7516__A1 _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8432_ _8431_/X _8782_/B _8496_/S vssd1 vssd1 vccd1 vccd1 _8432_/X sky130_fd_sc_hd__mux2_1
X_5644_ _5644_/A vssd1 vssd1 vccd1 vccd1 _7507_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8363_ _7956_/Y _8299_/A _8362_/X _8304_/A vssd1 vssd1 vccd1 vccd1 _8363_/X sky130_fd_sc_hd__a22o_1
X_5575_ _5575_/A vssd1 vssd1 vccd1 vccd1 _5575_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7314_ _7308_/X _4919_/X _7749_/S vssd1 vssd1 vccd1 vccd1 _7314_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4526_ _4526_/A _4526_/B vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8294_ _8567_/B vssd1 vssd1 vccd1 vccd1 _8564_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8557__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7245_ _7245_/A vssd1 vssd1 vccd1 vccd1 _7245_/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4457_ _4525_/A _4525_/C _4503_/B vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7176_ _7176_/A vssd1 vssd1 vccd1 vccd1 _7176_/X sky130_fd_sc_hd__buf_1
XANTENNA__6585__B _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4388_ _4392_/A _4393_/B _6231_/C vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__nand3_1
X_6127_ _6284_/A _7660_/A _5762_/A _6119_/Y _6126_/X vssd1 vssd1 vccd1 vccd1 _6128_/A
+ sky130_fd_sc_hd__o221ai_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8244__A2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5058__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6255__B2 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7452__B1 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6058_ _6058_/A vssd1 vssd1 vccd1 vccd1 _6058_/Y sky130_fd_sc_hd__inv_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _6470_/B _4986_/A _5008_/Y vssd1 vssd1 vccd1 vccd1 _6469_/B sky130_fd_sc_hd__o21ai_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6007__A1 _6007_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6007__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4569__A1 _4481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6106__A _6112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8704__B1 _8590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6540__S _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6715__C1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6730__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4741__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5297__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8235__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6246__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7443__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7994__B2 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5757__B1 _5788_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6016__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5221__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output490_A _7908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4980__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6182__B1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5360_ _6926_/A vssd1 vssd1 vccd1 vccd1 _6628_/B sky130_fd_sc_hd__buf_6
XFILLER_0_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4311_ _7847_/A _8180_/A vssd1 vssd1 vccd1 vccd1 _8185_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8377__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8960__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _6576_/B vssd1 vssd1 vccd1 vccd1 _5292_/A sky130_fd_sc_hd__inv_2
XFILLER_0_11_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6485__A1 _5064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7030_ _7029_/X _7332_/B _7097_/S vssd1 vssd1 vccd1 vccd1 _7031_/A sky130_fd_sc_hd__mux2_4
XANTENNA_hold23_A hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8226__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6237__A1 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7985__A1 _7985_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7985__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7932_ _7922_/Y _7874_/X _7923_/Y _7875_/X _7931_/Y vssd1 vssd1 vccd1 vccd1 _7932_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4934__A _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7310__A _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5460__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5749__B _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7863_ _7846_/X _7857_/Y _7760_/X _7862_/Y vssd1 vssd1 vccd1 vccd1 _7863_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_148_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6814_ _6801_/B _7536_/B _7707_/B _6828_/A vssd1 vssd1 vccd1 vccd1 _6815_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7794_ _7760_/X _7784_/X _7789_/X _7793_/X vssd1 vssd1 vccd1 vccd1 _7794_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_46_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6745_ _6906_/A _7529_/B _6743_/Y _6744_/Y vssd1 vssd1 vccd1 vccd1 _6746_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6960__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7683__C _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6676_ _7767_/A _7829_/A _8185_/B _5539_/X vssd1 vssd1 vccd1 vccd1 _6676_/X sky130_fd_sc_hd__or4b_1
X_8415_ _8555_/B _8413_/X _8414_/Y vssd1 vssd1 vccd1 vccd1 _8415_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5627_ _5601_/A _5102_/A _5602_/A _5191_/X _5626_/X vssd1 vssd1 vccd1 vccd1 _5628_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6712__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8346_ _8346_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5558_ _5505_/A _5102_/A _5506_/A _5191_/A _5557_/X vssd1 vssd1 vccd1 vccd1 _5558_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_130_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5920__B1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8287__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4509_ _4509_/A vssd1 vssd1 vccd1 vccd1 _7297_/B sky130_fd_sc_hd__buf_8
X_8277_ _8518_/B _8273_/X _8276_/Y vssd1 vssd1 vccd1 vccd1 _8277_/Y sky130_fd_sc_hd__a21oi_1
X_5489_ _5845_/B _5465_/Y _5484_/X _6133_/B _5488_/X vssd1 vssd1 vccd1 vccd1 _5490_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_112_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5279__A2 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6476__B2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7228_ _6192_/A _7004_/X _6931_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7228_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8217__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7159_ _5765_/X _7023_/X _7158_/X vssd1 vssd1 vccd1 vccd1 _7159_/X sky130_fd_sc_hd__o21a_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4844__A _8966_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5987__B1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5659__B _5827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7728__A1 _6326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6400__A1 _6400_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6400__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6951__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4962__A1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4962__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8153__A1 hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6164__B1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7900__A1 _7905_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7900__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5911__B1 _5937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7664__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8208__A2 _8198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6219__B2 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7967__B2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output503_A _6936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5442__A2 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _8934_/A _8934_/B _4860_/C vssd1 vssd1 vccd1 vccd1 _4861_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4791_ _4819_/A _4805_/B vssd1 vssd1 vccd1 vccd1 _4792_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6530_ _7368_/B _6925_/B _6563_/A _6871_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6530_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8144__A1 _8148_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6461_ _6461_/A vssd1 vssd1 vccd1 vccd1 _6462_/B sky130_fd_sc_hd__inv_2
XFILLER_0_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8200_ _8210_/A1 _6626_/B _8210_/B1 _6941_/A _8199_/X vssd1 vssd1 vccd1 vccd1 _8200_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5412_ _5412_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _5412_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6392_ _6401_/A1 _8516_/B input16/X _4913_/X _6391_/X vssd1 vssd1 vccd1 vccd1 _7754_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_113_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8131_ _8550_/A _7954_/X _8130_/Y _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8131_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _6780_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _5343_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7305__A _7532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7655__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8062_ _8067_/A1 _5146_/A _8067_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _8062_/Y sky130_fd_sc_hd__o22ai_2
X_5274_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__buf_6
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4648__B hold44/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4469__B1 hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7013_ _7013_/A vssd1 vssd1 vccd1 vccd1 _7761_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__7634__A2_N _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7407__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7958__A1 _7958_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7958__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8964_ _8967_/CLK hold28/X fanout733/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__5433__A2 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7915_ _7918_/A1 _5780_/X _7918_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7915_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8895_ _8894_/Y _4810_/A _8880_/Y vssd1 vssd1 vccd1 vccd1 _8898_/A sky130_fd_sc_hd__a21o_1
XANTENNA__4383__B _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7975__A _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7846_ _8315_/A _7872_/A _7975_/A vssd1 vssd1 vccd1 vccd1 _7846_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6918__C1 _6917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8383__A1 _7916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6394__B1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7777_ _7777_/A vssd1 vssd1 vccd1 vccd1 _7777_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4989_ _5056_/A _5174_/A _4986_/Y _4988_/X vssd1 vssd1 vccd1 vccd1 _4989_/X sky130_fd_sc_hd__a31o_1
XANTENNA__7186__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6728_ _5675_/Y _6912_/B _6724_/X _6726_/Y _6727_/Y vssd1 vssd1 vccd1 vccd1 _6729_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8135__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6659_ _7459_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6659_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7343__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7894__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8329_ _7886_/Y _8323_/X _8327_/X _8328_/Y vssd1 vssd1 vccd1 vccd1 _8329_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput680 _7291_/X vssd1 vssd1 vccd1 vccd1 sports_o[55] sky130_fd_sc_hd__buf_12
Xoutput691 _6534_/Y vssd1 vssd1 vccd1 vccd1 sports_o[65] sky130_fd_sc_hd__buf_12
XANTENNA__5121__A1 _5131_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8610__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__B _5425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8126__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput15 mports_i[112] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_2
Xwire730 _5132_/Y vssd1 vssd1 vccd1 vccd1 _6497_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput26 mports_i[122] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
Xinput37 mports_i[132] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6013__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 mports_i[142] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput59 mports_i[152] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7885__B1 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6948__B _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7125__A _7125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7101__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4468__B _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__A1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__A2 _5697_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8062__B1 _8067_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8601__A2 _8317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5415__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6612__A1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5299__B _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _5959_/X _6628_/B _5960_/Y vssd1 vssd1 vccd1 vccd1 _7619_/A sky130_fd_sc_hd__a21oi_2
X_7700_ _7701_/B _7700_/B vssd1 vssd1 vccd1 vccd1 _7700_/Y sky130_fd_sc_hd__nand2_1
X_4912_ _5191_/A vssd1 vssd1 vccd1 vccd1 _4913_/A sky130_fd_sc_hd__buf_8
XFILLER_0_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8680_ _8806_/A _8686_/B _8678_/X _8679_/Y vssd1 vssd1 vccd1 vccd1 _8680_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5892_ _6906_/A _5889_/Y _5891_/Y vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__8365__A1 _7906_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7168__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5179__A1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7631_ _7630_/Y _7297_/B _7575_/A _7385_/Y vssd1 vssd1 vccd1 vccd1 _7631_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5179__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4843_ hold10/X _8976_/D _4837_/A _4866_/A vssd1 vssd1 vccd1 vccd1 _4845_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8403__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7562_ _7767_/A _5750_/A _7561_/X vssd1 vssd1 vccd1 vccd1 _7562_/Y sky130_fd_sc_hd__o21ai_2
X_4774_ _5091_/A vssd1 vssd1 vccd1 vccd1 _8578_/A sky130_fd_sc_hd__inv_2
XANTENNA__8117__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6513_ _6513_/A vssd1 vssd1 vccd1 vccd1 _8163_/A sky130_fd_sc_hd__buf_12
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8668__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7493_ _7493_/A vssd1 vssd1 vccd1 vccd1 _7493_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6444_ _6946_/S vssd1 vssd1 vccd1 vccd1 _6968_/A sky130_fd_sc_hd__buf_6
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7340__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5351__A1 _6622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6375_ _6375_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5351__B2 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8114_ _8119_/A1 _5146_/A _8119_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _8114_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__7628__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5326_ input34/X _5111_/A _5326_/B1 _4931_/A _5325_/X vssd1 vssd1 vccd1 vccd1 _5328_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4378__B hold4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5103__A1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8045_ _8045_/A vssd1 vssd1 vccd1 vccd1 _8045_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5103__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5257_ _7422_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _5257_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8840__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5188_ _6593_/B _5184_/X _6547_/A vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__mux2_2
XANTENNA__8053__B1 _8458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7800__B1 _7802_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8947_ _8979_/CLK hold22/X fanout733/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8356__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8878_ hold18/X _8759_/A _8871_/A _8869_/B vssd1 vssd1 vccd1 vccd1 _8899_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_66_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7159__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7829_ _7829_/A _7829_/B vssd1 vssd1 vccd1 vccd1 _7829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8659__A2 _8068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5342__B2 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7095__A1 _5400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8292__B1 _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7095__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8831__A2 _8235_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8595__A1 _7784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6358__B1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4908__A1 _4876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4908__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6024__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4490_ hold15/X vssd1 vssd1 vccd1 vccd1 _4727_/C sky130_fd_sc_hd__clkinv_4
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4479__A _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5884__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6160_ _6157_/Y _4891_/X _6158_/Y _8455_/B _6159_/Y vssd1 vssd1 vccd1 vccd1 _6931_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5111_/A vssd1 vssd1 vccd1 vccd1 _8491_/B sky130_fd_sc_hd__buf_12
XANTENNA__7086__A1 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6088_/X _6095_/A _6224_/S vssd1 vssd1 vccd1 vccd1 _6092_/A sky130_fd_sc_hd__mux2_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6833__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5042_ _5106_/A _5042_/B vssd1 vssd1 vccd1 vccd1 _5042_/Y sky130_fd_sc_hd__nor2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8801_ _8833_/B _8107_/Y _8725_/A vssd1 vssd1 vccd1 vccd1 _8801_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6993_ _6993_/A vssd1 vssd1 vccd1 vccd1 _6993_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6061__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5944_ _5909_/B _5930_/Y _6851_/A _5174_/A vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__a22o_1
X_8732_ _7809_/X _8738_/A _7811_/X _8711_/A vssd1 vssd1 vccd1 vccd1 _8733_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8338__A1 _8352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8338__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6349__B1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8663_ _8662_/X _8476_/A _8690_/S vssd1 vssd1 vccd1 vccd1 _8664_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5875_ _6079_/A _6809_/B vssd1 vssd1 vccd1 vccd1 _5875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7010__A1 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7010__B2 _4408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7614_ _6841_/B _7542_/A _7694_/A _6854_/B _7613_/Y vssd1 vssd1 vccd1 vccd1 _7614_/Y
+ sky130_fd_sc_hd__o221ai_4
X_4826_ _8909_/S _4826_/B vssd1 vssd1 vccd1 vccd1 _4827_/B sky130_fd_sc_hd__nor2_1
X_8594_ _8593_/X _8272_/A _8621_/S vssd1 vssd1 vccd1 vccd1 _8594_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7561__A2 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7545_ _6747_/X _7361_/X _7543_/X _7754_/A _7544_/X vssd1 vssd1 vccd1 vccd1 _7545_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5572__A1 _5601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4757_ _4757_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4758_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5572__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7849__B1 _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7476_ _7476_/A _7476_/B vssd1 vssd1 vccd1 vccd1 _7476_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4688_ _4736_/A _4818_/B _4736_/B vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__nand3_2
X_6427_ _6448_/A vssd1 vssd1 vccd1 vccd1 _7001_/S sky130_fd_sc_hd__buf_8
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6358_ _6358_/A1 _4930_/X input13/X _4933_/X _6357_/X vssd1 vssd1 vccd1 vccd1 _6358_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__7077__A1 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8274__B1 _7788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5309_ _6875_/B _5306_/X _5308_/X vssd1 vssd1 vccd1 vccd1 _5310_/A sky130_fd_sc_hd__o21ai_1
Xinput205 mports_i[79] vssd1 vssd1 vccd1 vccd1 _5576_/A sky130_fd_sc_hd__buf_2
X_6289_ _6312_/A _7720_/B _6264_/X vssd1 vssd1 vccd1 vccd1 _6290_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__8813__A2 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput216 mports_i[89] vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_2_2__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__B1 _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput227 mports_i[99] vssd1 vssd1 vccd1 vccd1 _6141_/B1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5627__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6824__A1 _5860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput238 sports_i[107] vssd1 vssd1 vccd1 vccd1 _7840_/A sky130_fd_sc_hd__buf_1
X_8028_ _8028_/A vssd1 vssd1 vccd1 vccd1 _8028_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6824__B2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput249 sports_i[117] vssd1 vssd1 vccd1 vccd1 _7998_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5013__A _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5948__A _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6052__A2 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4852__A _8967_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8329__A1 _7886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7001__A1 _7756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7552__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5563__A1 _5635_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5563__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5315__A1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5315__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7068__A1 _5211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8804__A2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__buf_2
XANTENNA__4746__B _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6291__A2 _7720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output416_A _8096_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8568__A1 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5251__B1 _5266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7791__A2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4481__B _4481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5660_ _5660_/A _7384_/A vssd1 vssd1 vccd1 vccd1 _5660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8740__A1 _8315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7543__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4611_ _4611_/A _4611_/B vssd1 vssd1 vccd1 vccd1 _8846_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_154_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5591_ _5591_/A vssd1 vssd1 vccd1 vccd1 _5591_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_142_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7330_ _7330_/A vssd1 vssd1 vccd1 vccd1 _7756_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4542_ _8978_/Q vssd1 vssd1 vccd1 vccd1 _8181_/A sky130_fd_sc_hd__buf_8
XFILLER_0_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7261_ _6317_/X _7088_/A _6971_/X _7059_/A _7089_/A vssd1 vssd1 vccd1 vccd1 _7261_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5306__A1 _6578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5306__B2 _7413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4473_ _7818_/A vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__inv_2
X_6212_ _6212_/A _6212_/B vssd1 vssd1 vccd1 vccd1 _6212_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7192_ _7611_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7192_/X sky130_fd_sc_hd__and2_1
XFILLER_0_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6094_/X _6059_/B _8924_/B _6908_/A vssd1 vssd1 vccd1 vccd1 _6906_/B sky130_fd_sc_hd__a22o_1
XANTENNA__4937__A _4937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6806__A1 _6795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6074_/A vssd1 vssd1 vccd1 vccd1 _7209_/A sky130_fd_sc_hd__inv_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8008__B1 _8011_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6282__A2 _6283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _5010_/Y _5014_/Y _4925_/A _5017_/Y _5024_/Y vssd1 vssd1 vccd1 vccd1 _5025_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__7032__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8559__A1 _8217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8559__B2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6871__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6976_ _7266_/A _6994_/B _6333_/Y _6989_/B vssd1 vssd1 vccd1 vccd1 _6976_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7782__A2 _7763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5487__B _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8715_ _8738_/A vssd1 vssd1 vccd1 vccd1 _8803_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__5793__A1 _5722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5927_ _6628_/B _5925_/X _5926_/Y vssd1 vssd1 vccd1 vccd1 _7610_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__5793__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ _5928_/A1 _5090_/A input54/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5858_/X sky130_fd_sc_hd__o22a_1
X_8646_ _8412_/A _8577_/X _8644_/X _8645_/X vssd1 vssd1 vccd1 vccd1 _8646_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_36_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5545__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4809_ _4809_/A _4809_/B vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5789_ _5825_/A1 _5192_/X input51/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5789_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8577_ _8686_/B vssd1 vssd1 vccd1 vccd1 _8577_/X sky130_fd_sc_hd__buf_4
XFILLER_0_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7528_ _7606_/A _7528_/B vssd1 vssd1 vccd1 vccd1 _7528_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8495__B1 _8091_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7459_ _7459_/A _7696_/B vssd1 vssd1 vccd1 vccd1 _7459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5848__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5950__B _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6258__C1 _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6273__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__A3 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5481__B1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5233__B1 _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5397__B _5397_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4587__A2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5784__A1 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5784__B2 _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6981__B1 _6980_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7525__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5536__B2 _6679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7930__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput509 _6970_/X vssd1 vssd1 vccd1 vccd1 sports_o[106] sky130_fd_sc_hd__buf_12
XANTENNA_output366_A _7782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5839__A2 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5860__B _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8238__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4476__B _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7997__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7461__A1 _7458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8410__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6830_ _6798_/A _6829_/X _6870_/S vssd1 vssd1 vccd1 vccd1 _6831_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5224__B1 _5266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7764__A2 _7779_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5775__A1 _5741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6761_ _6761_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6761_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5775__B2 _5744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8500_ _8499_/Y _8476_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8500_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5712_ _6166_/B _5668_/X _5711_/X vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6692_ _5548_/X _6429_/S _6688_/X _6691_/X vssd1 vssd1 vccd1 vccd1 _6692_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_45_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8431_ _8426_/Y _8578_/B hold36/A _4727_/C _8430_/Y vssd1 vssd1 vccd1 vccd1 _8431_/X
+ sky130_fd_sc_hd__a41o_1
X_5643_ _5639_/Y _5642_/Y _8842_/B vssd1 vssd1 vccd1 vccd1 _5643_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5527__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8362_ _8713_/C _7901_/Y _8361_/Y _8513_/B vssd1 vssd1 vccd1 vccd1 _8362_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_72_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5574_ _5573_/X _5534_/A _6481_/B vssd1 vssd1 vccd1 vccd1 _5574_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6212__A _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7313_ _7715_/S vssd1 vssd1 vccd1 vccd1 _7749_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7027__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4525_ _4525_/A _4525_/B _4525_/C vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__nand3_1
X_8293_ _4933_/X _7821_/Y _4940_/X _7796_/X _8292_/X vssd1 vssd1 vccd1 vccd1 _8293_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7244_ _7243_/X _6248_/X _7249_/S vssd1 vssd1 vccd1 vccd1 _7245_/A sky130_fd_sc_hd__mux2_4
X_4456_ _4456_/A _4456_/B vssd1 vssd1 vccd1 vccd1 _4503_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7175_ _7174_/X _5824_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7176_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8139__A _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4387_ _4305_/Y _4377_/X _4300_/Y vssd1 vssd1 vccd1 vccd1 _4425_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__7043__A _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6126_ _6124_/X _5997_/B _6234_/B _6125_/Y vssd1 vssd1 vccd1 vccd1 _6126_/X sky130_fd_sc_hd__a211o_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4386__B _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__A2 _6262_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7452__A1 _6634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5058__A3 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6057_ _6133_/B _7648_/B _6055_/X _6233_/B _6056_/X vssd1 vssd1 vccd1 vccd1 _6057_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5008_ _5008_/A _6470_/B vssd1 vssd1 vccd1 vccd1 _5008_/Y sky130_fd_sc_hd__nand2_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6007__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5215__B1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7755__A2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4569__A2 _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5766__A1 _5765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6106__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6959_ _6467_/X _6261_/B _6450_/A vssd1 vssd1 vccd1 vccd1 _6959_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_49_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5010__B _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8704__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8629_ _8379_/X _8577_/X _8627_/X _8628_/Y vssd1 vssd1 vccd1 vccd1 _8629_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7435__A1_N _5094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7140__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6495__C _6497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6246__A2 _7707_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7443__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7994__A2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7400__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5206__B1 _7383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5757__A1 _5788_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5757__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6016__B _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4980__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6182__A1 _6182_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6182__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5871__A _5871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4310_ _4337_/A vssd1 vssd1 vccd1 vccd1 _7847_/A sky130_fd_sc_hd__inv_6
XANTENNA__7131__B1 _7130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5290_ _5159_/B _5239_/A _5125_/X _5241_/X _5289_/X vssd1 vssd1 vccd1 vccd1 _5290_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6178__S _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4496__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8393__S _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8631__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7985__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7931_ _7931_/A1 _7876_/X _7931_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7931_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_117_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7198__B1 _7197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7862_ _7862_/A vssd1 vssd1 vccd1 vccd1 _7862_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6207__A _6207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5111__A _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6813_ _6813_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6813_/Y sky130_fd_sc_hd__nand2_1
X_7793_ _7777_/X _8272_/A _7792_/X vssd1 vssd1 vccd1 vccd1 _7793_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4950__A _6359_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6744_ _6744_/A _6744_/B vssd1 vssd1 vccd1 vccd1 _6744_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_128_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6675_ _5496_/X _6429_/S _6674_/X vssd1 vssd1 vccd1 vccd1 _6675_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__8141__B _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5626_ _5640_/A1 _5192_/X input43/X _5193_/X vssd1 vssd1 vccd1 vccd1 _5626_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8414_ _8414_/A _8441_/B vssd1 vssd1 vccd1 vccd1 _8414_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5557_ _5557_/A1 _5192_/A input40/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5557_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5920__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8345_ _8345_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8345_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5381__C1 _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4508_ _8240_/A _4436_/A _4507_/Y _4506_/B vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8276_ _8299_/A _8274_/X _8275_/X _8304_/A _8496_/S vssd1 vssd1 vccd1 vccd1 _8276_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7122__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5488_ _6304_/A _6653_/A _7767_/A _5487_/Y _5715_/B vssd1 vssd1 vccd1 vccd1 _5488_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8965__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6088__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7227_ _7227_/A vssd1 vssd1 vccd1 vccd1 _7227_/X sky130_fd_sc_hd__buf_1
X_4439_ hold29/X vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__inv_2
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7158_ _7551_/A _7004_/X _5745_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7158_/X
+ sky130_fd_sc_hd__a221o_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7425__A1 _5356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6109_ _8150_/A _6914_/B _6108_/X vssd1 vssd1 vccd1 vccd1 _6110_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__7425__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7089_/A vssd1 vssd1 vccd1 vccd1 _7089_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5987__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8316__B _8364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7728__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5021__A _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6400__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4962__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6164__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7900__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8478__S _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5911__A1 _5936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5911__B2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7113__A0 _7112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7664__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6219__A2 _6185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8613__B1 _7890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7416__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7967__A2 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7411__A _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5978__A1 _5965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4754__B _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5978__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7719__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5866__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4790_ _4837_/A _4790_/B vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8144__A2 _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ _6994_/B vssd1 vssd1 vccd1 vccd1 _6899_/B sky130_fd_sc_hd__inv_6
XANTENNA__6155__A1 _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5411_ _6234_/B _7439_/B _5408_/Y _5410_/Y vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__a22o_1
X_6391_ _6400_/A1 _8716_/B input79/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6391_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5902__A1 _5902_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6697__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5902__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8130_ _8123_/Y _7769_/A _8124_/Y _6500_/A _8129_/Y vssd1 vssd1 vccd1 vccd1 _8130_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_101_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5342_ _5336_/Y _5299_/B _5390_/A _8140_/A vssd1 vssd1 vccd1 vccd1 _5342_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8061_ _8058_/Y _7013_/A _8059_/Y _5116_/A _8060_/Y vssd1 vssd1 vccd1 vccd1 _8491_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7655__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7305__B _7364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5273_ _5273_/A vssd1 vssd1 vccd1 vccd1 _5273_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7012_ _7009_/X _4919_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7012_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5106__A _5106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7407__A1 _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8604__B1 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5418__B1 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7958__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8080__A1 _8080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8963_ _8979_/CLK hold3/X fanout732/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__8080__B2 _7836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6091__A0 _6088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7914_ _7909_/Y _6965_/A _7910_/Y _8163_/A _7913_/Y vssd1 vssd1 vccd1 vccd1 _8352_/A
+ sky130_fd_sc_hd__a221oi_4
X_8894_ _8899_/B _8899_/C _8894_/C vssd1 vssd1 vccd1 vccd1 _8894_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7845_ _7840_/Y _7876_/A _7841_/Y _7835_/A _7844_/X vssd1 vssd1 vccd1 vccd1 _8315_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6394__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7776_ _7872_/A vssd1 vssd1 vccd1 vccd1 _7777_/A sky130_fd_sc_hd__inv_2
X_4988_ _7027_/A _5999_/B _5011_/A _6084_/B _6461_/A vssd1 vssd1 vccd1 vccd1 _4988_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7591__B1 _7587_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6727_ _6841_/A _6727_/B vssd1 vssd1 vccd1 vccd1 _6727_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8135__A2 _8523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6146__A1 _6135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6658_ _7470_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7894__A1 _8333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5609_ _6080_/A _5609_/B vssd1 vssd1 vccd1 vccd1 _5609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6589_ _6580_/Y _6450_/X _6583_/Y _6584_/Y _6588_/X vssd1 vssd1 vccd1 vccd1 _6589_/X
+ sky130_fd_sc_hd__a41o_1
X_8328_ _8333_/A _8518_/B _8323_/X vssd1 vssd1 vccd1 vccd1 _8328_/Y sky130_fd_sc_hd__a21oi_1
X_8259_ _8259_/A vssd1 vssd1 vccd1 vccd1 _8299_/A sky130_fd_sc_hd__inv_6
Xoutput670 _7245_/X vssd1 vssd1 vccd1 vccd1 sports_o[46] sky130_fd_sc_hd__buf_12
Xoutput681 _7296_/X vssd1 vssd1 vccd1 vccd1 sports_o[56] sky130_fd_sc_hd__buf_12
Xoutput692 _6556_/Y vssd1 vssd1 vccd1 vccd1 sports_o[66] sky130_fd_sc_hd__buf_12
XANTENNA__7231__A _7231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5686__A _5686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8950__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6281__S _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8126__A2 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 mports_i[113] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6137__A1 _6075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire731 _8094_/Y vssd1 vssd1 vccd1 vccd1 _8516_/A sky130_fd_sc_hd__clkbuf_4
Xinput27 mports_i[123] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
XFILLER_0_141_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput38 mports_i[133] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput49 mports_i[143] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7885__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6688__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output446_A _7839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output613_A _7025_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8062__A1 _8067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8062__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6980__A _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5960_ _6628_/B _5960_/B vssd1 vssd1 vccd1 vccd1 _5960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4911_ _8335_/B vssd1 vssd1 vccd1 vccd1 _8516_/B sky130_fd_sc_hd__clkbuf_16
X_5891_ _5891_/A _6906_/A vssd1 vssd1 vccd1 vccd1 _5891_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5596__A _5596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7630_ _7630_/A _7630_/B vssd1 vssd1 vccd1 vccd1 _7630_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5179__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4842_ _4842_/A _4842_/B vssd1 vssd1 vccd1 vccd1 _4866_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4773_ _4773_/A _4773_/B vssd1 vssd1 vccd1 vccd1 _4777_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7561_ _7560_/Y _7297_/B _7575_/A _7385_/Y vssd1 vssd1 vccd1 vccd1 _7561_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_71_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8117__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6512_ _6512_/A vssd1 vssd1 vccd1 vccd1 _6512_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7492_ _7491_/X _5548_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7493_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6443_ _6443_/A _6912_/B vssd1 vssd1 vccd1 vccd1 _6443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5535__S _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5887__B1 _5867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7316__A _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6374_ _6312_/A _7746_/B _6264_/X vssd1 vssd1 vccd1 vccd1 _6375_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5351__A2 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5325_ input93/X _4934_/A input30/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__o22a_1
X_8113_ _8110_/Y _7761_/A _8111_/Y _8857_/B _8112_/Y vssd1 vssd1 vccd1 vccd1 _8519_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7628__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5103__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5256_ _6440_/B vssd1 vssd1 vccd1 vccd1 _6544_/B sky130_fd_sc_hd__buf_8
X_8044_ _7975_/X _8439_/A _8040_/X _8043_/X vssd1 vssd1 vccd1 vccd1 _8044_/X sky130_fd_sc_hd__a22o_4
X_5187_ _6481_/B vssd1 vssd1 vccd1 vccd1 _6547_/A sky130_fd_sc_hd__buf_8
XANTENNA__8053__A1 _8455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8053__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7261__C1 _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7800__A1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6603__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8946_ _8979_/CLK _8946_/D fanout733/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__7800__B2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5811__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8877_ _8877_/A _8877_/B vssd1 vssd1 vccd1 vccd1 _8894_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8356__A2 _7945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7828_ _7836_/A vssd1 vssd1 vccd1 vccd1 _7828_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7564__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7759_ _7792_/A vssd1 vssd1 vccd1 vccd1 _7975_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8108__A2 _8107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6119__A1 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8967__D _8967_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7867__B2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5445__S _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5342__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8816__B1 _8169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8292__A1 _7763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7095__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6842__A2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8044__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7252__C1 _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5802__B1 _5801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6358__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8752__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4908__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6024__B _6074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6040__A _7660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6530__B2 _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5741_/B vssd1 vssd1 vccd1 vccd1 _5159_/B sky130_fd_sc_hd__buf_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6020_/A _5111_/A _6021_/A _4931_/A _6089_/X vssd1 vssd1 vccd1 vccd1 _6095_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6694__B _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6294__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _6507_/B vssd1 vssd1 vccd1 vccd1 _5042_/B sky130_fd_sc_hd__inv_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__A _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6186__S _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8035__B2 _7304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8800_ _8503_/A _8803_/B _8104_/Y _8711_/X _8788_/S vssd1 vssd1 vccd1 vccd1 _8800_/X
+ sky130_fd_sc_hd__a221o_1
X_6992_ _6991_/X _7746_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6993_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8731_ _8833_/B _8284_/B _8725_/X vssd1 vssd1 vccd1 vccd1 _8731_/Y sky130_fd_sc_hd__o21ai_1
X_5943_ _5942_/X _7592_/A _6711_/S vssd1 vssd1 vccd1 vccd1 _6851_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8338__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8662_ _8661_/X _8081_/Y _8689_/S vssd1 vssd1 vccd1 vccd1 _8662_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6215__A _7705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6349__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5874_ _5871_/Y _4886_/A _5872_/Y _4891_/A _5873_/Y vssd1 vssd1 vccd1 vccd1 _6809_/B
+ sky130_fd_sc_hd__o221a_2
XANTENNA__7546__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7010__A2 _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7613_ _7767_/A _5941_/A _7612_/X vssd1 vssd1 vccd1 vccd1 _7613_/Y sky130_fd_sc_hd__o21ai_1
X_4825_ _8869_/B _4825_/B vssd1 vssd1 vccd1 vccd1 _4826_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8593_ _7786_/X _8581_/A _7788_/X _8583_/A vssd1 vssd1 vccd1 vccd1 _8593_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7561__A3 _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7544_ _7544_/A _7696_/B vssd1 vssd1 vccd1 vccd1 _7544_/X sky130_fd_sc_hd__and2_1
XFILLER_0_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5572__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4756_ _4756_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7475_ _6671_/B _7660_/B _7473_/X _7348_/A _7474_/Y vssd1 vssd1 vccd1 vccd1 _7475_/X
+ sky130_fd_sc_hd__a221o_1
X_4687_ _4687_/A hold33/X vssd1 vssd1 vccd1 vccd1 _4736_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6426_ _6426_/A _6511_/A vssd1 vssd1 vccd1 vccd1 _6448_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6521__A1 _7356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6521__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6357_ _6357_/A1 _8706_/B input75/X _4940_/X vssd1 vssd1 vccd1 vccd1 _6357_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5308_ _6481_/B _5308_/B vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__or2_1
X_6288_ _6285_/X _6287_/X _6386_/S vssd1 vssd1 vccd1 vccd1 _6288_/X sky130_fd_sc_hd__mux2_1
Xinput206 mports_i[7] vssd1 vssd1 vccd1 vccd1 _5139_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5088__A1 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__B2 _5150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput217 mports_i[8] vssd1 vssd1 vccd1 vccd1 _5195_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput228 mports_i[9] vssd1 vssd1 vccd1 vccd1 _5208_/A1 sky130_fd_sc_hd__clkbuf_4
X_8027_ _7975_/X _8433_/A _8023_/X _8026_/X vssd1 vssd1 vccd1 vccd1 _8027_/X sky130_fd_sc_hd__a22o_4
XANTENNA__6824__A2 _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput239 sports_i[108] vssd1 vssd1 vccd1 vccd1 _7877_/A1 sky130_fd_sc_hd__clkbuf_4
X_5239_ _5239_/A _5361_/A vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__and2_1
XANTENNA__8026__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__B2 _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6037__B1 _5989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5013__B _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6588__A1 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7785__B1 _7304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6588__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6052__A3 _6897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8929_ _8929_/A _8929_/B vssd1 vssd1 vccd1 vccd1 _8930_/C sky130_fd_sc_hd__nor2_1
XANTENNA__4852__B _8966_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8329__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6125__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7537__B1 _7535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5964__A _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5563__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5315__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8017__A1 _8024_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8017__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8568__A2 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8515__A _8515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output409_A _8014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5251__B2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6200__B1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8740__A2 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4610_ _4610_/A _4610_/B vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5590_ _5590_/A vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__buf_1
XFILLER_0_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4541_ _4557_/B _4591_/B vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7260_ _7260_/A vssd1 vssd1 vccd1 vccd1 _7260_/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5306__A2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4472_ _4331_/B _4518_/A _4611_/B _6440_/B vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6211_ _6211_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _6211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_150_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7191_ _7191_/A vssd1 vssd1 vccd1 vccd1 _7191_/X sky130_fd_sc_hd__buf_1
XFILLER_0_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6185_/A _8924_/B _6059_/B _7683_/A vssd1 vssd1 vccd1 vccd1 _6217_/B sky130_fd_sc_hd__a22o_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6547_/A _6133_/A _6072_/Y vssd1 vssd1 vccd1 vccd1 _6912_/A sky130_fd_sc_hd__o21ai_2
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6806__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5762_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5024_/Y sky130_fd_sc_hd__nor2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8008__A1 _8011_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8008__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8559__A2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4953__A _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _6975_/A vssd1 vssd1 vccd1 vccd1 _6975_/X sky130_fd_sc_hd__buf_2
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8714_ _8714_/A vssd1 vssd1 vccd1 vccd1 _8738_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5926_ _6628_/B _5926_/B vssd1 vssd1 vccd1 vccd1 _5926_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5793__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7519__B1 _5628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8645_ _8698_/B _8012_/Y _8590_/X vssd1 vssd1 vccd1 vccd1 _8645_/X sky130_fd_sc_hd__o21a_1
X_5857_ _6811_/B vssd1 vssd1 vccd1 vccd1 _5857_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8731__A2 _8284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4808_ _4808_/A _7511_/B vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__nand2_1
XANTENNA__8160__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5545__A2 _5544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8576_ _8690_/S vssd1 vssd1 vccd1 vccd1 _8686_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6742__A1 _5741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5788_ _5788_/A1 _8271_/A _5788_/B1 _4913_/A _5787_/X vssd1 vssd1 vccd1 vccd1 _6770_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6742__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7527_ _6731_/B _7361_/X _7525_/X _7326_/A _7526_/Y vssd1 vssd1 vccd1 vccd1 _7527_/X
+ sky130_fd_sc_hd__a221o_1
X_4739_ _6342_/A vssd1 vssd1 vccd1 vccd1 _6980_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8495__A1 _8511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8495__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7458_ _5423_/X _7680_/B _7457_/X vssd1 vssd1 vccd1 vccd1 _7458_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5008__B _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6409_ _6434_/B _7302_/B vssd1 vssd1 vccd1 vccd1 _6475_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7389_ _7389_/A vssd1 vssd1 vccd1 vccd1 _7696_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8798__A2 _8516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5024__A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5481__A1 _5738_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5481__B2 _7551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8335__A _8335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5233__A1 _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6981__A1 _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6981__B2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__B1 _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7930__B1 _7929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7289__A2 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8238__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7997__B1 _8424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7461__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5472__A1 _5637_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5472__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6464__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8410__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5224__B2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6760_ _6760_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6760_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6972__A1 _6317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5775__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6972__B2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5711_ _6711_/S _5752_/B vssd1 vssd1 vccd1 vccd1 _5711_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6691_ _5558_/X _6801_/A _6924_/A _6690_/Y _6450_/A vssd1 vssd1 vccd1 vccd1 _6691_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7295__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8430_ _8428_/X _8513_/B _8429_/Y vssd1 vssd1 vccd1 vccd1 _8430_/Y sky130_fd_sc_hd__a21oi_1
X_5642_ _5679_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5642_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5527__A2 _5498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8361_ _8361_/A vssd1 vssd1 vccd1 vccd1 _8361_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5573_ _5552_/X _7299_/A _6281_/S _5659_/A vssd1 vssd1 vccd1 vccd1 _5573_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6212__B _6212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5109__A _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7312_ _7681_/A _7673_/A vssd1 vssd1 vccd1 vccd1 _7715_/S sky130_fd_sc_hd__nand2_4
X_4524_ _4524_/A _4549_/A vssd1 vssd1 vccd1 vccd1 _4839_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8292_ _7763_/X hold31/A _8759_/B vssd1 vssd1 vccd1 vccd1 _8292_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7243_ _7707_/D _7138_/X _7241_/X _7242_/X vssd1 vssd1 vccd1 vccd1 _7243_/X sky130_fd_sc_hd__o22a_1
X_4455_ _4455_/A _4455_/B vssd1 vssd1 vccd1 vccd1 _4456_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4948__A _5893_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5160__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4386_ _4386_/A _7510_/B vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__nand2_1
X_7174_ _6788_/B _7138_/X _7172_/X _7173_/X vssd1 vssd1 vccd1 vccd1 _7174_/X sky130_fd_sc_hd__o22a_2
X_6125_ _6304_/A _6897_/A vssd1 vssd1 vccd1 vccd1 _6125_/Y sky130_fd_sc_hd__nor2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6056_ _6016_/A _5845_/B _6386_/S vssd1 vssd1 vccd1 vccd1 _6056_/X sky130_fd_sc_hd__a21o_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7452__A2 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5463__A1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5463__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5007_ _6965_/A _6474_/A vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__nor2_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5215__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6963__A1 _7720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6958_ _6958_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5909_ _7183_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5909_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6889_ _6889_/A _6933_/A vssd1 vssd1 vccd1 vccd1 _6889_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8704__A2 _8252_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8628_ _8381_/Y _8685_/B _8686_/B vssd1 vssd1 vccd1 vccd1 _8628_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6715__A1 _5628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7218__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6122__B _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8559_ _8217_/X _8304_/X _8219_/X _8299_/X _8496_/S vssd1 vssd1 vccd1 vccd1 _8559_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6191__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7140__A1 _5659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8640__A1 _8403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7443__A2 _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8640__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5689__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5206__A1 _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5206__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5757__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4965__B1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8156__B1 _8158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7409__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6706__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6182__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7131__A1 _5562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7682__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8631__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8092__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7930_ _8359_/A _7768_/X _7929_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7930_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7861_ _7840_/Y _4947_/B _7841_/Y _5123_/A _7860_/X vssd1 vssd1 vccd1 vccd1 _7862_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_77_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7198__A1 _6868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6207__B _6868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6812_ _7584_/A _6912_/B _6808_/Y _6810_/Y _6811_/Y vssd1 vssd1 vccd1 vccd1 _6813_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_147_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7792_ _7792_/A vssd1 vssd1 vccd1 vccd1 _7792_/X sky130_fd_sc_hd__buf_4
XANTENNA__6945__A1 _6234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6945__B2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6743_ _6743_/A _8924_/B vssd1 vssd1 vccd1 vccd1 _6743_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8147__B1 _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6674_ _6667_/X _6871_/B _6672_/X _6467_/X _6673_/Y vssd1 vssd1 vccd1 vccd1 _6674_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8413_ _8412_/Y _8390_/Y _8875_/B vssd1 vssd1 vccd1 vccd1 _8413_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5625_ _5625_/A vssd1 vssd1 vccd1 vccd1 _7526_/B sky130_fd_sc_hd__inv_2
XFILLER_0_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8344_ _7932_/Y _8564_/B _8343_/X vssd1 vssd1 vccd1 vccd1 _8344_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__5381__B1 _5400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5556_ _5550_/X _6233_/B _6170_/A _5555_/X vssd1 vssd1 vccd1 vccd1 _5556_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5920__A2 _5885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5781__B _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4507_ _6440_/B _6342_/A vssd1 vssd1 vccd1 vccd1 _4507_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8275_ _7786_/X _8257_/C _8579_/C _8232_/X vssd1 vssd1 vccd1 vccd1 _8275_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7122__A1 _6679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5487_ _5487_/A _6837_/A vssd1 vssd1 vccd1 vccd1 _5487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7226_ _7225_/X _7683_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7227_/A sky130_fd_sc_hd__mux2_2
XANTENNA__6476__A3 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4438_ _8945_/Q vssd1 vssd1 vccd1 vccd1 _8584_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4397__B _7683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7157_ _7157_/A vssd1 vssd1 vccd1 vccd1 _7157_/X sky130_fd_sc_hd__buf_1
X_4369_ hold34/X vssd1 vssd1 vccd1 vccd1 _4715_/B sky130_fd_sc_hd__inv_2
XANTENNA__8622__A1 _7912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7425__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6108_ _8151_/B _6108_/B vssd1 vssd1 vccd1 vccd1 _6108_/X sky130_fd_sc_hd__or2_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7088_/A vssd1 vssd1 vccd1 vccd1 _7088_/X sky130_fd_sc_hd__buf_6
X_6039_ _6047_/A _5080_/A _6048_/A _5089_/X _6038_/X vssd1 vssd1 vccd1 vccd1 _7660_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5987__A2 _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7189__A1 _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8386__B1 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6936__A1 _6185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8689__A1 _8211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5911__A2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6787__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7113__A1 _5464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5124__B1 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7664__A2 _6094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5675__A1 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6872__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8613__A1 _7888_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7416__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8613__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5427__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5427__B2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5978__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5212__A _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8523__A _8523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6927__A1 _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output593_A _5290_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8129__B1 _8132_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5410_ _5011_/Y _5409_/Y _5013_/Y vssd1 vssd1 vccd1 vccd1 _5410_/Y sky130_fd_sc_hd__o21ai_1
X_6390_ _6386_/X _6402_/A _6389_/Y vssd1 vssd1 vccd1 vccd1 _6390_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5902__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6697__B _6697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5341_ _6024_/A _7094_/A vssd1 vssd1 vccd1 vccd1 _5390_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8060_ _8067_/A1 _4946_/A _8067_/B1 _5119_/A vssd1 vssd1 vccd1 vccd1 _8060_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__7655__A2 _6095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5272_ _5272_/A vssd1 vssd1 vccd1 vccd1 _5272_/Y sky130_fd_sc_hd__inv_2
X_7011_ _7089_/A vssd1 vssd1 vccd1 vccd1 _7012_/S sky130_fd_sc_hd__buf_8
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8604__A1 _7837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7407__A2 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5418__A1 _5440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5418__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7812__C1 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8962_ _8979_/CLK hold6/X fanout732/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfstp_1
XANTENNA__8080__A2 _7876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5122__A _7352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6091__A1 _6095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7913_ _7918_/A1 _5146_/A _7918_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _7913_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8893_ _8893_/A _8893_/B vssd1 vssd1 vccd1 vccd1 _8899_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7844_ _7842_/Y _7843_/Y hold12/A vssd1 vssd1 vccd1 vccd1 _7844_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_66_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8433__A _8433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5776__B _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7775_ _7765_/X _7768_/X _7771_/X _7772_/X _7774_/X vssd1 vssd1 vccd1 vccd1 _7775_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6394__A2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ _7384_/A _5096_/A vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6726_ _6432_/X _6725_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6726_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6146__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6657_ _6655_/X _6933_/A _6968_/A _6656_/X vssd1 vssd1 vccd1 vccd1 _6657_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_6_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7343__B2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5608_ _5600_/Y _8140_/A _6456_/B _5607_/Y vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__a31o_1
XANTENNA__7894__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6588_ _5239_/A _6510_/A _6587_/Y _6512_/X vssd1 vssd1 vccd1 vccd1 _6588_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8327_ _7888_/Y _8304_/X _7890_/Y _8299_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8327_/X
+ sky130_fd_sc_hd__a221o_1
X_5539_ _6470_/B _5514_/Y _5538_/Y vssd1 vssd1 vccd1 vccd1 _5539_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_131_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8258_ _8429_/A vssd1 vssd1 vccd1 vccd1 _8304_/A sky130_fd_sc_hd__buf_6
Xoutput660 _7204_/X vssd1 vssd1 vccd1 vccd1 sports_o[37] sky130_fd_sc_hd__buf_12
Xoutput671 _7250_/X vssd1 vssd1 vccd1 vccd1 sports_o[47] sky130_fd_sc_hd__buf_12
X_7209_ _7209_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7209_/X sky130_fd_sc_hd__and2_1
XFILLER_0_111_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput682 _6430_/X vssd1 vssd1 vccd1 vccd1 sports_o[57] sky130_fd_sc_hd__buf_12
Xoutput693 _6572_/X vssd1 vssd1 vccd1 vccd1 sports_o[67] sky130_fd_sc_hd__buf_12
X_8189_ _8189_/A _8189_/B _8189_/C vssd1 vssd1 vccd1 vccd1 _8189_/X sky130_fd_sc_hd__and3_1
XANTENNA__7512__A _7512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4871__A _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5593__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 mports_i[114] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
XFILLER_0_25_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 mports_i[124] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_2
XFILLER_0_107_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 mports_i[134] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5896__A1 _5962_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5896__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8834__A1 _8226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7422__A _7422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4765__B _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8598__B1 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output606_A _5650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8062__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6073__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4484__C _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4910_ _5102_/A vssd1 vssd1 vccd1 vccd1 _8335_/B sky130_fd_sc_hd__buf_12
XFILLER_0_87_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _5824_/X _7316_/A _8924_/B _5853_/X vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4841_ _4841_/A _4841_/B vssd1 vssd1 vccd1 vccd1 _4842_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_114_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7560_ _7560_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7560_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4772_ _4772_/A vssd1 vssd1 vccd1 vccd1 _4773_/B sky130_fd_sc_hd__inv_2
XFILLER_0_117_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6781__C1 _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6511_ _6511_/A vssd1 vssd1 vccd1 vccd1 _6512_/A sky130_fd_sc_hd__inv_2
XFILLER_0_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7491_ _7487_/X _7488_/Y _7489_/X _7490_/X vssd1 vssd1 vccd1 vccd1 _7491_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_43_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6442_ _6876_/C vssd1 vssd1 vccd1 vccd1 _6912_/B sky130_fd_sc_hd__buf_6
XFILLER_0_130_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5887__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5887__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6373_ _6170_/A _6364_/X _6372_/X vssd1 vssd1 vccd1 vccd1 _6373_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5117__A _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8112_ _8119_/A1 _4947_/B _8119_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _8112_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_140_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8825__A1 _8200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5324_ _7415_/B _6181_/B vssd1 vssd1 vccd1 vccd1 _5324_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7628__A2 _6059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8043_ _7777_/X _8042_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _8043_/X sky130_fd_sc_hd__o21ba_1
X_5255_ _5272_/A _4953_/X _5273_/A _5089_/X _5254_/X vssd1 vssd1 vccd1 vccd1 _7422_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__4956__A _4956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7332__A _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5186_ _6793_/S vssd1 vssd1 vccd1 vccd1 _6481_/B sky130_fd_sc_hd__inv_6
XANTENNA__8053__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7800__A2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8945_ _8978_/CLK _8945_/D fanout732/X vssd1 vssd1 vccd1 vccd1 _8945_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6890__B _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5811__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7478__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8163__A _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8876_ _8875_/Y _4811_/B _8870_/B vssd1 vssd1 vccd1 vccd1 _8877_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7827_ _7827_/A vssd1 vssd1 vccd1 vccd1 _7827_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7564__A1 _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7758_ _8759_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _7792_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_19_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6709_ _5568_/Y _6924_/A _6704_/X _6708_/X vssd1 vssd1 vccd1 vccd1 _6709_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7689_ _7687_/X _7754_/A _7688_/X vssd1 vssd1 vccd1 vccd1 _7689_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_144_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7867__A2 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6411__A _6411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5878__A1 _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5878__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8816__A1 _8165_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput490 _7908_/X vssd1 vssd1 vccd1 vccd1 mports_o[8] sky130_fd_sc_hd__buf_12
XANTENNA__7242__A _7242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8044__A2 _8439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6055__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6055__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5802__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6358__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8752__B1 _8386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5869__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6040__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6530__A2 _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8807__A1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output723_A _6874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5371__S _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__A1 _6336_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5131_/A2 _8335_/B _5131_/B2 _4913_/A _5039_/X vssd1 vssd1 vccd1 vccd1 _6507_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6294__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__B _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8035__A2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6991_ _6990_/X _6364_/X _7000_/S vssd1 vssd1 vccd1 vccd1 _6991_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7794__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8730_ _7796_/X _8806_/B _8728_/X _8729_/Y vssd1 vssd1 vccd1 vccd1 _8730_/X sky130_fd_sc_hd__a22o_1
X_5942_ _8140_/A _5970_/A _5941_/Y vssd1 vssd1 vccd1 vccd1 _5942_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5400__A _5400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8661_ _8483_/A _8581_/A _8480_/A _8583_/A vssd1 vssd1 vccd1 vccd1 _8661_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6349__A2 _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5873_ _5274_/X _5902_/A1 _5275_/X input53/X vssd1 vssd1 vccd1 vccd1 _5873_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__7546__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6215__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7612_ _7611_/Y _7297_/B _7694_/A _7385_/Y vssd1 vssd1 vccd1 vccd1 _7612_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5557__B1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4824_ _8877_/B _4824_/B _8870_/B vssd1 vssd1 vccd1 vccd1 _4825_/B sky130_fd_sc_hd__nand3_1
X_8592_ _7763_/X _8577_/X _8588_/X _8591_/X vssd1 vssd1 vccd1 vccd1 _8592_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7543_ _5482_/X _7680_/B _7541_/X _7640_/B _7542_/Y vssd1 vssd1 vccd1 vccd1 _7543_/X
+ sky130_fd_sc_hd__a221o_2
X_4755_ _8240_/A _8256_/A _4754_/Y _4752_/B vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6231__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7474_ _7575_/A _7474_/B vssd1 vssd1 vccd1 vccd1 _7474_/Y sky130_fd_sc_hd__nor2_1
X_4686_ _8239_/A _4686_/B vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6425_ _8857_/B _8574_/B vssd1 vssd1 vccd1 vccd1 _6511_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6521__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6356_ _6353_/X _6355_/X _6356_/S vssd1 vssd1 vccd1 vccd1 _6356_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5307_ _7422_/A _7299_/A _6281_/S _5094_/A vssd1 vssd1 vccd1 vccd1 _5308_/B sky130_fd_sc_hd__a22o_1
XANTENNA__8274__A2 _8230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4686__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ _6287_/A1 _8516_/B input7/X _4913_/X _6286_/X vssd1 vssd1 vccd1 vccd1 _6287_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__8158__A _8158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput207 mports_i[80] vssd1 vssd1 vccd1 vccd1 _5592_/A sky130_fd_sc_hd__buf_2
XANTENNA__6285__A1 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__A2 _6499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput218 mports_i[90] vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6285__B2 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8026_ _7777_/X _8782_/B _7792_/X vssd1 vssd1 vccd1 vccd1 _8026_/X sky130_fd_sc_hd__o21ba_1
Xinput229 nrst_i vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_8
X_5238_ _7316_/A vssd1 vssd1 vccd1 vccd1 _6059_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__4835__A2 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8026__A2 _8782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5169_ _6558_/B vssd1 vssd1 vccd1 vccd1 _7071_/A sky130_fd_sc_hd__inv_2
XANTENNA__6037__A1 _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6037__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7785__A1 _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6588__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7785__B2 _7790_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8928_ _4848_/A _4847_/A hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__o21ai_1
XANTENNA__6406__A _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7001__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6125__B _6897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8859_ _8856_/Y _4601_/A _8858_/X vssd1 vssd1 vccd1 vccd1 _8969_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__7537__A1 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5548__B1 _5506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5980__A _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6276__A1 _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6276__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8017__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6579__A2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8515__B _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5251__A2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6200__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4540_ _4863_/B vssd1 vssd1 vccd1 vccd1 _8945_/D sky130_fd_sc_hd__inv_2
XFILLER_0_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4471_ _7852_/A _8189_/B vssd1 vssd1 vccd1 vccd1 _6440_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8963__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6210_ _6870_/S _6204_/Y _6209_/Y vssd1 vssd1 vccd1 vccd1 _6211_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7190_ _7189_/X _5899_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7191_/A sky130_fd_sc_hd__mux2_2
X_6141_ _6141_/A1 _4929_/A _6141_/B1 _4932_/A _6140_/X vssd1 vssd1 vccd1 vccd1 _7683_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6197__S _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6072_/A _6481_/B vssd1 vssd1 vccd1 vccd1 _6072_/Y sky130_fd_sc_hd__nand2_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _8189_/A _5060_/B _5022_/X vssd1 vssd1 vccd1 vccd1 _5024_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__8008__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8706__A _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7216__A0 _7215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6974_ _6973_/X _7729_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6226__A _7705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5130__A _5130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8713_ _8755_/A _8755_/C _8713_/C vssd1 vssd1 vccd1 vccd1 _8714_/A sky130_fd_sc_hd__and3_1
XFILLER_0_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5925_ _5923_/Y _5924_/Y _8842_/B vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6990__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7519__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8644_ _8416_/A _8581_/X _8009_/Y _8583_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8644_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6660__S _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5856_ _5856_/A _6481_/B vssd1 vssd1 vccd1 vccd1 _5863_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8959__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4807_ _4607_/A _4748_/B _8584_/A _4793_/Y _4806_/B vssd1 vssd1 vccd1 vccd1 _4808_/A
+ sky130_fd_sc_hd__a41o_1
X_8575_ _8590_/A vssd1 vssd1 vccd1 vccd1 _8690_/S sky130_fd_sc_hd__inv_2
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5787_ _5787_/A1 _8271_/B input50/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5787_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8160__B _8172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6742__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7526_ _7681_/A _7526_/B vssd1 vssd1 vccd1 vccd1 _7526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4738_ _4738_/A _4738_/B vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7457_ _6648_/B _7660_/B _7456_/X _7640_/B vssd1 vssd1 vccd1 vccd1 _7457_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8495__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4669_ _4372_/A _4668_/B _4406_/A vssd1 vssd1 vccd1 vccd1 _4670_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6408_ _6415_/A vssd1 vssd1 vccd1 vccd1 _6994_/B sky130_fd_sc_hd__buf_8
XFILLER_0_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7388_ _6550_/A _7542_/A _6560_/B _7694_/A _7387_/X vssd1 vssd1 vccd1 vccd1 _7388_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6339_ _6312_/A _7733_/B _6264_/X vssd1 vssd1 vccd1 vccd1 _6340_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5305__A _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6258__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7455__B1 _6630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8009_ _8002_/Y _7769_/X _8003_/Y _6500_/X _8008_/Y vssd1 vssd1 vccd1 vccd1 _8009_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7207__A0 _7206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7520__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5481__A2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8335__B _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6966__C1 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5233__A2 _6566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6981__A2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__A1 _4975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8351__A _8351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4992__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8183__A1 _8189_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8183__B2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6194__B1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7930__A1 _8359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7930__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8497__S _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8238__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6249__A1 _6248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7997__A1 _8403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7997__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output421_A _8177_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5472__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8410__A2 _7999_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5224__A2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6972__A2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5710_ _5689_/Y _5523_/A _8160_/A vssd1 vssd1 vccd1 vccd1 _5752_/B sky130_fd_sc_hd__mux2_1
X_6690_ _7483_/B vssd1 vssd1 vccd1 vccd1 _6690_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6709__C1 _6708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ _5601_/A _4929_/A _5602_/A _4932_/A _5640_/X vssd1 vssd1 vccd1 vccd1 _5679_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7921__A1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8360_ _8358_/Y _8359_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8361_/A sky130_fd_sc_hd__mux2_1
X_5572_ _5601_/A _4953_/X _5602_/A _5089_/X _5571_/X vssd1 vssd1 vccd1 vccd1 _5659_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_122_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7311_ _7311_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _7673_/A sky130_fd_sc_hd__nand2_8
X_4523_ _4603_/B _4602_/B vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5109__B _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8291_ _8555_/B vssd1 vssd1 vccd1 vccd1 _8759_/B sky130_fd_sc_hd__clkinv_4
XFILLER_0_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7134__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7242_ _7242_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7242_/X sky130_fd_sc_hd__and2_1
X_4454_ _4454_/A _4454_/B vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5160__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7173_ _5827_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7173_/X sky130_fd_sc_hd__a21o_1
X_4385_ _8239_/A _7304_/A _4412_/C vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__nand3_1
XANTENNA__5125__A _5893_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6124_ _6053_/Y _6123_/Y _6166_/B vssd1 vssd1 vccd1 vccd1 _6124_/X sky130_fd_sc_hd__mux2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7988__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _5909_/B _7639_/A _6054_/X _5997_/B vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__a22o_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5006_ _5003_/Y _4891_/X _5004_/Y _8455_/B _5005_/Y vssd1 vssd1 vccd1 vccd1 _6474_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__5463__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6957_ _6252_/X _6933_/A _6956_/X vssd1 vssd1 vccd1 vccd1 _6958_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5908_ _6809_/B vssd1 vssd1 vccd1 vccd1 _7183_/A sky130_fd_sc_hd__inv_2
XANTENNA__8171__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6888_ _7209_/A _6475_/X _6026_/X _6694_/B vssd1 vssd1 vccd1 vccd1 _6889_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5839_ _6811_/B _8188_/S _5682_/B _5879_/A vssd1 vssd1 vccd1 vccd1 _5839_/X sky130_fd_sc_hd__a22o_1
X_8627_ _8384_/X _8583_/A _8386_/X _8581_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8627_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6715__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7912__B2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8558_ _8558_/A vssd1 vssd1 vccd1 vccd1 _8558_/X sky130_fd_sc_hd__buf_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5019__B _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7509_ _7509_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _7509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8489_ _8323_/X _8479_/Y _8487_/X _8488_/X vssd1 vssd1 vccd1 vccd1 _8489_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6479__A1 _5028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7140__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7979__B2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4874__A _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6100__B1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8346__A _8346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8640__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7250__A _7250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6651__B2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5689__B _6737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4593__B _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5206__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4965__A1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4965__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8156__A1 _8172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8156__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6706__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7903__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7131__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5142__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7419__B1 _7359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8092__B1 _8091_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8631__A2 _8765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7860_ _7858_/Y _7859_/Y hold44/A vssd1 vssd1 vccd1 vccd1 _7860_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7198__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6811_ _6841_/A _6811_/B vssd1 vssd1 vccd1 vccd1 _6811_/Y sky130_fd_sc_hd__nor2_1
X_7791_ _7791_/A1 _8174_/A _7791_/B1 _5230_/B _7790_/X vssd1 vssd1 vccd1 vccd1 _8272_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6945__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6742_ _5741_/A _6908_/B _5720_/X _6512_/X _6741_/X vssd1 vssd1 vccd1 vccd1 _6742_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6504__A _6528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8147__A1 _8151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6673_ _6506_/A _5498_/X _6449_/A vssd1 vssd1 vccd1 vccd1 _6673_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5624_ _5596_/A _5102_/A _5597_/A _5191_/A _5623_/X vssd1 vssd1 vccd1 vccd1 _5625_/A
+ sky130_fd_sc_hd__o221a_4
X_8412_ _8412_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8412_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8343_ _8359_/A _8304_/A _7929_/Y _8299_/A _8496_/S vssd1 vssd1 vccd1 vccd1 _8343_/X
+ sky130_fd_sc_hd__a221o_1
X_5555_ _5845_/B _5500_/X _5554_/X _6133_/B vssd1 vssd1 vccd1 vccd1 _5555_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5381__A1 _6634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5381__B2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5554__S _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4506_ _4506_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7658__B1 _7654_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8274_ _8578_/A _8230_/Y _7788_/X vssd1 vssd1 vccd1 vccd1 _8274_/X sky130_fd_sc_hd__a21o_1
X_5486_ _5405_/Y _5444_/Y _6470_/B vssd1 vssd1 vccd1 vccd1 _5487_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7122__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7225_ _6180_/A _7138_/X _7223_/X _7224_/X vssd1 vssd1 vccd1 vccd1 _7225_/X sky130_fd_sc_hd__o22a_1
X_4437_ _4437_/A vssd1 vssd1 vccd1 vccd1 _8977_/D sky130_fd_sc_hd__buf_1
X_7156_ _7155_/X _5741_/A _7175_/S vssd1 vssd1 vccd1 vccd1 _7157_/A sky130_fd_sc_hd__mux2_1
X_4368_ _4706_/B _4810_/B vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6107_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6108_/B sky130_fd_sc_hd__nand2_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _7087_/A vssd1 vssd1 vccd1 vccd1 _7087_/X sky130_fd_sc_hd__buf_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4395_/B _4394_/B vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__nand2_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6104_/A1 _8709_/B input61/X _5091_/X vssd1 vssd1 vccd1 vccd1 _6038_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7830__B1 _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7920__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8386__A1 _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7189__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8386__B2 _8404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6397__B1 _6400_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8974__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7989_ _7989_/A vssd1 vssd1 vccd1 vccd1 _7989_/Y sky130_fd_sc_hd__inv_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5729__S _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6936__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6133__B _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4869__A _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7245__A _7245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7649__B1 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5124__A1 _7356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5124__B2 _7345_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6872__A1 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8613__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6624__A1 _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5427__A2 _7451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6624__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6388__B1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8523__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8129__A1 _8132_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8129__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7139__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output586_A _5127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5340_ _5337_/Y _4885_/A _5338_/Y _4890_/A _5339_/Y vssd1 vssd1 vccd1 vccd1 _7094_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8082__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5115__A1 _5139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5115__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5271_ _6081_/S vssd1 vssd1 vccd1 vccd1 _7829_/A sky130_fd_sc_hd__buf_8
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7010_ _7874_/A _8584_/B _7510_/A _4408_/B vssd1 vssd1 vccd1 vccd1 _7089_/A sky130_fd_sc_hd__a22o_4
XANTENNA__5418__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6615__A1 _6608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7812__B1 _7811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8961_ _8979_/CLK _8961_/D fanout732/X vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfrtp_4
X_7912_ _7909_/Y _7761_/A _7910_/Y _8857_/B _7911_/Y vssd1 vssd1 vccd1 vccd1 _7912_/Y
+ sky130_fd_sc_hd__a221oi_4
X_8892_ _8892_/A _8892_/B vssd1 vssd1 vccd1 vccd1 _8973_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7843_ _8181_/A _7859_/B vssd1 vssd1 vccd1 vccd1 _7843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8433__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6918__A2 _6511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6234__A _6234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4986_ _4986_/A _6470_/B vssd1 vssd1 vccd1 vccd1 _4986_/Y sky130_fd_sc_hd__nand2_1
X_7774_ _7872_/A vssd1 vssd1 vccd1 vccd1 _7774_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7591__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6725_ _6852_/A _7532_/B vssd1 vssd1 vccd1 vccd1 _6725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6656_ _5465_/A _6913_/B _5423_/X _6912_/B vssd1 vssd1 vccd1 vccd1 _6656_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7343__A2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5607_ _5607_/A vssd1 vssd1 vccd1 vccd1 _5607_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5354__A1 _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6587_ _6587_/A vssd1 vssd1 vccd1 vccd1 _6587_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8326_ _7867_/Y _8323_/X _8324_/X _8325_/X vssd1 vssd1 vccd1 vccd1 _8326_/X sky130_fd_sc_hd__a22o_1
X_5538_ _5538_/A vssd1 vssd1 vccd1 vccd1 _5538_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8595__S _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8257_ _8259_/A _8755_/C _8257_/C vssd1 vssd1 vccd1 vccd1 _8429_/A sky130_fd_sc_hd__and3_2
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5469_ _6671_/B _5077_/A _6017_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput650 _7161_/X vssd1 vssd1 vccd1 vccd1 sports_o[28] sky130_fd_sc_hd__buf_12
Xoutput661 _7208_/X vssd1 vssd1 vccd1 vccd1 sports_o[38] sky130_fd_sc_hd__buf_12
X_7208_ _7208_/A vssd1 vssd1 vccd1 vccd1 _7208_/X sky130_fd_sc_hd__buf_1
Xoutput672 _7256_/X vssd1 vssd1 vccd1 vccd1 sports_o[48] sky130_fd_sc_hd__buf_12
Xoutput683 _6452_/X vssd1 vssd1 vccd1 vccd1 sports_o[58] sky130_fd_sc_hd__buf_12
X_8188_ _8180_/A _8192_/A _8188_/S vssd1 vssd1 vccd1 vccd1 _8188_/X sky130_fd_sc_hd__mux2_1
Xoutput694 _6589_/X vssd1 vssd1 vccd1 vccd1 sports_o[68] sky130_fd_sc_hd__buf_12
X_7139_ _7514_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7139_/X sky130_fd_sc_hd__and2_1
XANTENNA__6409__A _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7803__B1 _7803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6606__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6128__B _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__B1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7582__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5593__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5593__B2 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6790__B1 _5824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 mports_i[115] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__8531__A1 _8137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6798__B _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 mports_i[125] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5896__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8819__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5648__A2 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8518__B _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7422__B _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8598__A1 _8297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output501_A _7921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4840_ _4839_/Y hold1/X _7309_/B vssd1 vssd1 vccd1 vccd1 _4841_/A sky130_fd_sc_hd__a21o_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4771_ _4771_/A _4771_/B vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__nand2_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6510_ _6510_/A vssd1 vssd1 vccd1 vccd1 _6908_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7490_ _5558_/X _7389_/A _6701_/B _7476_/B vssd1 vssd1 vccd1 vccd1 _7490_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6441_ _6854_/A vssd1 vssd1 vccd1 vccd1 _6876_/C sky130_fd_sc_hd__inv_6
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5887__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6372_ _6234_/B _6367_/Y _5762_/A _6370_/X _6371_/X vssd1 vssd1 vccd1 vccd1 _6372_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4302__A _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8111_ _8111_/A vssd1 vssd1 vccd1 vccd1 _8111_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5323_ _5323_/A vssd1 vssd1 vccd1 vccd1 _7415_/B sky130_fd_sc_hd__inv_2
XFILLER_0_140_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8709__A _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8042_ _8028_/Y _5230_/B _8029_/Y _7536_/B _8041_/X vssd1 vssd1 vccd1 vccd1 _8042_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__6836__A1 _5899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5254_ input94/X _8709_/B input31/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5254_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7332__B _7332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5185_ _5185_/A _7769_/A vssd1 vssd1 vccd1 vccd1 _6793_/S sky130_fd_sc_hd__nor2_4
XANTENNA__5133__A _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7261__A1 _6317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7261__B2 _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8944_ _8978_/CLK _8944_/D fanout732/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__8444__A _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5811__A2 _5825_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4691__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8875_ _8875_/A _8875_/B vssd1 vssd1 vccd1 vccd1 _8875_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8210__B1 _8210_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7826_ _7826_/A vssd1 vssd1 vccd1 vccd1 _7826_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7564__A2 _5770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4969_ _4978_/B _5090_/A _4977_/B _4874_/A vssd1 vssd1 vccd1 vccd1 _4969_/X sky130_fd_sc_hd__o22a_1
X_7757_ _7755_/X _7332_/A _7756_/Y vssd1 vssd1 vccd1 vccd1 _7757_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6708_ _6706_/X _6899_/B _7000_/S _6707_/X vssd1 vssd1 vccd1 vccd1 _6708_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7688_ _7673_/A _6179_/A _6212_/B _7389_/A vssd1 vssd1 vccd1 vccd1 _7688_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6639_ _6632_/Y _6467_/X _6633_/Y _6634_/Y _6638_/X vssd1 vssd1 vccd1 vccd1 _6639_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_62_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5308__A _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8309_ _4891_/X _7851_/Y _4894_/A _7809_/X _8308_/X vssd1 vssd1 vccd1 vccd1 _8309_/X
+ sky130_fd_sc_hd__o221a_2
Xoutput480 _8632_/X vssd1 vssd1 vccd1 vccd1 mports_o[80] sky130_fd_sc_hd__buf_12
Xoutput491 _8667_/X vssd1 vssd1 vccd1 vccd1 mports_o[90] sky130_fd_sc_hd__buf_12
XANTENNA__7242__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7252__B2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5802__A2 _5770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8201__B1 _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5015__B1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8752__A1 _8384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8752__B2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6763__B1 _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6321__B _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5218__A _5218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5869__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4776__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7243__A1 _7707_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8264__A _8264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6990_ _7743_/A _6994_/B _6989_/X vssd1 vssd1 vccd1 vccd1 _6990_/X sky130_fd_sc_hd__a21o_1
XANTENNA__7794__A2 _7784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _5941_/A vssd1 vssd1 vccd1 vccd1 _5941_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_88_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5872_ _5872_/A vssd1 vssd1 vccd1 vccd1 _5872_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_125_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8660_ _8491_/A _8577_/X _8658_/X _8659_/X vssd1 vssd1 vccd1 vccd1 _8660_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7546__A2 _5741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4823_ _8887_/A _4823_/B _8887_/B vssd1 vssd1 vccd1 vccd1 _8870_/B sky130_fd_sc_hd__nand3_1
X_7611_ _7611_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7611_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5557__A1 _5557_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5557__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8591_ _8698_/B _8295_/A _8590_/X vssd1 vssd1 vccd1 vccd1 _8591_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4754_ hold32/A _6342_/A vssd1 vssd1 vccd1 vccd1 _4754_/Y sky130_fd_sc_hd__nor2_1
X_7542_ _7542_/A _7542_/B vssd1 vssd1 vccd1 vccd1 _7542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5309__A1 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7473_ _7115_/A _7630_/B _5538_/Y _8755_/C vssd1 vssd1 vccd1 vccd1 _7473_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6231__B _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4685_ _4685_/A _7272_/B vssd1 vssd1 vccd1 vccd1 _4686_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7703__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5128__A _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6424_ _6510_/A vssd1 vssd1 vccd1 vccd1 _6426_/A sky130_fd_sc_hd__inv_2
XFILLER_0_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6355_ _6358_/A1 _8516_/B input13/X _4913_/X _6354_/X vssd1 vssd1 vccd1 vccd1 _6355_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8439__A _8439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5306_ _6578_/B _5682_/B _8188_/S _7413_/A vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__a22o_1
X_6286_ _6286_/A1 _8716_/B input70/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6286_/X sky130_fd_sc_hd__o22a_1
Xinput208 mports_i[81] vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__buf_2
XANTENNA__7482__A1 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5237_ _5237_/A vssd1 vssd1 vccd1 vccd1 _7316_/A sky130_fd_sc_hd__clkbuf_16
X_8025_ _8015_/Y _7874_/X _8016_/Y _7875_/X _8024_/Y vssd1 vssd1 vccd1 vccd1 _8782_/B
+ sky130_fd_sc_hd__a221oi_4
Xinput219 mports_i[91] vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__buf_2
XANTENNA__5493__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5168_ input28/X _4896_/A input91/X _4893_/A _5167_/X vssd1 vssd1 vccd1 vccd1 _6558_/B
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__6037__A2 _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8174__A _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5099_ _6489_/A _5845_/B _6386_/S vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5245__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7785__A2 _7790_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8927_ _8927_/A vssd1 vssd1 vccd1 vccd1 _8959_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__6406__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8858_ _4600_/A _4600_/B _8857_/Y _6264_/X vssd1 vssd1 vccd1 vccd1 _8858_/X sky130_fd_sc_hd__a31o_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8734__A1 _7807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5548__A1 _5505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7809_ _7814_/A1 _5171_/B _7814_/B1 _5299_/B _7808_/X vssd1 vssd1 vccd1 vccd1 _7809_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5548__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8789_ _8502_/Y _8759_/Y _8788_/X _8725_/X vssd1 vssd1 vccd1 vccd1 _8789_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6568__S _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__A1 _6743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4877__A _6312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8349__A _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__B2 _5741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4596__B _4596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6276__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7473__B2 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__buf_2
XANTENNA__7225__A1 _6180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7700__B _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5236__B1 _5266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5787__A1 _5787_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5787__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5539__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6736__B1 _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output499_A _8694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7428__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6051__B _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4470_ _8189_/B _8166_/A vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_111_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6140_ _6140_/A1 _4935_/A input63/X _4939_/A vssd1 vssd1 vccd1 vccd1 _6140_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_21_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7464__A1 _5460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6676__D_N _5539_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6071_ _6116_/B _6040_/Y _8189_/A vssd1 vssd1 vccd1 vccd1 _6133_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8661__B1 _8480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _8188_/S _5022_/B vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__or2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8706__B _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7216__A1 _6094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7610__B _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6507__A _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5227__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6973_ _6326_/X _6467_/X _6972_/X vssd1 vssd1 vccd1 vccd1 _6973_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8712_ _8712_/A vssd1 vssd1 vccd1 vccd1 _8755_/A sky130_fd_sc_hd__inv_2
X_5924_ _5924_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5924_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8722__A _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8643_ _8643_/A vssd1 vssd1 vccd1 vccd1 _8643_/X sky130_fd_sc_hd__buf_1
XFILLER_0_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5855_ _5855_/A vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__inv_2
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4806_ _4806_/A _4806_/B vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__nand2_1
X_8574_ _8574_/A _8574_/B vssd1 vssd1 vccd1 vccd1 _8590_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5786_ _5780_/X _5782_/Y _6284_/A _6758_/B _5785_/X vssd1 vssd1 vccd1 vccd1 _5786_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7525_ _5674_/X _7680_/B _7523_/X _7348_/A _7524_/X vssd1 vssd1 vccd1 vccd1 _7525_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4737_ _4737_/A vssd1 vssd1 vccd1 vccd1 _4738_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7456_ _7105_/A _7668_/B _5487_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _7456_/X sky130_fd_sc_hd__a22o_1
X_4668_ _4668_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4670_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6407_ _6462_/A _6854_/A vssd1 vssd1 vccd1 vccd1 _6415_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_141_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4599_ _4599_/A _7309_/B vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__nand2_1
X_7387_ _6557_/A _7638_/B _7386_/X vssd1 vssd1 vccd1 vccd1 _7387_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6338_ _6335_/X _6337_/X _6386_/S vssd1 vssd1 vccd1 vccd1 _6338_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6258__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6269_ _6286_/A1 _8706_/B input70/X _4940_/A vssd1 vssd1 vccd1 vccd1 _6269_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8652__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7455__B2 _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8008_ _8011_/A1 _5780_/X _8011_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _8008_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__7207__A1 _6058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6417__A _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7012__S _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5769__A1 _5792_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5769__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8351__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8183__A2 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6194__A1 _6229_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6194__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7930__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5457__B1 _5402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7997__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output414_A _8070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8261__B _8584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5640_ _5640_/A1 _4935_/A input43/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_116_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7921__A2 _7912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5571_ _5640_/A1 _8709_/B input43/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5571_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_143_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4522_ _4596_/B _4601_/B vssd1 vssd1 vccd1 vccd1 _4602_/B sky130_fd_sc_hd__nand2_1
X_7310_ _7389_/A vssd1 vssd1 vccd1 vccd1 _7681_/A sky130_fd_sc_hd__inv_4
XFILLER_0_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8290_ _8491_/B _8368_/A vssd1 vssd1 vccd1 vccd1 _8555_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7241_ _6241_/X _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7241_/X sky130_fd_sc_hd__a21o_1
X_4453_ _4453_/A _7852_/A vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__nand2_1
XANTENNA__8882__B1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7685__B2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7172_ _7172_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7172_/X sky130_fd_sc_hd__and2_1
XANTENNA__5160__A2 _5195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4384_ _8160_/A _6231_/C vssd1 vssd1 vccd1 vccd1 _7304_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6123_ _7829_/A _7678_/B _6122_/Y vssd1 vssd1 vccd1 vccd1 _6123_/Y sky130_fd_sc_hd__o21ai_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7437__A1 _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8717__A _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5448__B1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7988__A2 _8390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6054_ _5995_/X _6053_/Y _6780_/A vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__mux2_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _4893_/A input83/X _4896_/A input20/X vssd1 vssd1 vccd1 vccd1 _5005_/Y sky130_fd_sc_hd__a22oi_1
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6956_ _6456_/B _7246_/A _6851_/B _6955_/Y vssd1 vssd1 vccd1 vccd1 _6956_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5907_ _7767_/A _6780_/A _6807_/B vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__or3_1
XFILLER_0_49_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6887_ _6058_/A _6908_/B _6884_/X _6886_/Y vssd1 vssd1 vccd1 vccd1 _6887_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8626_ _8372_/X _8577_/X _8624_/X _8625_/X vssd1 vssd1 vccd1 vccd1 _8626_/X sky130_fd_sc_hd__a22o_1
X_5838_ _5804_/A _4868_/A _5805_/A _5089_/A _5837_/X vssd1 vssd1 vccd1 vccd1 _5879_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7912__A2 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8557_ _8554_/X _8556_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8558_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5769_ _5792_/A1 _4934_/A input49/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5769_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_133_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7508_ _5651_/X _7619_/B _7505_/X _7506_/X _7507_/Y vssd1 vssd1 vccd1 vccd1 _7508_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8488_ _8564_/B _8081_/Y _8497_/S vssd1 vssd1 vccd1 vccd1 _8488_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6479__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7676__A1 _7683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7439_ _7542_/A _7439_/B vssd1 vssd1 vccd1 vccd1 _7439_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7676__B2 _7359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5687__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5316__A _6102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8625__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7979__A2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6100__A1 _6136_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6100__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8346__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6651__A2 _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6403__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8953__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4890__A _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4965__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8156__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6167__A1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7903__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5925__S _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7116__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7667__A1 _7663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5678__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5142__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output629_A _6220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7441__A _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8092__A1 _8511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8092__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8256__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6810_ _6432_/X _6809_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6810_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__8272__A _8272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7790_ _7874_/A _7790_/A2 _7311_/A _7790_/B2 vssd1 vssd1 vccd1 vccd1 _7790_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6741_ _5704_/Y _6924_/A _6736_/X _6740_/X vssd1 vssd1 vccd1 vccd1 _6741_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8147__A2 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6672_ _5454_/B _6876_/C _6668_/Y _6670_/Y _6671_/Y vssd1 vssd1 vccd1 vccd1 _6672_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8411_ _8323_/X _8402_/X _8409_/X _8410_/X vssd1 vssd1 vccd1 vccd1 _8411_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_45_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5623_ _5637_/A1 _5192_/A input44/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8342_ _8342_/A vssd1 vssd1 vccd1 vccd1 _8342_/X sky130_fd_sc_hd__buf_1
XFILLER_0_143_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5554_ _5501_/X _5553_/X _6593_/A vssd1 vssd1 vccd1 vccd1 _5554_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5381__A2 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7658__A1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4505_ _4505_/A vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__inv_2
X_8273_ _4917_/X _8235_/Y _8364_/A _8316_/A vssd1 vssd1 vccd1 vccd1 _8273_/X sky130_fd_sc_hd__o22a_1
X_5485_ _5485_/A vssd1 vssd1 vccd1 vccd1 _7767_/A sky130_fd_sc_hd__buf_8
XANTENNA__5136__A _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4436_ _4436_/A _4436_/B vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__or2_1
X_7224_ _7678_/B _7288_/B vssd1 vssd1 vccd1 vccd1 _7224_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4975__A _4975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4367_ hold35/X vssd1 vssd1 vccd1 vccd1 _4706_/B sky130_fd_sc_hd__inv_2
X_7155_ _7544_/A _7138_/X _7153_/X _7154_/X vssd1 vssd1 vccd1 vccd1 _7155_/X sky130_fd_sc_hd__o22a_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8083__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6112_/B _6868_/B vssd1 vssd1 vccd1 vccd1 _6914_/B sky130_fd_sc_hd__nand2_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7085_/X _5362_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7087_/A sky130_fd_sc_hd__mux2_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4416_/B _4601_/B vssd1 vssd1 vccd1 vccd1 _4394_/B sky130_fd_sc_hd__nand2_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ _5988_/A _8491_/B _5989_/A _4933_/A _6036_/X vssd1 vssd1 vccd1 vccd1 _6058_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8386__A2 _8351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6397__A1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6397__B2 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7988_ _7975_/X _8390_/A _7984_/X _7987_/X vssd1 vssd1 vccd1 vccd1 _7988_/X sky130_fd_sc_hd__a22o_2
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7594__B1 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6939_ _7696_/A _6517_/B _6938_/X vssd1 vssd1 vccd1 vccd1 _6939_/X sky130_fd_sc_hd__o21a_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8609_ _8609_/A vssd1 vssd1 vccd1 vccd1 _8609_/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7526__A _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6430__A _6430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7649__A1 _7532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5046__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5124__A2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4885__A _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6872__A2 _6867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8074__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6624__A2 _6510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _8979_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6388__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7585__B1 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8129__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8820__A _8820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7888__A1 _7881_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7888__B2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8837__B1 _4662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _7847_/A vssd1 vssd1 vccd1 vccd1 _6081_/S sky130_fd_sc_hd__buf_8
XANTENNA__5115__A2 _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6994__B _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6486__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6863__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7171__A _7171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8065__B2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7812__A1 _7809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7812__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8960_ _8979_/CLK hold9/X fanout732/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfrtp_1
X_7911_ _7918_/A1 _4947_/B _7918_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _7911_/Y sky130_fd_sc_hd__o22ai_2
X_8891_ _4824_/B _8890_/X _8888_/Y vssd1 vssd1 vccd1 vccd1 _8892_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7842_ _8150_/A _7858_/B vssd1 vssd1 vccd1 vccd1 _7842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6234__B _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7773_ _8716_/A _8516_/B vssd1 vssd1 vccd1 vccd1 _7872_/A sky130_fd_sc_hd__nor2_8
X_4985_ _8140_/A vssd1 vssd1 vccd1 vccd1 _6470_/B sky130_fd_sc_hd__buf_8
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6724_ _6724_/A _6724_/B vssd1 vssd1 vccd1 vccd1 _6724_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7879__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6655_ _7110_/A _6475_/X _6654_/X _6851_/B vssd1 vssd1 vccd1 vccd1 _6655_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6000__B1 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5606_ _5606_/A _6081_/S vssd1 vssd1 vccd1 vccd1 _5607_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6586_ _6906_/A _5241_/X _6585_/Y vssd1 vssd1 vccd1 vccd1 _6587_/A sky130_fd_sc_hd__o21ai_1
X_8325_ _8564_/B _7878_/Y _8349_/A vssd1 vssd1 vccd1 vccd1 _8325_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5537_ _5537_/A _6081_/S vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_103_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8256_ _8256_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _8259_/A sky130_fd_sc_hd__nand2_2
X_5468_ _5510_/A _4868_/A _5511_/A _5089_/A _5467_/X vssd1 vssd1 vccd1 vccd1 _6679_/B
+ sky130_fd_sc_hd__o221a_4
Xoutput640 _6360_/X vssd1 vssd1 vccd1 vccd1 sports_o[224] sky130_fd_sc_hd__buf_12
XANTENNA__7500__B1 _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput651 _7165_/X vssd1 vssd1 vccd1 vccd1 sports_o[29] sky130_fd_sc_hd__buf_12
Xoutput662 _7213_/X vssd1 vssd1 vccd1 vccd1 sports_o[39] sky130_fd_sc_hd__buf_12
X_7207_ _7206_/X _6058_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7208_/A sky130_fd_sc_hd__mux2_2
Xoutput673 _7260_/X vssd1 vssd1 vccd1 vccd1 sports_o[49] sky130_fd_sc_hd__buf_12
X_4419_ _4456_/B _4455_/B vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__nand2_1
Xoutput684 _6466_/X vssd1 vssd1 vccd1 vccd1 sports_o[59] sky130_fd_sc_hd__buf_12
X_8187_ _8189_/C _6456_/B _8196_/B1 _6495_/B _8186_/X vssd1 vssd1 vccd1 vccd1 _8187_/X
+ sky130_fd_sc_hd__o221a_4
X_5399_ _5031_/X _6611_/A _5397_/X _5398_/X vssd1 vssd1 vccd1 vccd1 _5399_/X sky130_fd_sc_hd__a22o_1
Xoutput695 _6600_/X vssd1 vssd1 vccd1 vccd1 sports_o[69] sky130_fd_sc_hd__buf_12
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8056__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7138_ _7138_/A vssd1 vssd1 vccd1 vccd1 _7138_/X sky130_fd_sc_hd__buf_8
XANTENNA__6067__B1 _6057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7803__A1 _4566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6606__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7803__B2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7069_ _7069_/A vssd1 vssd1 vccd1 vccd1 _7069_/X sky130_fd_sc_hd__buf_1
XFILLER_0_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6425__A _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8764__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5593__A2 _5635_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6790__B2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 mports_i[116] vssd1 vssd1 vccd1 vccd1 _4977_/B sky130_fd_sc_hd__buf_2
XANTENNA__8531__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7256__A _7256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4599__B _7309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8819__B1 _8190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5504__A _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8047__A1 _8054_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8047__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5281__A1 _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5569__C1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5033__A1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5033__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8550__A _8550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _4770_/A _4770_/B _4770_/C vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__nand3_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6989__B _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8507__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5893__B _5893_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8522__A2 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6440_ _6440_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _6443_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6533__A1 _5159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6533__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6371_ _6284_/A _7743_/A _6261_/A vssd1 vssd1 vccd1 vccd1 _6371_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8110_ _8110_/A vssd1 vssd1 vccd1 vccd1 _8110_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_140_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8286__A1 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5322_ _6609_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _5322_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8709__B _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8041_ _7874_/X _8030_/Y _7875_/X _8031_/Y vssd1 vssd1 vccd1 vccd1 _8041_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6836__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5253_ _5218_/A _7299_/A _6281_/S _6578_/B vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8038__B2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5184_ _6544_/A _5682_/B _6526_/A _8188_/S vssd1 vssd1 vccd1 vccd1 _5184_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6049__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7797__B1 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7261__A2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8943_ _8942_/A _4553_/B hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8874_ _8893_/A _8874_/B vssd1 vssd1 vccd1 vccd1 _8886_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_94_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8210__A1 _8210_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7825_ _7827_/A _5780_/X _7836_/A _5079_/X _7824_/X vssd1 vssd1 vccd1 vccd1 _7825_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8210__B2 _5106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7756_ _7756_/A _7756_/B vssd1 vssd1 vccd1 vccd1 _7756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _4968_/A vssd1 vssd1 vccd1 vccd1 _4968_/X sky130_fd_sc_hd__buf_1
XANTENNA__6772__A1 _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6899__B _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6707_ _5552_/X _6549_/A _5554_/X _6876_/C vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7687_ _6156_/Y _7680_/B _7685_/X _7640_/B _7686_/Y vssd1 vssd1 vccd1 vccd1 _7687_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4899_ _4899_/A vssd1 vssd1 vccd1 vccd1 _4899_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6638_ _6635_/Y _6925_/B _6637_/Y _6882_/B _7001_/S vssd1 vssd1 vccd1 vccd1 _6638_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6569_ _6628_/B _6569_/B vssd1 vssd1 vccd1 vccd1 _6569_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8277__A1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8308_ _7786_/X hold26/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8308_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8239_ _8239_/A vssd1 vssd1 vccd1 vccd1 _8239_/Y sky130_fd_sc_hd__inv_2
Xoutput470 _8602_/X vssd1 vssd1 vccd1 vccd1 mports_o[71] sky130_fd_sc_hd__buf_12
XFILLER_0_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput481 _8636_/X vssd1 vssd1 vccd1 vccd1 mports_o[81] sky130_fd_sc_hd__buf_12
Xoutput492 _8670_/X vssd1 vssd1 vccd1 vccd1 mports_o[91] sky130_fd_sc_hd__buf_12
XANTENNA__7237__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7788__B1 _7790_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7252__A2 _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__B1_N _5153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5263__A1 _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8201__A1 _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__A1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8752__A2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6763__A1 _5744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6763__B2 _5770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4403__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7712__B1 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6279__B1 _6314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output444_A _8399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7228__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output611_A _5779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7779__B1 _7779_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7243__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8264__B _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5254__A1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6451__B1 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5940_ _8160_/A _6231_/C _6839_/B vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__or3_1
XANTENNA__8728__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5871_ _5871_/A vssd1 vssd1 vccd1 vccd1 _5871_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5006__B2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8743__A2 _7878_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7610_ _7610_/A _7619_/B vssd1 vssd1 vccd1 vccd1 _7610_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4822_ _4607_/A _4748_/B _4793_/Y _4821_/Y _4758_/A vssd1 vssd1 vccd1 vccd1 _8887_/B
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5557__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8590_ _8590_/A vssd1 vssd1 vccd1 vccd1 _8590_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__6754__A1 _5744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6754__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7541_ _7153_/A _7668_/B _5711_/X _7638_/B vssd1 vssd1 vccd1 vccd1 _7541_/X sky130_fd_sc_hd__a22o_1
X_4753_ _5089_/A vssd1 vssd1 vccd1 vccd1 _8256_/A sky130_fd_sc_hd__inv_2
XFILLER_0_145_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5409__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7472_ _7466_/X _7471_/X _5464_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7472_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4684_ _4684_/A _4684_/B vssd1 vssd1 vccd1 vccd1 _7272_/B sky130_fd_sc_hd__nand2_4
XANTENNA__6231__C _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6423_ _6434_/B _7372_/B vssd1 vssd1 vccd1 vccd1 _6510_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6354_ _6357_/A1 _8716_/B input75/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6354_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8439__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5305_ _6593_/A vssd1 vssd1 vccd1 vccd1 _6875_/B sky130_fd_sc_hd__buf_8
XFILLER_0_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6285_ _5128_/A _6272_/X _6282_/X _6133_/B _6284_/Y vssd1 vssd1 vccd1 vccd1 _6285_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5144__A _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8024_ _8024_/A1 _7876_/X _8024_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _8024_/Y sky130_fd_sc_hd__o22ai_2
Xinput209 mports_i[82] vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__buf_2
X_5236_ _5265_/A _4931_/A _5266_/A _5111_/A _5235_/X vssd1 vssd1 vccd1 vccd1 _5239_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5493__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5167_ _8444_/A input12/X _5130_/A _5222_/B1 vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__a22o_1
XANTENNA__8455__A _8455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5798__B _6211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5098_ _6356_/S vssd1 vssd1 vccd1 vccd1 _6386_/S sky130_fd_sc_hd__buf_8
XANTENNA__5245__A1 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5245__B2 _5356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8926_ _8850_/B hold44/X _8926_/S vssd1 vssd1 vccd1 vccd1 _8927_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8857_ _8857_/A _8857_/B vssd1 vssd1 vccd1 vccd1 _8857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8195__B1 hold44/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7808_ _6080_/A _7813_/A2 _6513_/A _7813_/B2 vssd1 vssd1 vccd1 vccd1 _7808_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5548__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8788_ _8787_/X _8055_/Y _8788_/S vssd1 vssd1 vccd1 vccd1 _8788_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6745__A1 _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7739_ _6349_/X _7753_/B _7278_/A _7349_/A _7715_/S vssd1 vssd1 vccd1 vccd1 _7739_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5705__C1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5181__B1 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5720__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4877__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5054__A _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8670__A1 _8499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7473__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5989__A _5989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4893__A _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8422__A1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7225__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5236__B2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6433__B1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5787__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__B1 _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6613__A _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6717__A1_N _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8489__A1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6913_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _6116_/B sky130_fd_sc_hd__nand2_1
XANTENNA__8661__A1 _8483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7464__A2 _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8661__B2 _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5475__A1 _5661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5899__A _5899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5475__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _6281_/S vssd1 vssd1 vccd1 vccd1 _8188_/S sky130_fd_sc_hd__buf_8
XANTENNA__5227__A1 _5248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6507__B _6507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5227__B2 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6972_ _6317_/X _6989_/B _6971_/X _6994_/B _7000_/S vssd1 vssd1 vccd1 vccd1 _6972_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8711_ _8711_/A vssd1 vssd1 vccd1 vccd1 _8711_/X sky130_fd_sc_hd__buf_4
XFILLER_0_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5923_ _5923_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _5923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8642_ _8641_/X _8400_/A _8690_/S vssd1 vssd1 vccd1 vccd1 _8643_/A sky130_fd_sc_hd__mux2_1
X_5854_ _5827_/A _5077_/A _6017_/A _5879_/A vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_146_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7924__B1 _7931_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4805_ _4813_/B _4805_/B _4813_/C vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8573_ _8573_/A vssd1 vssd1 vccd1 vccd1 _8573_/X sky130_fd_sc_hd__buf_1
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5785_ _7629_/B _6837_/A _6780_/B _5784_/X _5013_/Y vssd1 vssd1 vccd1 vccd1 _5785_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5139__A _5139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7524_ _7524_/A _7660_/B vssd1 vssd1 vccd1 vccd1 _7524_/X sky130_fd_sc_hd__and2_1
XFILLER_0_133_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4736_ _4736_/A _4736_/B vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7455_ _7449_/Y _7454_/X _6630_/A _7741_/S vssd1 vssd1 vccd1 vccd1 _7455_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4978__A hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4667_ _4693_/B hold39/A vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6406_ _6500_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5163__B1 _5161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7386_ _7383_/Y _7297_/B _7575_/A _7385_/Y vssd1 vssd1 vccd1 vccd1 _7386_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_102_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4598_ _4607_/A _8174_/A _4607_/B _4596_/B vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6337_ input10/X _4913_/X _6337_/B1 _8516_/B _6336_/X vssd1 vssd1 vccd1 vccd1 _6337_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__8652__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6268_ _6258_/X _6261_/X _6267_/Y _6224_/S _6263_/X vssd1 vssd1 vccd1 vccd1 _6268_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__8968__RESET_B input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8007_ _8002_/Y _6080_/A _8003_/Y _6513_/A _8006_/Y vssd1 vssd1 vccd1 vccd1 _8416_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__6663__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5219_ _6233_/B _5219_/B vssd1 vssd1 vccd1 vccd1 _5219_/Y sky130_fd_sc_hd__nor2_1
X_6199_ _7767_/A _7829_/A _6231_/C _6931_/A vssd1 vssd1 vccd1 vccd1 _6199_/X sky130_fd_sc_hd__or4_1
XANTENNA__6417__B _7309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5769__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6966__B2 _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8909_ _8874_/B hold30/X _8909_/S vssd1 vssd1 vccd1 vccd1 _8910_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8168__B1 _8162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7529__A _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6718__A1 _7524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7915__B1 _7918_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6718__B2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6194__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6152__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7391__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7679__C1 _7334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8340__B1 _7912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8891__A1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8794__S _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5457__A1 _5401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5457__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7203__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5209__A1 _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output407_A _7988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7439__A _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ _5031_/X _5548_/X _5556_/X _5569_/X vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_25_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4521_ _4521_/A _4521_/B vssd1 vssd1 vccd1 vccd1 _4596_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7134__A1 _5552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8331__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7134__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7240_ _7240_/A vssd1 vssd1 vccd1 vccd1 _7240_/X sky130_fd_sc_hd__buf_1
XANTENNA__8882__A1 _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4452_ _8166_/A vssd1 vssd1 vccd1 vccd1 _7852_/A sky130_fd_sc_hd__inv_6
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold44_A hold44/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7171_ _7171_/A vssd1 vssd1 vccd1 vccd1 _7172_/A sky130_fd_sc_hd__inv_2
XFILLER_0_22_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4383_ hold32/X _8709_/A vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6122_ _6122_/A _7829_/A vssd1 vssd1 vccd1 vccd1 _6122_/Y sky130_fd_sc_hd__nand2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8634__A1 _7972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7437__A2 _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5448__A1 _6634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5448__B2 _6648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A vssd1 vssd1 vccd1 vccd1 _6053_/Y sky130_fd_sc_hd__inv_2
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7113__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5422__A _6634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5004_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5004_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8398__B1 _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6952__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7070__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6852_/A _6257_/A _6899_/B vssd1 vssd1 vccd1 vccd1 _6955_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7349__A _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5906_ _6470_/B _5875_/Y _5905_/Y vssd1 vssd1 vccd1 vccd1 _6807_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6886_ _6886_/A _6940_/A vssd1 vssd1 vccd1 vccd1 _6886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8625_ _8698_/B _8366_/X _8590_/X vssd1 vssd1 vccd1 vccd1 _8625_/X sky130_fd_sc_hd__o21a_1
X_5837_ _5881_/A1 _4871_/A input52/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8570__B1 _8249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8556_ _4940_/X _8157_/X _4933_/X _8200_/X _8555_/Y vssd1 vssd1 vccd1 vccd1 _8556_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_106_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5768_ _6744_/A vssd1 vssd1 vccd1 vccd1 _6906_/A sky130_fd_sc_hd__buf_4
XFILLER_0_44_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7507_ _7507_/A _7507_/B vssd1 vssd1 vccd1 vccd1 _7507_/Y sky130_fd_sc_hd__nor2_1
X_4719_ _5274_/A _4719_/B vssd1 vssd1 vccd1 vccd1 _4720_/A sky130_fd_sc_hd__nand2_1
X_8487_ _8299_/X _8482_/Y _8486_/Y _8304_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8487_/X
+ sky130_fd_sc_hd__a221o_1
X_5699_ _5718_/A1 _8271_/B input47/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5699_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7438_ _7094_/Y _7630_/B _5391_/Y _8755_/C vssd1 vssd1 vccd1 vccd1 _7438_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5687__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7369_ _6553_/A _7361_/X _7367_/X _7326_/A _7368_/Y vssd1 vssd1 vccd1 vccd1 _7369_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8625__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6636__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7531__B _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7833__C1 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6428__A _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6100__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6939__A1 _7696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7600__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8010__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7116__A1 _6671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8313__B1 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__A _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5678__B2 _5628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8092__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5242__A _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7052__A0 _7051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5063__C1 _5062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6595__A1_N _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6740_ _6738_/X _6899_/B _7000_/S _6739_/X vssd1 vssd1 vccd1 vccd1 _6740_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6671_ _6841_/A _6671_/B vssd1 vssd1 vccd1 vccd1 _6671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_128_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8552__B1 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8410_ _8564_/B _7999_/Y _8497_/S vssd1 vssd1 vccd1 vccd1 _8410_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5622_ _5618_/X _6233_/B _6170_/A _5621_/X vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6801__A _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8341_ _8339_/X _8340_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8342_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7107__A1 _7459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5553_ _6697_/B _7299_/A _6281_/S _5552_/X vssd1 vssd1 vccd1 vccd1 _5553_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7108__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4504_ _4504_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4505_/A sky130_fd_sc_hd__nand2_1
X_8272_ _8272_/A _8336_/S vssd1 vssd1 vccd1 vccd1 _8316_/A sky130_fd_sc_hd__nand2_1
X_5484_ _7474_/B _5707_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7223_ _6115_/A _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7223_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6866__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4435_ _4420_/Y _4430_/Y _8913_/A vssd1 vssd1 vccd1 vccd1 _4436_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__6330__A2 _7729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7632__A _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7154_ _5738_/C _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7154_/X sky130_fd_sc_hd__a21o_1
X_4366_ _4696_/B _4823_/B vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6618__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6105_ _6047_/A _8335_/B _6048_/A _4913_/A _6104_/X vssd1 vssd1 vccd1 vccd1 _6112_/B
+ sky130_fd_sc_hd__o221a_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8083__A2 _8476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _5356_/B _7026_/X _7083_/X _7084_/X vssd1 vssd1 vccd1 vccd1 _7085_/X sky130_fd_sc_hd__o22a_1
X_4297_ _6434_/B vssd1 vssd1 vccd1 vccd1 _4416_/B sky130_fd_sc_hd__inv_2
XANTENNA__6094__A1 _6047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6094__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6061_/A1 _8368_/A input59/X _4940_/A vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__o22a_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6397__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _7777_/X _8772_/B _7792_/X vssd1 vssd1 vccd1 vccd1 _7987_/X sky130_fd_sc_hd__o21ba_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7594__A1 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _6221_/Y _6989_/B _6937_/X _6994_/B _6946_/S vssd1 vssd1 vccd1 vccd1 _6938_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6869_ _6867_/Y _6868_/Y _8150_/A vssd1 vssd1 vccd1 vccd1 _6869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8608_ _8607_/X _7862_/Y _8686_/B vssd1 vssd1 vccd1 vccd1 _8609_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6554__C1 _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8539_ _8564_/B _8538_/X _8349_/A vssd1 vssd1 vccd1 vccd1 _8539_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7649__A2 _6074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6857__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7542__A _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6158__A _6158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8074__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6085__A1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__A _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7282__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6085__B2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6388__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7585__A1 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7337__A1 _5028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8820__B _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7888__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7436__B _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6340__B _6375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4571__A1 _5106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8837__B2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5520__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8065__A2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7273__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7812__A2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5823__A1 _5825_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5823__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7910_ _7910_/A vssd1 vssd1 vccd1 vccd1 _7910_/Y sky130_fd_sc_hd__inv_2
X_8890_ _4661_/A _4578_/Y _8264_/A _8759_/A vssd1 vssd1 vccd1 vccd1 _8890_/X sky130_fd_sc_hd__a31o_1
X_7841_ _7841_/A vssd1 vssd1 vccd1 vccd1 _7841_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7576__A1 _5827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7576__B2 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7772_ _7826_/A vssd1 vssd1 vccd1 vccd1 _7772_/X sky130_fd_sc_hd__clkbuf_8
X_4984_ _8160_/A vssd1 vssd1 vccd1 vccd1 _8140_/A sky130_fd_sc_hd__buf_6
XFILLER_0_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6723_ _6719_/X _6450_/X _6720_/Y _6721_/Y _6722_/X vssd1 vssd1 vccd1 vccd1 _6723_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5339__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7879__A2 _7878_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6654_ _5487_/A _6780_/A _5426_/Y vssd1 vssd1 vccd1 vccd1 _6654_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5605_ _6024_/A _5658_/A vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6585_ _6585_/A _6906_/A vssd1 vssd1 vccd1 vccd1 _6585_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8324_ _7869_/Y _8304_/X _7871_/Y _8299_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8324_/X
+ sky130_fd_sc_hd__a221o_1
X_5536_ _6133_/B _5535_/X _6284_/A _6679_/B vssd1 vssd1 vccd1 vccd1 _5536_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__8828__A1 _8222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8255_ _8584_/A _8222_/X _8295_/A _8261_/A vssd1 vssd1 vccd1 vccd1 _8255_/X sky130_fd_sc_hd__a22o_1
X_5467_ _5543_/A1 _4871_/A input39/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5467_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_112_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8458__A _8458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput630 _6225_/X vssd1 vssd1 vccd1 vccd1 sports_o[215] sky130_fd_sc_hd__buf_12
XFILLER_0_112_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput641 _6376_/X vssd1 vssd1 vccd1 vccd1 sports_o[225] sky130_fd_sc_hd__buf_12
XFILLER_0_111_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7362__A _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput652 _7031_/X vssd1 vssd1 vccd1 vccd1 sports_o[2] sky130_fd_sc_hd__buf_12
X_7206_ _6063_/A _7026_/X _7205_/X vssd1 vssd1 vccd1 vccd1 _7206_/X sky130_fd_sc_hd__o21a_1
Xoutput663 _7036_/X vssd1 vssd1 vccd1 vccd1 sports_o[3] sky130_fd_sc_hd__buf_12
X_4418_ _4515_/A _4601_/B _4515_/B vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__nand3_1
Xoutput674 _7042_/X vssd1 vssd1 vccd1 vccd1 sports_o[4] sky130_fd_sc_hd__buf_12
X_8186_ _6470_/B _8192_/A _8185_/Y vssd1 vssd1 vccd1 vccd1 _8186_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_111_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5398_ _6202_/B _5317_/A _5136_/X vssd1 vssd1 vccd1 vccd1 _5398_/X sky130_fd_sc_hd__o21a_1
Xoutput685 _7048_/X vssd1 vssd1 vccd1 vccd1 sports_o[5] sky130_fd_sc_hd__buf_12
Xoutput696 _7053_/X vssd1 vssd1 vccd1 vccd1 sports_o[6] sky130_fd_sc_hd__buf_12
XANTENNA__8056__A2 _8055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7137_ _7137_/A vssd1 vssd1 vccd1 vccd1 _7137_/X sky130_fd_sc_hd__buf_1
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4349_ _4349_/A vssd1 vssd1 vccd1 vccd1 _8512_/S sky130_fd_sc_hd__buf_8
XANTENNA__8461__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7803__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7068_ _7067_/X _5211_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__mux2_1
X_6019_ _6072_/A _5982_/A _6481_/B vssd1 vssd1 vccd1 vccd1 _7637_/B sky130_fd_sc_hd__mux2_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5290__A2 _5239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__B _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6441__A _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8819__A1 _8187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8819__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4896__A _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8368__A _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4305__A1 _5827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8047__A2 _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5281__A2 _5333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5569__B1 _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5033__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6230__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8550__B _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6781__A2 _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7447__A _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6070__B _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8966__CLK _8967_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6533__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6370_ _6349_/X _5682_/B _8188_/S _7743_/A vssd1 vssd1 vccd1 vccd1 _6370_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_125_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5321_ _6870_/S _5227_/X _7424_/A vssd1 vssd1 vccd1 vccd1 _6609_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__6297__A1 _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7182__A _7182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6297__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8040_ _8036_/Y _7954_/X _8468_/A _7826_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _8040_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7494__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5252_ _6793_/S vssd1 vssd1 vccd1 vccd1 _6593_/A sky130_fd_sc_hd__buf_8
XFILLER_0_139_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8038__A2 _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5183_ _5195_/A1 _4953_/X _5195_/B1 _4870_/A _5182_/X vssd1 vssd1 vccd1 vccd1 _6526_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6049__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7797__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7797__B2 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4843__A1_N hold10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8942_ _8942_/A hold12/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__nand2_1
XANTENNA__6526__A _6526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8873_ _8893_/B vssd1 vssd1 vccd1 vccd1 _8874_/B sky130_fd_sc_hd__inv_2
XFILLER_0_64_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8210__A2 _6102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7824_ _7823_/Y _4474_/Y hold23/A vssd1 vssd1 vccd1 vccd1 _7824_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_148_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7755_ _7752_/Y _7754_/A _7753_/Y _7754_/Y vssd1 vssd1 vccd1 vccd1 _7755_/X sky130_fd_sc_hd__a31o_1
X_4967_ _4964_/X _4966_/X _6224_/S vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6261__A _6261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6706_ _5595_/Y _6475_/A _6705_/X _6694_/B vssd1 vssd1 vccd1 vccd1 _6706_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7686_ _7686_/A _7686_/B vssd1 vssd1 vccd1 vccd1 _7686_/Y sky130_fd_sc_hd__nor2_1
X_4898_ _4883_/Y _8550_/B _4888_/Y _4891_/X _4897_/Y vssd1 vssd1 vccd1 vccd1 _4899_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6637_ _6637_/A vssd1 vssd1 vccd1 vccd1 _6637_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6568_ _6535_/Y _6567_/Y _8924_/B vssd1 vssd1 vccd1 vccd1 _6568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _5519_/A vssd1 vssd1 vccd1 vccd1 _5519_/Y sky130_fd_sc_hd__inv_2
X_8307_ _8349_/A _8293_/X _8298_/Y _8306_/X vssd1 vssd1 vccd1 vccd1 _8307_/X sky130_fd_sc_hd__o22a_2
XFILLER_0_131_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6499_ _6499_/A vssd1 vssd1 vccd1 vccd1 _6543_/A sky130_fd_sc_hd__inv_2
XANTENNA__5605__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8238_ _4607_/A _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _8238_/Y sky130_fd_sc_hd__a21oi_1
Xoutput460 _8544_/X vssd1 vssd1 vccd1 vccd1 mports_o[62] sky130_fd_sc_hd__buf_12
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput471 _8605_/X vssd1 vssd1 vccd1 vccd1 mports_o[72] sky130_fd_sc_hd__buf_12
Xoutput482 _8639_/X vssd1 vssd1 vccd1 vccd1 mports_o[82] sky130_fd_sc_hd__buf_12
XANTENNA__5324__B _6181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput493 _8673_/X vssd1 vssd1 vccd1 vccd1 mports_o[92] sky130_fd_sc_hd__buf_12
X_8169_ _8169_/A vssd1 vssd1 vccd1 vccd1 _8169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7788__A1 _7790_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7788__B2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6436__A _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8201__A2 _8198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6870__S _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5486__S _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7960__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6763__A2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4403__B _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6515__A2 _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7712__A1 _7532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6279__A1 _6315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6279__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7779__B2 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output604_A _5570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__A2 _8709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6451__A1 _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8728__B1 _7800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5870_ _6079_/A _5930_/A vssd1 vssd1 vccd1 vccd1 _5870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5006__A2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4821_ _4821_/A _5191_/A vssd1 vssd1 vccd1 vccd1 _4821_/Y sky130_fd_sc_hd__nor2_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6754__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7951__B2 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7540_ _5654_/Y _7332_/A _7539_/X vssd1 vssd1 vccd1 vccd1 _7540_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4752_ _4752_/A _4752_/B vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5409__B _7094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7471_ _6667_/X _7673_/A _7749_/S _7469_/X _7470_/Y vssd1 vssd1 vccd1 vccd1 _7471_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4683_ _5129_/A _4719_/B vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7703__A1 _6234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6231__D _6944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7703__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6422_ _6416_/X _4919_/X _7000_/S vssd1 vssd1 vccd1 vccd1 _6422_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_141_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8500__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6353_ _6349_/X _6234_/B _7278_/A _5128_/A vssd1 vssd1 vccd1 vccd1 _6353_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5425__A _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5304_ _5909_/B _5280_/A _5303_/Y _5997_/B vssd1 vssd1 vccd1 vccd1 _5304_/X sky130_fd_sc_hd__a22o_1
X_6284_ _6284_/A _7251_/B vssd1 vssd1 vccd1 vccd1 _6284_/Y sky130_fd_sc_hd__nor2_1
X_8023_ _8427_/A _7954_/X _8423_/A _7826_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _8023_/X
+ sky130_fd_sc_hd__a221o_1
X_5235_ input92/X _4934_/A input29/X _4938_/A vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5493__A2 _7470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7219__B1 _7061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5166_ _5166_/A vssd1 vssd1 vccd1 vccd1 _7383_/A sky130_fd_sc_hd__inv_2
XANTENNA__4983__B _6456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8455__B _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8431__A2 _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5097_ _6084_/B vssd1 vssd1 vccd1 vccd1 _5845_/B sky130_fd_sc_hd__buf_8
XANTENNA__5245__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8925_ _8926_/S _8861_/A _8924_/Y vssd1 vssd1 vccd1 vccd1 _8958_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__8719__B1 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8856_ _8865_/A _8856_/B vssd1 vssd1 vccd1 vccd1 _8856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7807_ _7814_/A1 _5359_/B _7814_/B1 _7316_/A _7806_/X vssd1 vssd1 vccd1 vccd1 _7807_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _7620_/A _5999_/B vssd1 vssd1 vccd1 vccd1 _5999_/Y sky130_fd_sc_hd__nand2_1
X_8787_ _8458_/A _8711_/A _8506_/Y _8770_/B vssd1 vssd1 vccd1 vccd1 _8787_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7942__B2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5953__B1 _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7738_ _7736_/Y _7332_/A _7737_/Y vssd1 vssd1 vccd1 vccd1 _7738_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7669_ _7668_/Y _7297_/B _7694_/A _7385_/Y vssd1 vssd1 vccd1 vccd1 _7669_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4508__A1 _8240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5705__B1 _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6902__C1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5181__A1 _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5181__B2 _5218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5335__A _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6130__B1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8670__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5070__A _5070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5236__A2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4995__A1 _4975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__B2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8186__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7933__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6736__A2 _7544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7933__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7725__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7444__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output721_A _6850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6121__B1 _6140_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8661__A2 _8581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5475__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _6017_/A vssd1 vssd1 vccd1 vccd1 _6281_/S sky130_fd_sc_hd__buf_8
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5899__B _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5227__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7621__B1 _7385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6971_ _6971_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _6971_/X sky130_fd_sc_hd__and2_1
XFILLER_0_45_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8710_ _8712_/A vssd1 vssd1 vccd1 vccd1 _8711_/A sky130_fd_sc_hd__buf_4
X_5922_ _5931_/A _4929_/A _5932_/A _4932_/A _5921_/X vssd1 vssd1 vccd1 vccd1 _5923_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__8291__A _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8177__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5853_ _5804_/A _4929_/A _5805_/A _4932_/A _5852_/X vssd1 vssd1 vccd1 vccd1 _5853_/X
+ sky130_fd_sc_hd__o221a_4
X_8641_ _8640_/X _7999_/Y _8689_/S vssd1 vssd1 vccd1 vccd1 _8641_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7619__B _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7924__A1 _7931_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4804_ _4801_/Y _4802_/Y _4803_/Y vssd1 vssd1 vccd1 vccd1 _4813_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8572_ _8571_/X _8244_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8573_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5784_ _5999_/B _7560_/A _5782_/Y _7266_/B vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4735_ _4770_/A _4750_/C _4770_/C vssd1 vssd1 vccd1 vccd1 _4738_/A sky130_fd_sc_hd__nand3_1
X_7523_ _5600_/Y _7630_/B _5667_/Y _8755_/C vssd1 vssd1 vccd1 vccd1 _7523_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7454_ _6635_/Y _7681_/A _6643_/X _7673_/A _7453_/X vssd1 vssd1 vccd1 vccd1 _7454_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__7688__B1 _6212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4666_ _8880_/A hold7/X vssd1 vssd1 vccd1 vccd1 _8909_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4978__B _4978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6405_ _6549_/A vssd1 vssd1 vccd1 vccd1 _6462_/A sky130_fd_sc_hd__inv_2
XANTENNA__5163__A1 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5163__B2 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7385_ _7497_/B vssd1 vssd1 vccd1 vccd1 _7385_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4597_ _4597_/A vssd1 vssd1 vccd1 vccd1 _8174_/A sky130_fd_sc_hd__buf_12
XFILLER_0_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6336_ _6336_/A1 _8716_/B input73/X _4917_/X vssd1 vssd1 vccd1 vccd1 _6336_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8637__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8101__A1 _8106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6267_ _6267_/A _6375_/B vssd1 vssd1 vccd1 vccd1 _6267_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8652__A2 _8042_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7370__A _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6663__A1 _7470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8006_ _8011_/A1 _5146_/A _8011_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _8006_/Y sky130_fd_sc_hd__o22ai_2
X_5218_ _5218_/A vssd1 vssd1 vccd1 vccd1 _5219_/B sky130_fd_sc_hd__inv_2
XANTENNA__7860__B1 hold44/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6198_ _7680_/A _6197_/X _6593_/A vssd1 vssd1 vccd1 vccd1 _7694_/B sky130_fd_sc_hd__mux2_1
XANTENNA__8185__B _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5149_ _6261_/A vssd1 vssd1 vccd1 vccd1 _6128_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7612__B1 _7385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6966__A2 _6475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8908_ _8908_/A vssd1 vssd1 vccd1 vccd1 _8948_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__8405__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8168__A1 _8175_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8168__B2 _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8839_ _8833_/B _8252_/X _8725_/A vssd1 vssd1 vccd1 vccd1 _8839_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7915__A1 _7918_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6718__A2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7915__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7391__A2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7679__B1 _7347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8340__A1 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5154__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6351__B1 _6357_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5065__A _6359_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8376__A _8376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5457__A2 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7603__B1 _7334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8800__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6957__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6709__A2 _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7906__B2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5393__A1 _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520_ _4520_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _4521_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8331__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7134__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4451_ _8950_/Q vssd1 vssd1 vccd1 vccd1 _8166_/A sky130_fd_sc_hd__buf_8
XFILLER_0_123_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8882__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6893__A1 _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7170_ _7170_/A vssd1 vssd1 vccd1 vccd1 _7170_/X sky130_fd_sc_hd__buf_1
XFILLER_0_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4382_ _8977_/Q vssd1 vssd1 vccd1 vccd1 _8709_/A sky130_fd_sc_hd__inv_4
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6121_ input63/X _4896_/A _6140_/A1 _4893_/A _6120_/X vssd1 vssd1 vccd1 vccd1 _7678_/B
+ sky130_fd_sc_hd__a221oi_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5448__A2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6052_ _6081_/S _6080_/A _6897_/A _7650_/B vssd1 vssd1 vccd1 vccd1 _6053_/A sky130_fd_sc_hd__o31a_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5003_ _5003_/A vssd1 vssd1 vccd1 vccd1 _5003_/Y sky130_fd_sc_hd__inv_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5422__B _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8398__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7070__A1 _5218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4959__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6954_ _6954_/A vssd1 vssd1 vccd1 vccd1 _6954_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5905_ _5905_/A vssd1 vssd1 vccd1 vccd1 _5905_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6885_ _6941_/A _6060_/Y _8574_/B vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8624_ _7929_/Y _8583_/X _8362_/X _8581_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8624_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5836_ _5871_/A _4953_/A _5872_/A _5089_/A _5835_/X vssd1 vssd1 vccd1 vccd1 _6811_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8570__A1 _8247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8570__B2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8555_ _8555_/A _8555_/B vssd1 vssd1 vccd1 vccd1 _8555_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5767_ _6926_/A vssd1 vssd1 vccd1 vccd1 _6744_/A sky130_fd_sc_hd__inv_2
XFILLER_0_133_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7506_ _7754_/A _5634_/B _7330_/A vssd1 vssd1 vccd1 vccd1 _7506_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4718_ _8300_/B vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__inv_6
X_5698_ _5661_/A _8335_/B _5662_/A _4913_/A _5697_/X vssd1 vssd1 vccd1 vccd1 _6732_/A
+ sky130_fd_sc_hd__o221a_4
X_8486_ _8486_/A vssd1 vssd1 vccd1 vccd1 _8486_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4649_ _4946_/A vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__inv_8
X_7437_ _6611_/A _7741_/S _7430_/X _7436_/Y vssd1 vssd1 vccd1 vccd1 _7437_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_102_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5687__A2 _5718_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6884__A1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7368_ _7681_/A _7368_/B vssd1 vssd1 vccd1 vccd1 _7368_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8086__B1 _8093_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6319_ input10/X _4870_/X _6337_/B1 _8480_/B _6318_/X vssd1 vssd1 vccd1 vccd1 _7266_/A
+ sky130_fd_sc_hd__o221a_2
XANTENNA__8625__A2 _8366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7299_ _7299_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _7575_/A sky130_fd_sc_hd__nand2_8
XANTENNA__6636__A1 _6622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5613__A _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7833__B1 _7832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6636__B2 _6635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8389__A1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5072__B1 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8010__B1 _8009_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8561__A1 _8215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4899__A _4899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5375__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5375__B2 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8313__A1 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7116__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8313__B2 _7811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6324__B1 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8864__A2 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4411__B _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7824__B1 hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output517_A _7002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput360 sports_i[95] vssd1 vssd1 vccd1 vccd1 _8158_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5669__S _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7052__A1 _7352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6670_ _6432_/X _6669_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6670_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__8552__A1 _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8552__B2 _8203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5621_ _5845_/B _5552_/X _5620_/X _6133_/B vssd1 vssd1 vccd1 vccd1 _5621_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_144_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5366__A1 _5337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5366__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6801__B _6801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5552_ _5591_/A _4953_/X _5592_/A _5089_/X _5551_/X vssd1 vssd1 vccd1 vccd1 _5552_/X
+ sky130_fd_sc_hd__o221a_4
X_8340_ _4940_/X _7886_/Y _7912_/Y vssd1 vssd1 vccd1 vccd1 _8340_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7107__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4503_ _4514_/A _4503_/B _4525_/C vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__nand3_1
X_8271_ _8271_/A _8271_/B vssd1 vssd1 vccd1 vccd1 _8364_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5483_ _6593_/A _5674_/B _5482_/X vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7222_ _7222_/A vssd1 vssd1 vccd1 vccd1 _7222_/X sky130_fd_sc_hd__buf_1
X_4434_ _7384_/A hold10/X vssd1 vssd1 vccd1 vccd1 _8913_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7153_ _7153_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7153_/X sky130_fd_sc_hd__and2_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4365_ _8973_/Q vssd1 vssd1 vccd1 vccd1 _4696_/B sky130_fd_sc_hd__inv_2
XFILLER_0_111_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7124__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6104_ _6104_/A1 _8271_/B input61/X _4917_/A vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__o22a_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6618__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7815__B1 _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7084_ _7422_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7084_/X sky130_fd_sc_hd__a21o_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _8969_/Q vssd1 vssd1 vccd1 vccd1 _6434_/B sky130_fd_sc_hd__clkbuf_16
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6094__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6035_ _6035_/A vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__buf_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6963__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6264__A _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7986_ _7976_/Y _7875_/X _7977_/Y _7874_/X _7985_/Y vssd1 vssd1 vccd1 vccd1 _8772_/B
+ sky130_fd_sc_hd__a221oi_4
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7594__A2 _6811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _6937_/A _7266_/B vssd1 vssd1 vccd1 vccd1 _6937_/X sky130_fd_sc_hd__and2_1
XFILLER_0_138_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4801__B1 _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6868_ _6868_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6868_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7346__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5357__A1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8607_ _8315_/Y _8589_/A _8606_/X vssd1 vssd1 vccd1 vccd1 _8607_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5357__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5819_ _6234_/B _7568_/B _5816_/Y _5818_/Y vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6799_ _6870_/S _6772_/Y _6798_/Y vssd1 vssd1 vccd1 vccd1 _7577_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8538_ _8518_/A _8364_/A _8537_/X vssd1 vssd1 vccd1 vccd1 _8538_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8469_ _8469_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8469_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8919__A _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6857__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6857__B2 _6868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6439__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5343__A _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7806__B1 _5117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8952__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__B _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5997__B _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8231__B1 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7585__A2 _5879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8534__A1 _8157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6621__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5518__A _5518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4422__A _5145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8298__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7733__A _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5520__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5520__B2 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7273__A1 _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5823__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput190 mports_i[65] vssd1 vssd1 vccd1 vccd1 _5195_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__7025__A1 _4966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8222__B1 _8222_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6084__A _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7840_ _7840_/A vssd1 vssd1 vccd1 vccd1 _7840_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7576__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5587__A1 _5587_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5587__B2 _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7771_ _7779_/B1 _7769_/X _4476_/A _6500_/X _7770_/X vssd1 vssd1 vccd1 vccd1 _7771_/X
+ sky130_fd_sc_hd__a221o_4
X_4983_ _7027_/A _6456_/B vssd1 vssd1 vccd1 vccd1 _4986_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4316__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6722_ _5655_/A _6510_/A _5648_/Y _6512_/X vssd1 vssd1 vccd1 vccd1 _6722_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7328__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5339__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5339__B2 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6653_ _6653_/A vssd1 vssd1 vccd1 vccd1 _7110_/A sky130_fd_sc_hd__inv_2
XFILLER_0_128_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5604_ _5601_/Y _4885_/A _5602_/Y _4890_/A _5603_/Y vssd1 vssd1 vccd1 vccd1 _5658_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6584_ _6584_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8323_ _8572_/S vssd1 vssd1 vccd1 vccd1 _8323_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5535_ _7488_/A _5470_/Y _6547_/A vssd1 vssd1 vccd1 vccd1 _5535_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8254_ _7975_/A _8244_/X _8250_/X _8253_/X vssd1 vssd1 vccd1 vccd1 _8254_/X sky130_fd_sc_hd__a22o_2
X_5466_ _5466_/A vssd1 vssd1 vccd1 vccd1 _5466_/Y sky130_fd_sc_hd__inv_2
Xoutput620 _5987_/X vssd1 vssd1 vccd1 vccd1 sports_o[206] sky130_fd_sc_hd__buf_12
XANTENNA__4986__B _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput631 _6237_/Y vssd1 vssd1 vccd1 vccd1 sports_o[216] sky130_fd_sc_hd__buf_12
XFILLER_0_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8458__B _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput642 _6390_/Y vssd1 vssd1 vccd1 vccd1 sports_o[226] sky130_fd_sc_hd__buf_12
XFILLER_0_112_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4417_ _4417_/A hold40/A vssd1 vssd1 vccd1 vccd1 _4515_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7205_ _6016_/A _7004_/X _7639_/A _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7205_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput653 _7170_/X vssd1 vssd1 vccd1 vccd1 sports_o[30] sky130_fd_sc_hd__buf_12
Xoutput664 _7217_/X vssd1 vssd1 vccd1 vccd1 sports_o[40] sky130_fd_sc_hd__buf_12
X_8185_ _8185_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _8185_/Y sky130_fd_sc_hd__nand2_1
X_5397_ _6170_/A _5397_/B vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__or2_1
Xoutput675 _7265_/X vssd1 vssd1 vccd1 vccd1 sports_o[50] sky130_fd_sc_hd__buf_12
Xoutput686 _6479_/X vssd1 vssd1 vccd1 vccd1 sports_o[60] sky130_fd_sc_hd__buf_12
Xoutput697 _6605_/X vssd1 vssd1 vccd1 vccd1 sports_o[70] sky130_fd_sc_hd__buf_12
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7136_ _7135_/X _5644_/A _7175_/S vssd1 vssd1 vccd1 vccd1 _7137_/A sky130_fd_sc_hd__mux2_1
X_4348_ _4348_/A _4348_/B vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__and2_1
XANTENNA__7264__A1 _7729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6067__A2 _6058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7067_ _6551_/A _7023_/X _7066_/X vssd1 vssd1 vccd1 vccd1 _7067_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6693__S _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6018_ _8189_/A _6013_/Y _6017_/X vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5610__B _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4507__A _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__B1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8764__A1 _7956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7567__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5578__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7969_ _7962_/Y _7769_/X _7963_/Y _6500_/X _7968_/Y vssd1 vssd1 vccd1 vccd1 _7969_/Y
+ sky130_fd_sc_hd__a221oi_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6775__B1 _5803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7818__A _7818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8413__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8819__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7272__B _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4305__A2 _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7255__A1 _7720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6616__B _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8204__B1 _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5569__A1 _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6230__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8507__A1 _8104_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8507__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5248__A _5248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7730__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5320_ _5320_/A _6870_/S vssd1 vssd1 vccd1 vccd1 _7424_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5251_ _5265_/A _5089_/X _5266_/A _5080_/A _5250_/X vssd1 vssd1 vccd1 vccd1 _6578_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6297__A2 _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7494__A1 _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6079__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5182_ input88/X _5090_/A input26/X _4874_/A vssd1 vssd1 vccd1 vccd1 _5182_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6049__A2 _6104_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8294__A _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8443__B1 _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6807__A _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7797__A2 _7802_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5711__A _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8941_ _8941_/A vssd1 vssd1 vccd1 vccd1 _8978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8872_ _8872_/A _8872_/B vssd1 vssd1 vccd1 vccd1 _8893_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8746__A1 _8334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7823_ _7823_/A _8189_/A vssd1 vssd1 vccd1 vccd1 _7823_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6757__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7754_ _7754_/A _7754_/B vssd1 vssd1 vccd1 vccd1 _7754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4966_ _4956_/A _4930_/X _4957_/A _4933_/X _4965_/X vssd1 vssd1 vccd1 vccd1 _4966_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_19_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6705_ _5613_/B _5516_/B _6837_/A vssd1 vssd1 vccd1 vccd1 _6705_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6261__B _6261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7685_ _7364_/A _6167_/Y _6931_/Y _7630_/B vssd1 vssd1 vccd1 vccd1 _7685_/X sky130_fd_sc_hd__a2bb2o_1
X_4897_ _8713_/C input80/X _8579_/C input17/X vssd1 vssd1 vccd1 vccd1 _4897_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_129_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5158__A _5159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6636_ _6622_/A _5197_/X _8151_/B _6635_/A vssd1 vssd1 vccd1 vccd1 _6637_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7721__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5732__A1 _5792_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5732__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8469__A _8469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6567_ _6567_/A _6626_/B vssd1 vssd1 vccd1 vccd1 _6567_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7373__A _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8306_ _8306_/A _8564_/B vssd1 vssd1 vccd1 vccd1 _8306_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5518_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5518_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8131__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6498_ _6432_/X _6497_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6498_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__7485__A1 _5530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5605__B _5658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8682__B1 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8237_ _7975_/A _8226_/X _8233_/X _8236_/Y vssd1 vssd1 vccd1 vccd1 _8237_/X sky130_fd_sc_hd__a22o_2
X_5449_ _5497_/A1 _4871_/A input38/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5449_/X sky130_fd_sc_hd__o22a_1
Xoutput450 _8463_/X vssd1 vssd1 vccd1 vccd1 mports_o[53] sky130_fd_sc_hd__buf_12
Xoutput461 _8558_/X vssd1 vssd1 vccd1 vccd1 mports_o[63] sky130_fd_sc_hd__buf_12
XANTENNA__5496__B1 _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput472 _8609_/X vssd1 vssd1 vccd1 vccd1 mports_o[73] sky130_fd_sc_hd__buf_12
Xoutput483 _8643_/X vssd1 vssd1 vccd1 vccd1 mports_o[83] sky130_fd_sc_hd__buf_12
Xoutput494 _8677_/X vssd1 vssd1 vccd1 vccd1 mports_o[93] sky130_fd_sc_hd__buf_12
X_8168_ _8175_/A1 _6440_/B _8162_/A _4518_/A _8167_/X vssd1 vssd1 vccd1 vccd1 _8169_/A
+ sky130_fd_sc_hd__o221ai_2
XANTENNA__7237__A1 _6234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7119_ _7119_/A vssd1 vssd1 vccd1 vccd1 _7119_/X sky130_fd_sc_hd__buf_1
XANTENNA__7237__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8099_ _8106_/A1 _4947_/B _8106_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _8099_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__7788__A2 _7299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8737__A1 _7821_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6748__B1 _6449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5420__B1 _5402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7960__A2 _8765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7173__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6515__A3 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6920__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4700__A _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6279__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7228__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8318__S _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7779__A2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6451__A2 _4963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8728__A1 _7798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8728__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _8261_/A vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__inv_8
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7951__A2 _7013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7177__B _7246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5962__A1 _5962_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4751_ _4751_/A _4751_/B vssd1 vssd1 vccd1 vccd1 _4752_/B sky130_fd_sc_hd__and2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5962__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4682_ _4682_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4736_/A sky130_fd_sc_hd__nand2_1
X_7470_ _7470_/A _7696_/B vssd1 vssd1 vccd1 vccd1 _7470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7703__A2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6421_ _6946_/S vssd1 vssd1 vccd1 vccd1 _7000_/S sky130_fd_sc_hd__buf_6
XANTENNA__5714__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8289__A _8497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5714__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6352_ _6352_/A vssd1 vssd1 vccd1 vccd1 _7278_/A sky130_fd_sc_hd__inv_2
XFILLER_0_113_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5303_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5303_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5425__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6283_ _6283_/A vssd1 vssd1 vccd1 vccd1 _7251_/B sky130_fd_sc_hd__inv_2
XANTENNA__7467__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5478__B1 _5686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8022_ _8015_/Y _7769_/A _8016_/Y _6500_/A _8021_/Y vssd1 vssd1 vccd1 vccd1 _8423_/A
+ sky130_fd_sc_hd__a221oi_4
X_5234_ _5031_/X _6567_/A _5220_/X _5233_/X vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__a22o_2
XANTENNA__7640__B _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5165_ input90/X _4893_/A input27/X _4896_/A _5164_/X vssd1 vssd1 vccd1 vccd1 _5166_/A
+ sky130_fd_sc_hd__a221oi_2
XANTENNA__7132__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5441__A _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5096_ _5096_/A vssd1 vssd1 vccd1 vccd1 _6133_/B sky130_fd_sc_hd__buf_8
X_8924_ _8926_/S _8924_/B vssd1 vssd1 vccd1 vccd1 _8924_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8719__A1 _8297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8855_ _8855_/A _8861_/A vssd1 vssd1 vccd1 vccd1 _8865_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7368__A _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7806_ _7761_/A _7813_/A2 _5117_/A _7813_/B2 vssd1 vssd1 vccd1 vccd1 _7806_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8786_ _8494_/Y _8759_/Y _8785_/X _8725_/X vssd1 vssd1 vccd1 vccd1 _8786_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _6852_/B vssd1 vssd1 vccd1 vccd1 _7620_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7942__A2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7737_ _7756_/A _7737_/B vssd1 vssd1 vccd1 vccd1 _7737_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4949_ _4949_/A _6266_/A vssd1 vssd1 vccd1 vccd1 _6359_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_62_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7668_ _7668_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7668_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5705__A1 _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6619_ _7439_/B _6994_/B _6616_/Y _6618_/Y vssd1 vssd1 vccd1 vccd1 _6620_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6902__B1 _6528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7599_ _7701_/A _7599_/B vssd1 vssd1 vccd1 vccd1 _7599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5181__A2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5469__B1 _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6130__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6166__B _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6969__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__A2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8186__A2 _8192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7933__A2 _7932_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5944__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5944__B2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7146__A0 _7145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8343__C1 _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7697__A1 _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7725__B _7725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6121__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6121__B2 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6672__A2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6970_ _7725_/B _6429_/S _6968_/X _6969_/X vssd1 vssd1 vccd1 vccd1 _6970_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _6007_/A1 _4935_/A input57/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8177__A2 _8157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8640_ _8403_/A _8581_/A _8426_/Y _8583_/A vssd1 vssd1 vccd1 vccd1 _8640_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_48_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5852_ _5881_/A1 _4935_/A input52/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4803_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4803_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8571_ _8252_/X _8567_/B _8570_/X vssd1 vssd1 vccd1 vccd1 _8571_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_17_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5783_ _6756_/B vssd1 vssd1 vccd1 vccd1 _7560_/A sky130_fd_sc_hd__inv_2
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7522_ _7510_/B _5655_/A _7398_/A vssd1 vssd1 vccd1 vccd1 _7528_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_43_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4734_ _4734_/A _4734_/B vssd1 vssd1 vccd1 vccd1 _4770_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_44_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7453_ _7640_/B _7450_/Y _7451_/Y _7452_/Y vssd1 vssd1 vccd1 vccd1 _7453_/X sky130_fd_sc_hd__a31o_1
XANTENNA__7688__B2 _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4665_ hold18/X _8574_/B vssd1 vssd1 vccd1 vccd1 _8880_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5436__A _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6404_ _6434_/B _7297_/B vssd1 vssd1 vccd1 vccd1 _6549_/A sky130_fd_sc_hd__nor2_4
X_7384_ _7384_/A _7510_/B vssd1 vssd1 vccd1 vccd1 _7497_/B sky130_fd_sc_hd__nand2_2
X_4596_ _4596_/A _4596_/B vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6335_ _7266_/A _6084_/B _5128_/A _6333_/Y _6334_/Y vssd1 vssd1 vccd1 vccd1 _6335_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8637__B1 _7983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8101__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6266_ _6266_/A _7372_/B vssd1 vssd1 vccd1 vccd1 _6375_/B sky130_fd_sc_hd__nand2_4
X_8005_ _8002_/Y _7013_/A _8003_/Y _5116_/A _8004_/Y vssd1 vssd1 vccd1 vccd1 _8412_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6663__A2 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8979__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5217_ _5909_/B _7071_/A _6590_/B _5997_/B vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__a22o_1
X_6197_ _6149_/Y _6196_/Y _6281_/S vssd1 vssd1 vccd1 vccd1 _6197_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5171__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5148_ _5148_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _5148_/Y sky130_fd_sc_hd__nand2_1
X_5079_ _5079_/A vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__clkbuf_16
X_8907_ _8899_/A hold31/X _8909_/S vssd1 vssd1 vccd1 vccd1 _8908_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8168__A2 _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8838_ _8247_/Y _8711_/X _8249_/X _8803_/B _8788_/S vssd1 vssd1 vccd1 vccd1 _8838_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8977__RESET_B input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7915__A2 _5780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8769_ _8436_/Y _8759_/Y _8768_/X _8725_/X vssd1 vssd1 vccd1 vccd1 _8769_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7679__A1 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8340__A2 _7886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6351__A1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__A2 _7356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6351__B2 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8628__B1 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8376__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6654__A2 _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7603__A1 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8800__B1 _8104_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7906__A2 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5917__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8867__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5256__A _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8331__A2 _7906_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4450_ _4430_/Y _4449_/Y _4420_/Y vssd1 vssd1 vccd1 vccd1 _4525_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__8882__A3 _4662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4353__B1 _4674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _8967_/D sky130_fd_sc_hd__buf_2
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6120_ _8444_/A _6141_/A1 _8257_/C _6141_/B1 vssd1 vssd1 vccd1 vccd1 _6120_/X sky130_fd_sc_hd__a22o_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6051_/A _6081_/S vssd1 vssd1 vccd1 vccd1 _7650_/B sky130_fd_sc_hd__nand2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__A1 _5359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5853__B1 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__B2 _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _6080_/A vssd1 vssd1 vccd1 vccd1 _6965_/A sky130_fd_sc_hd__buf_12
XANTENNA__5422__C hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8398__A2 _8772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6815__A _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7070__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4959__A2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6953_ _6952_/X _6248_/X _7001_/S vssd1 vssd1 vccd1 vccd1 _6954_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5081__A1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6026__S _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5904_ _5904_/A _7829_/A vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6884_ _8574_/B _8857_/B _6060_/Y _6883_/X vssd1 vssd1 vccd1 vccd1 _6884_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8623_ _8623_/A vssd1 vssd1 vccd1 vccd1 _8623_/X sky130_fd_sc_hd__buf_1
XFILLER_0_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5835_ _5902_/A1 _4871_/A input53/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5835_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_119_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8570__A2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7646__A _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8554_ _8567_/B _8547_/Y _8553_/X vssd1 vssd1 vccd1 vccd1 _8554_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_17_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6550__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5766_ _5763_/X _5765_/X _6386_/S vssd1 vssd1 vccd1 vccd1 _5766_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_146_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7505_ _7749_/S _7505_/B vssd1 vssd1 vccd1 vccd1 _7505_/X sky130_fd_sc_hd__or2_1
XANTENNA__8858__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4717_ hold26/A hold41/A vssd1 vssd1 vccd1 vccd1 _8300_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_17_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8485_ _8484_/X _8428_/X _8755_/B vssd1 vssd1 vccd1 vccd1 _8486_/A sky130_fd_sc_hd__mux2_1
X_5697_ _5697_/A1 _8271_/B input46/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5697_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_115_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7436_ _7436_/A _7723_/B vssd1 vssd1 vccd1 vccd1 _7436_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4648_ _8958_/Q hold44/A vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6884__A2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7367_ _6573_/B _7680_/B _7365_/X _7348_/A _7366_/Y vssd1 vssd1 vccd1 vccd1 _7367_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4579_ _8336_/S vssd1 vssd1 vccd1 vccd1 _8904_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7381__A _7686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8086__A1 _8093_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6318_ _6336_/A1 _8310_/B input73/X _4874_/X vssd1 vssd1 vccd1 vccd1 _6318_/X sky130_fd_sc_hd__o22a_1
X_7298_ _7660_/B vssd1 vssd1 vccd1 vccd1 _7686_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__6097__B1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7833__A1 _7825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6636__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6249_ _6246_/X _6248_/X _6359_/S vssd1 vssd1 vccd1 vccd1 _6250_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7833__B2 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8924__B _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8389__A2 _8379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6725__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7597__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5072__A1 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5072__B2 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8010__A1 _8416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8010__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8561__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7556__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6460__A _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5375__A2 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6324__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5127__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6324__B2 _6317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7291__A _7291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5804__A _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8077__A1 _8080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8077__B2 _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5523__B _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput350 sports_i[86] vssd1 vssd1 vccd1 vccd1 _8029_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput361 sports_i[96] vssd1 vssd1 vccd1 vccd1 _8180_/A sky130_fd_sc_hd__buf_2
XANTENNA_output412_A _8057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6635__A _6635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7588__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7230__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5063__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6260__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8001__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8552__A2 _8165_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5620_ _5619_/X _5553_/X _6547_/A vssd1 vssd1 vccd1 vccd1 _5620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5366__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5551_ _5635_/A1 _8709_/B input42/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5551_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_42_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4502_ _4502_/A hold10/A vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__and2_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8270_ _8496_/S vssd1 vssd1 vccd1 vccd1 _8518_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5482_ _6481_/B _5482_/B vssd1 vssd1 vccd1 vccd1 _5482_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7221_ _7220_/X _6908_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7222_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4433_ _8578_/B _4689_/B vssd1 vssd1 vccd1 vccd1 _7384_/A sky130_fd_sc_hd__nor2_8
XANTENNA__6866__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7152_ _7152_/A vssd1 vssd1 vccd1 vccd1 _7152_/X sky130_fd_sc_hd__buf_1
XANTENNA__8068__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4364_ _4693_/B _4719_/B vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7815__A1 _8284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6099_/Y _6102_/Y _8150_/A vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__mux2_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7083_ _7083_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7083_/X sky130_fd_sc_hd__and2_1
X_4295_ _4408_/B _4611_/B vssd1 vssd1 vccd1 vccd1 _4395_/B sky130_fd_sc_hd__nand2_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5826__B1 _5810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6033_/X _6059_/A _6224_/S vssd1 vssd1 vccd1 vccd1 _6035_/A sky130_fd_sc_hd__mux2_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7579__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7985_ _7985_/A1 _7876_/X _7985_/B1 _7836_/B vssd1 vssd1 vccd1 vccd1 _7985_/Y sky130_fd_sc_hd__o22ai_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6251__B1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8791__A2 _8068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _6185_/A _6429_/S _6934_/X _6935_/X vssd1 vssd1 vccd1 vccd1 _6936_/X sky130_fd_sc_hd__a22o_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6867_ _6867_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_147_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7376__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8606_ _7851_/Y _8581_/A _7856_/Y _8583_/A _8689_/S vssd1 vssd1 vccd1 vccd1 _8606_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5818_ _5011_/Y _5817_/Y _5013_/Y vssd1 vssd1 vccd1 vccd1 _5818_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5357__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6798_ _6798_/A _6870_/S vssd1 vssd1 vccd1 vccd1 _6798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8537_ _8261_/A _8820_/A _8153_/X _8584_/A vssd1 vssd1 vccd1 vccd1 _8537_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_134_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4512__B _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5749_ _5749_/A _7847_/A vssd1 vssd1 vccd1 vccd1 _5750_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6306__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8468_ _8468_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8468_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6306__B2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7503__B1 _7640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8919__B hold10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7419_ _7701_/A _7418_/A _7359_/A _5364_/Y vssd1 vssd1 vccd1 vccd1 _7419_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__7823__B _8189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6857__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8399_ _8323_/X _8393_/X _8397_/X _8398_/X vssd1 vssd1 vccd1 vccd1 _8399_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6439__B _6440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7267__C1 _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7806__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__C _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7282__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5293__A1 _5280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7034__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8231__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8231__B2 _8234_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__A1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6242__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7286__A _7286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8534__A2 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8298__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5520__A2 _5764_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7273__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8564__B _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput180 mports_i[56] vssd1 vssd1 vccd1 vccd1 _6401_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput191 mports_i[66] vssd1 vssd1 vccd1 vccd1 _5208_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__8222__A1 _4312_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7025__A2 _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8222__B2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6084__B _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7430__C1 _7756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7770_ _5185_/A _4318_/B _4481_/B _5682_/B vssd1 vssd1 vccd1 vccd1 _7770_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5587__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4982_ _6024_/A vssd1 vssd1 vccd1 vccd1 _6456_/B sky130_fd_sc_hd__inv_6
XFILLER_0_19_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6721_ _7526_/B _6925_/B vssd1 vssd1 vccd1 vccd1 _6721_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7196__A _7196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5709__A _7532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5339__A2 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6652_ _5460_/X _6429_/S _6651_/X vssd1 vssd1 vccd1 vccd1 _6652_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5603_ _5274_/A _5640_/A1 _5275_/X input43/X vssd1 vssd1 vccd1 vccd1 _5603_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6583_ _7396_/B _6871_/B vssd1 vssd1 vccd1 vccd1 _6583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8322_ _8322_/A vssd1 vssd1 vccd1 vccd1 _8322_/X sky130_fd_sc_hd__buf_1
XFILLER_0_54_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5534_ _5534_/A vssd1 vssd1 vccd1 vccd1 _7488_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8253_ _7777_/A _8252_/X _7792_/A vssd1 vssd1 vccd1 vccd1 _8253_/X sky130_fd_sc_hd__o21ba_1
Xoutput610 _5742_/X vssd1 vssd1 vccd1 vccd1 sports_o[198] sky130_fd_sc_hd__buf_12
X_5465_ _5465_/A vssd1 vssd1 vccd1 vccd1 _5465_/Y sky130_fd_sc_hd__inv_2
Xoutput621 _6010_/X vssd1 vssd1 vccd1 vccd1 sports_o[207] sky130_fd_sc_hd__buf_12
XFILLER_0_111_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5444__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput632 _6250_/X vssd1 vssd1 vccd1 vccd1 sports_o[217] sky130_fd_sc_hd__buf_12
X_7204_ _7204_/A vssd1 vssd1 vccd1 vccd1 _7204_/X sky130_fd_sc_hd__buf_1
Xoutput643 _6403_/Y vssd1 vssd1 vccd1 vccd1 sports_o[227] sky130_fd_sc_hd__buf_12
X_4416_ _4416_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__nand2_1
X_8184_ _8820_/A _7872_/A _7975_/A vssd1 vssd1 vccd1 vccd1 _8184_/X sky130_fd_sc_hd__a21o_1
Xoutput654 _7176_/X vssd1 vssd1 vccd1 vccd1 sports_o[31] sky130_fd_sc_hd__buf_12
XFILLER_0_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput665 _7222_/X vssd1 vssd1 vccd1 vccd1 sports_o[41] sky130_fd_sc_hd__buf_12
X_5396_ _6284_/A _5094_/A _5762_/A _6633_/A _5395_/X vssd1 vssd1 vccd1 vccd1 _5397_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput676 _7271_/X vssd1 vssd1 vccd1 vccd1 sports_o[51] sky130_fd_sc_hd__buf_12
XANTENNA__6974__S _7001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput687 _6487_/X vssd1 vssd1 vccd1 vccd1 sports_o[61] sky130_fd_sc_hd__buf_12
X_7135_ _5634_/B _7023_/X _7134_/X vssd1 vssd1 vccd1 vccd1 _7135_/X sky130_fd_sc_hd__o21a_1
Xoutput698 _6615_/X vssd1 vssd1 vccd1 vccd1 sports_o[71] sky130_fd_sc_hd__buf_12
X_4347_ _5129_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__nand2_1
X_7066_ _6550_/A _7059_/X _7383_/A _7246_/B _7061_/X vssd1 vssd1 vccd1 vccd1 _7066_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__8461__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6472__B1 _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6017_ _6017_/A _6017_/B vssd1 vssd1 vccd1 vccd1 _6017_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8749__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8213__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__A1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6224__A0 _6223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4507__B _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__B2 _4940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8490__A _8490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5578__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7968_ _7971_/A1 _5780_/X _7971_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7968_/Y sky130_fd_sc_hd__o22ai_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6775__B2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7818__B _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6919_ _6919_/A _7678_/B vssd1 vssd1 vccd1 vccd1 _6919_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7899_ _7896_/Y _7013_/A _7897_/Y _5117_/A _7898_/Y vssd1 vssd1 vccd1 vccd1 _8346_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_119_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6527__B2 _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7272__C _7272_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6185__A _6185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8204__A1 _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5569__A2 _5558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6766__A1 _6926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6632__B _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8507__A2 _8299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6124__S _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4433__A _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6518__B2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7463__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5250_ input92/X _8310_/B input29/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7494__A2 _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8575__A _8590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5181_ _6550_/A _5682_/B _8188_/S _5218_/A vssd1 vssd1 vccd1 vccd1 _6593_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8443__A1 _8042_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6454__B1 _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold12_A hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8940_ _4595_/B _7707_/B _8942_/A vssd1 vssd1 vccd1 vccd1 _8941_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4608__A _6102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6095__A _6095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8871_ _8871_/A vssd1 vssd1 vccd1 vccd1 _8872_/B sky130_fd_sc_hd__inv_2
XANTENNA__5009__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4327__B _7818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7403__C1 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7822_ _7829_/B vssd1 vssd1 vccd1 vccd1 _7823_/A sky130_fd_sc_hd__inv_2
XANTENNA__6757__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7753_ _7753_/A _7753_/B vssd1 vssd1 vccd1 vccd1 _7753_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7638__B _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4965_ input81/X _8706_/B input18/X _4940_/X vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6542__B _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5439__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6704_ _6506_/A _5634_/B _6449_/A vssd1 vssd1 vccd1 vccd1 _6704_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4343__A hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7684_ _6144_/X _7619_/B _7682_/X _7756_/A _7683_/X vssd1 vssd1 vccd1 vccd1 _7684_/X
+ sky130_fd_sc_hd__a221o_1
X_4896_ _4896_/A vssd1 vssd1 vccd1 vccd1 _8579_/C sky130_fd_sc_hd__buf_12
XFILLER_0_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6635_ _6635_/A vssd1 vssd1 vccd1 vccd1 _6635_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6566_ _6801_/A _6566_/B vssd1 vssd1 vccd1 vccd1 _6566_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5732__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8469__B _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8305_ _7825_/X _8299_/X _8303_/X _8304_/X vssd1 vssd1 vccd1 vccd1 _8306_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5517_ _6780_/A _5445_/X _5516_/X vssd1 vssd1 vccd1 vccd1 _5517_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8131__B1 _8130_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6497_ _6852_/A _6497_/B vssd1 vssd1 vccd1 vccd1 _6497_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5174__A _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8236_ _8235_/Y _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _8236_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5448_ _6634_/A _5077_/A _6017_/A _6648_/B vssd1 vssd1 vccd1 vccd1 _6644_/A sky130_fd_sc_hd__a22o_1
Xoutput440 _8350_/Y vssd1 vssd1 vccd1 vccd1 mports_o[44] sky130_fd_sc_hd__buf_12
XANTENNA__5496__A1 _5435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput451 _8475_/X vssd1 vssd1 vccd1 vccd1 mports_o[54] sky130_fd_sc_hd__buf_12
XANTENNA__6693__A0 _5539_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5496__B2 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput462 _8561_/X vssd1 vssd1 vccd1 vccd1 mports_o[64] sky130_fd_sc_hd__buf_12
Xoutput473 _8612_/X vssd1 vssd1 vccd1 vccd1 mports_o[74] sky130_fd_sc_hd__buf_12
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput484 _8646_/X vssd1 vssd1 vccd1 vccd1 mports_o[84] sky130_fd_sc_hd__buf_12
X_8167_ _6017_/A _8172_/B _8189_/B _8166_/Y vssd1 vssd1 vccd1 vccd1 _8167_/X sky130_fd_sc_hd__a211o_1
X_5379_ input96/X _8310_/B input33/X _4874_/X vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__o22a_1
Xoutput495 _8680_/X vssd1 vssd1 vccd1 vccd1 mports_o[94] sky130_fd_sc_hd__buf_12
XFILLER_0_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7118_ _7117_/X _5496_/X _7175_/S vssd1 vssd1 vccd1 vccd1 _7119_/A sky130_fd_sc_hd__mux2_2
XANTENNA__7237__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8098_ _8098_/A vssd1 vssd1 vccd1 vccd1 _8098_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6445__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7049_ _7272_/A _6499_/A _7138_/A vssd1 vssd1 vccd1 vccd1 _7049_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4518__A _4518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8737__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7829__A _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5420__A1 _5401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5420__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5708__C1 _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7173__A1 _5827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5184__B1 _6526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6920__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7283__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8673__A1 _8519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6684__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6908__A _6908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7228__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7779__A3 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6987__A1 _6358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8842__B _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8728__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6739__A1 _5738_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6739__B2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5411__A1 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750_ _4761_/A _4770_/A _4750_/C vssd1 vssd1 vccd1 vccd1 _4752_/A sky130_fd_sc_hd__nand3_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5962__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6789__S _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4681_ _4681_/A _4681_/B vssd1 vssd1 vccd1 vccd1 _4682_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7164__A1 _5770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5693__S _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7474__A _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6420_ _6506_/A _6528_/A vssd1 vssd1 vccd1 vccd1 _6946_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_114_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6351_ input75/X _8579_/C _6357_/A1 _8713_/C _6350_/X vssd1 vssd1 vccd1 vccd1 _6352_/A
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_141_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8113__B1 _8111_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5302_ _6780_/A _6591_/B _5301_/X vssd1 vssd1 vccd1 vccd1 _5303_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7467__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5425__C _5425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6282_ _5185_/A _6283_/A _6322_/B _6875_/B vssd1 vssd1 vccd1 vccd1 _6282_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5478__A1 _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5478__B2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8021_ _8024_/A1 _5780_/A _8024_/B1 _5079_/A vssd1 vssd1 vccd1 vccd1 _8021_/Y sky130_fd_sc_hd__o22ai_2
X_5233_ _6212_/A _6566_/B _5108_/A _6597_/B _5136_/X vssd1 vssd1 vccd1 vccd1 _5233_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5722__A _5722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7219__A2 _7059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5164_ _8444_/A _5208_/A1 _8257_/C _5208_/B1 vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__a22o_1
X_5095_ _5682_/B _5088_/X _5094_/Y vssd1 vssd1 vccd1 vccd1 _5095_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8923_ _8922_/A _4760_/B hold16/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8719__A2 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5650__A1 _5622_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8854_ _7372_/B _8852_/X _8853_/X vssd1 vssd1 vccd1 vccd1 _8968_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7805_ _7760_/X _7796_/X _7801_/X _7804_/Y vssd1 vssd1 vccd1 vccd1 _7805_/X sky130_fd_sc_hd__a22o_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8785_ _8784_/X _8042_/Y _8788_/S vssd1 vssd1 vccd1 vccd1 _8785_/X sky130_fd_sc_hd__mux2_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _5997_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5997_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5169__A _6558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7736_ _4793_/A _7723_/B _7735_/X vssd1 vssd1 vccd1 vccd1 _7736_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4948_ _5893_/B vssd1 vssd1 vccd1 vccd1 _6266_/A sky130_fd_sc_hd__inv_2
XANTENNA__5953__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7155__A1 _7544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7667_ _7663_/X _7665_/Y _7666_/Y vssd1 vssd1 vccd1 vccd1 _7667_/X sky130_fd_sc_hd__a21o_1
X_4879_ _8709_/A _5780_/A vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7384__A _7384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6618_ _6432_/X _6617_/Y _6436_/A vssd1 vssd1 vccd1 vccd1 _6618_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5705__A2 _5625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7598_ _7599_/B _7691_/B vssd1 vssd1 vccd1 vccd1 _7598_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6902__A1 _6112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6549_ _6549_/A vssd1 vssd1 vccd1 vccd1 _6913_/B sky130_fd_sc_hd__buf_6
XANTENNA__4520__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8655__A1 _8055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7458__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5469__A1 _6671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5469__B2 _6679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8219_ _4478_/B _6500_/X _8221_/A2 _7769_/X _8218_/X vssd1 vssd1 vccd1 vccd1 _8219_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6130__A2 _6094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6969__A1 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5641__A1 _5601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7918__B1 _7918_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7278__B _7288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8040__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8591__B1 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5079__A _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5944__A2 _5930_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7146__A1 _5655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8343__B1 _7929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5526__B _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8646__A1 _8412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6657__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6121__A2 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5880__A1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5880__B2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7621__A2 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5632__A1 _6870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5920_ _5159_/B _5885_/X _5125_/X _5901_/X _5919_/X vssd1 vssd1 vccd1 vccd1 _5920_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5851_ _5159_/B _5824_/X _5846_/X _5847_/X _5850_/Y vssd1 vssd1 vccd1 vccd1 _5851_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4802_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8570_ _8247_/Y _8299_/A _8249_/X _8304_/A _8269_/A vssd1 vssd1 vccd1 vccd1 _8570_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5396__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5782_ _5782_/A _8578_/B vssd1 vssd1 vccd1 vccd1 _5782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7521_ _5648_/Y _7619_/B _7517_/X _7519_/X _7520_/Y vssd1 vssd1 vccd1 vccd1 _7521_/X
+ sky130_fd_sc_hd__a221o_2
X_4733_ _4733_/A _4733_/B vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7452_ _6634_/A _7542_/A _7694_/A _6644_/A _7326_/A vssd1 vssd1 vccd1 vccd1 _7452_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4664_ hold20/X vssd1 vssd1 vccd1 vccd1 _8574_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5699__A1 _5718_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6403_ _6399_/Y _6402_/A _6402_/Y vssd1 vssd1 vccd1 vccd1 _6403_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__5699__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7383_ _7383_/A _7630_/B vssd1 vssd1 vccd1 vccd1 _7383_/Y sky130_fd_sc_hd__nand2_1
X_4595_ _4604_/A _4595_/B _4612_/B vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6334_ _6321_/A _6547_/A _5762_/A vssd1 vssd1 vccd1 vccd1 _6334_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__8637__A1 _8394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8637__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6265_ _6312_/A _6263_/X _6264_/X vssd1 vssd1 vccd1 vccd1 _6267_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8004_ _8011_/A1 _4946_/A _8011_/B1 _5119_/A vssd1 vssd1 vccd1 vccd1 _8004_/Y sky130_fd_sc_hd__o22ai_2
X_5216_ input12/X _4929_/A _5222_/B1 _4932_/A _5215_/X vssd1 vssd1 vccd1 vccd1 _6567_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6267__B _6375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6196_ _6234_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6196_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5171__B _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5147_ _7055_/A _5909_/B _5146_/Y _7629_/B vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__a22o_1
XANTENNA__7073__A0 _7072_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7612__A2 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5078_ _7299_/A vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__buf_8
XANTENNA__5623__A1 _5637_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5623__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6283__A _6283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8906_ _4821_/A _4819_/C hold21/X _8904_/B vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8837_ _8835_/Y _8836_/X _4662_/C _8806_/B vssd1 vssd1 vccd1 vccd1 _8837_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5387__B1 _5275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8768_ _8767_/X _7972_/Y _8788_/S vssd1 vssd1 vccd1 vccd1 _8768_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7719_ _6287_/X _7723_/B _7718_/X vssd1 vssd1 vccd1 vccd1 _7719_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__7128__A1 _5548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8325__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7318__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8699_ _8695_/X _8698_/Y _8226_/X _8590_/X vssd1 vssd1 vccd1 vccd1 _8699_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7679__A2 _7686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8946__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5346__B _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6351__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7842__A _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8628__A1 _8381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6458__A _6724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5362__A _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7064__A0 _7063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8800__A1 _8503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7603__A2 _5860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8800__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__A1 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7367__B2 _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5378__B1 _5386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8867__A1 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8619__A1 _8346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5550__B1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4380_ hold46/X _4380_/B vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__or2_1
XANTENNA__8567__B _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8095__A2 _8516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5272__A _5272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6047_/Y _4886_/A _6048_/Y _4891_/A _6049_/Y vssd1 vssd1 vccd1 vccd1 _6897_/A
+ sky130_fd_sc_hd__o221a_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__A1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__A2 _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5001_ _6024_/A vssd1 vssd1 vccd1 vccd1 _6080_/A sky130_fd_sc_hd__buf_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8583__A _8583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6952_ _6951_/X _7707_/D _7000_/S vssd1 vssd1 vccd1 vccd1 _6952_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5081__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5903_ _5871_/A _8335_/B _5872_/A _4913_/A _5902_/X vssd1 vssd1 vccd1 vccd1 _6828_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__4335__B _7847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6883_ _6063_/A _6506_/A _6968_/A _6879_/X _6882_/Y vssd1 vssd1 vccd1 vccd1 _6883_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8622_ _8621_/X _7912_/Y _8686_/B vssd1 vssd1 vccd1 vccd1 _8623_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5834_ _5011_/Y _5828_/Y _5832_/Y _7629_/B _5833_/Y vssd1 vssd1 vccd1 vccd1 _5834_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6030__A1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6030__B2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5765_ _5518_/A _5102_/A _5519_/A _5191_/A _5764_/X vssd1 vssd1 vccd1 vccd1 _5765_/X
+ sky130_fd_sc_hd__o221a_4
X_8553_ _8549_/X _8299_/A _8552_/X _8304_/A _8269_/A vssd1 vssd1 vccd1 vccd1 _8553_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6550__B _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4716_ _4716_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4351__A _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7504_ _5552_/X _7686_/A _7694_/A _5573_/X _7503_/Y vssd1 vssd1 vccd1 vccd1 _7505_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8484_ _8483_/Y _8455_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8484_/X sky130_fd_sc_hd__mux2_1
X_5696_ _6170_/A _5696_/B vssd1 vssd1 vccd1 vccd1 _5696_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7435_ _5094_/A _7640_/B _7431_/X _7434_/Y vssd1 vssd1 vccd1 vccd1 _7436_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6977__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4647_ _8958_/Q hold44/A vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_32_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8946__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7530__A1 _7683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7366_ _7686_/A _7366_/B vssd1 vssd1 vccd1 vccd1 _7366_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_114_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _4823_/B vssd1 vssd1 vccd1 vccd1 _4578_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6317_ _6326_/A1 _8444_/A input9/X _8257_/C _6316_/Y vssd1 vssd1 vccd1 vccd1 _6317_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_40_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7297_ _7510_/B _7297_/B vssd1 vssd1 vccd1 vccd1 _7660_/B sky130_fd_sc_hd__nor2_8
XANTENNA__6278__A _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6097__A1 _6140_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6097__B2 _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6248_ _6248_/A1 _4930_/X input5/X _4933_/X _6247_/X vssd1 vssd1 vccd1 vccd1 _6248_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__7833__A2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6179_ _6179_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _6179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7597__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6725__B _7532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5072__A2 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8432__S _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8010__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6572__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6324__A2 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8077__A2 _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6188__A _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6088__A1 _6107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5835__A1 _5902_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5835__B2 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput340 sports_i[77] vssd1 vssd1 vccd1 vccd1 _7918_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__5820__A _5820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput351 sports_i[87] vssd1 vssd1 vccd1 vccd1 _8054_/B1 sky130_fd_sc_hd__buf_2
Xinput362 sports_i[97] vssd1 vssd1 vccd1 vccd1 _8198_/B sky130_fd_sc_hd__buf_2
XANTENNA__7588__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6260__B2 _4913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8537__B1 _8153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8001__A2 _8400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6012__A1 _6020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6012__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7466__B _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8969__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _5516_/B _7629_/B _6837_/A _5909_/B _5549_/Y vssd1 vssd1 vccd1 vccd1 _5550_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4501_ _4551_/B vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__inv_2
XFILLER_0_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5481_ _5738_/C _5077_/A _6017_/A _7551_/A vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7220_ _6102_/A _7138_/X _7218_/X _7219_/X vssd1 vssd1 vccd1 vccd1 _7220_/X sky130_fd_sc_hd__o22a_2
X_4432_ hold32/X vssd1 vssd1 vccd1 vccd1 _4689_/B sky130_fd_sc_hd__inv_2
XFILLER_0_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7151_ _7150_/X _6743_/A _7175_/S vssd1 vssd1 vccd1 vccd1 _7152_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8068__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ _4681_/B _4818_/B vssd1 vssd1 vccd1 vccd1 _4693_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6102_ _6102_/A _6102_/B vssd1 vssd1 vccd1 vccd1 _6102_/Y sky130_fd_sc_hd__nand2_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7815__A2 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7082_ _7082_/A vssd1 vssd1 vccd1 vccd1 _7082_/X sky130_fd_sc_hd__buf_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _8968_/Q vssd1 vssd1 vccd1 vccd1 _4408_/B sky130_fd_sc_hd__clkinv_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5826__A1 _5809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5826__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6033_ _6030_/X _6867_/A _6356_/S vssd1 vssd1 vccd1 vccd1 _6033_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6003__B1_N _5013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7028__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5730__A _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7579__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7984_ _8394_/A _7954_/X _7983_/Y _7772_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _7984_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6251__A1 _6262_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6251__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6935_ _6958_/B _6212_/B _6450_/A vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5876__S _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4801__A2 _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7657__A _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6866_ _6864_/X _6933_/A _6968_/A _6865_/X vssd1 vssd1 vccd1 vccd1 _6866_/X sky130_fd_sc_hd__a211o_2
XFILLER_0_92_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8605_ _7821_/Y _8577_/X _8603_/X _8604_/Y vssd1 vssd1 vccd1 vccd1 _8605_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5817_ _6304_/A _5829_/C vssd1 vssd1 vccd1 vccd1 _5817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6797_ _6797_/A vssd1 vssd1 vccd1 vccd1 _6798_/A sky130_fd_sc_hd__inv_2
XFILLER_0_146_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6554__A2 _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8536_ _4933_/X _8821_/A _4940_/X _8137_/X _8535_/Y vssd1 vssd1 vccd1 vccd1 _8806_/A
+ sky130_fd_sc_hd__o221a_1
X_5748_ _5829_/C vssd1 vssd1 vccd1 vccd1 _7167_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6306__A2 _6277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8467_ _8513_/B _8418_/Y _8304_/A _8466_/Y vssd1 vssd1 vccd1 vccd1 _8467_/X sky130_fd_sc_hd__o211a_1
X_5679_ _5679_/A _5741_/B vssd1 vssd1 vccd1 vccd1 _5679_/X sky130_fd_sc_hd__and2_1
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8700__B1 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7418_ _7418_/A _7691_/B vssd1 vssd1 vccd1 vccd1 _7418_/Y sky130_fd_sc_hd__nand2_1
X_8398_ _8564_/B _8772_/B _8497_/S vssd1 vssd1 vccd1 vccd1 _8398_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7349_ _7349_/A vssd1 vssd1 vccd1 vccd1 _7349_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7806__A2 _7813_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__D _5062_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5293__A2 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7535__A2_N _7348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8767__B1 _7969_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8231__A2 _8234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6242__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6242__B2 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8961__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5087__A _6489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8298__A2 _8297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6646__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8207__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput170 mports_i[47] vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__clkbuf_2
Xinput181 mports_i[57] vssd1 vssd1 vccd1 vccd1 _4888_/A sky130_fd_sc_hd__clkbuf_2
Xinput192 mports_i[67] vssd1 vssd1 vccd1 vccd1 _5222_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__8222__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7430__B1 _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4981_ _4981_/A vssd1 vssd1 vccd1 vccd1 _7027_/A sky130_fd_sc_hd__inv_2
XANTENNA__7981__B2 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4795__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6720_ _6720_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6651_ _6643_/X _6871_/B _6649_/X _6467_/X _6650_/Y vssd1 vssd1 vccd1 vccd1 _6651_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5602_ _5602_/A vssd1 vssd1 vccd1 vccd1 _5602_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5744__B1 _5519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6582_ _6689_/S _5246_/X _6581_/Y vssd1 vssd1 vccd1 vccd1 _7396_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8321_ _8318_/X _8320_/X _8572_/S vssd1 vssd1 vccd1 vccd1 _8322_/A sky130_fd_sc_hd__mux2_1
X_5533_ _5500_/X _7299_/A _6281_/S _6697_/B vssd1 vssd1 vccd1 vccd1 _5534_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8252_ _8252_/A1 _7536_/B _8252_/B1 _5230_/B _8251_/X vssd1 vssd1 vccd1 vccd1 _8252_/X
+ sky130_fd_sc_hd__a221o_4
X_5464_ _5440_/A _8523_/B _5441_/A _4933_/A _5463_/X vssd1 vssd1 vccd1 vccd1 _5464_/X
+ sky130_fd_sc_hd__o221a_4
Xoutput600 _5494_/X vssd1 vssd1 vccd1 vccd1 sports_o[189] sky130_fd_sc_hd__buf_12
Xoutput611 _5779_/X vssd1 vssd1 vccd1 vccd1 sports_o[199] sky130_fd_sc_hd__buf_12
XFILLER_0_42_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput622 _6035_/X vssd1 vssd1 vccd1 vccd1 sports_o[208] sky130_fd_sc_hd__buf_12
XFILLER_0_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7203_ _7202_/X _6059_/A _7249_/S vssd1 vssd1 vccd1 vccd1 _7204_/A sky130_fd_sc_hd__mux2_2
Xoutput633 _6268_/X vssd1 vssd1 vccd1 vccd1 sports_o[218] sky130_fd_sc_hd__buf_12
XFILLER_0_1_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5444__B _6653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4415_ _4415_/A _4425_/B _4425_/A vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__nand3_1
X_8183_ _8189_/C _7874_/A _8196_/B1 _8174_/A _8182_/X vssd1 vssd1 vccd1 vccd1 _8820_/A
+ sky130_fd_sc_hd__a221oi_4
Xoutput644 _7133_/X vssd1 vssd1 vccd1 vccd1 sports_o[22] sky130_fd_sc_hd__buf_12
XFILLER_0_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5395_ _5909_/B _5336_/Y _5394_/Y _5997_/B _6234_/B vssd1 vssd1 vccd1 vccd1 _5395_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput655 _7182_/X vssd1 vssd1 vccd1 vccd1 sports_o[32] sky130_fd_sc_hd__buf_12
XFILLER_0_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput666 _7227_/X vssd1 vssd1 vccd1 vccd1 sports_o[42] sky130_fd_sc_hd__buf_12
XANTENNA__7946__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput677 _7276_/X vssd1 vssd1 vccd1 vccd1 sports_o[52] sky130_fd_sc_hd__buf_12
X_7134_ _5552_/X _7004_/X _5595_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7134_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_100_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4346_ _4346_/A vssd1 vssd1 vccd1 vccd1 _4818_/B sky130_fd_sc_hd__buf_6
Xoutput688 _6493_/X vssd1 vssd1 vccd1 vccd1 sports_o[62] sky130_fd_sc_hd__buf_12
Xoutput699 _6625_/X vssd1 vssd1 vccd1 vccd1 sports_o[72] sky130_fd_sc_hd__buf_12
X_7065_ _7065_/A vssd1 vssd1 vccd1 vccd1 _7065_/X sky130_fd_sc_hd__buf_1
XANTENNA__8461__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7151__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6016_ _6016_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _6017_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4483__B1 _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8749__B1 _8362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8213__A2 _8200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__A2 _8706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6224__A1 _6941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8490__B _8491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7967_ _7962_/Y _6080_/A _7963_/Y _6513_/A _7966_/Y vssd1 vssd1 vccd1 vccd1 _8404_/A
+ sky130_fd_sc_hd__a221oi_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7972__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6918_ _6907_/Y _6511_/A _6908_/Y _6917_/X vssd1 vssd1 vccd1 vccd1 _6918_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7898_ _7905_/A1 _4946_/A _7905_/B1 _5119_/A vssd1 vssd1 vccd1 vccd1 _7898_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6849_ _5924_/A _6510_/A _5901_/X _6512_/A vssd1 vssd1 vccd1 vccd1 _6849_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7724__A1 _6310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8519_ _8519_/A _8523_/B vssd1 vssd1 vccd1 vccd1 _8519_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6466__A _6466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5370__A _6611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6463__B2 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6185__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8204__A2 _8198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6913__B _6913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7297__A _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7715__A1 _6261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6151__B1 _6158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7760__A _7975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5180_ input12/X _5080_/A _5222_/B1 _5089_/X _5179_/X vssd1 vssd1 vccd1 vccd1 _5218_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__8443__A2 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5280__A _5280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6454__A1 _4876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6095__B _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4465__B1 _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8870_ _8877_/B _8870_/B vssd1 vssd1 vccd1 vccd1 _8871_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6206__B2 _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7403__B1 _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7821_ _7821_/A vssd1 vssd1 vccd1 vccd1 _7821_/Y sky130_fd_sc_hd__inv_2
X_7752_ _7694_/A _6395_/A _7542_/A _7306_/A _6397_/X vssd1 vssd1 vccd1 vccd1 _7752_/Y
+ sky130_fd_sc_hd__o2111ai_1
X_4964_ _4961_/X _4963_/X _6356_/S vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6703_ _6699_/Y _6701_/X _6702_/X _5645_/A _6429_/S vssd1 vssd1 vccd1 vccd1 _6703_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5439__B _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4895_ _5275_/A vssd1 vssd1 vccd1 vccd1 _4896_/A sky130_fd_sc_hd__buf_8
XANTENNA__6509__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7683_ _7683_/A _7683_/B _7683_/C vssd1 vssd1 vccd1 vccd1 _7683_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5717__B1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6634_ _6634_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6565_ _6565_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6565_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7146__S _7175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8304_ _8304_/A vssd1 vssd1 vccd1 vccd1 _8304_/X sky130_fd_sc_hd__clkbuf_8
X_5516_ _6711_/S _5516_/B vssd1 vssd1 vccd1 vccd1 _5516_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6496_ _6919_/A vssd1 vssd1 vccd1 vccd1 _6852_/A sky130_fd_sc_hd__buf_6
XFILLER_0_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8131__A1 _8550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8131__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8235_ _8235_/A1 _7536_/B _8235_/B1 _5230_/B _8234_/X vssd1 vssd1 vccd1 vccd1 _8235_/Y
+ sky130_fd_sc_hd__a221oi_4
X_5447_ _5999_/B _7105_/A _6668_/A _5174_/A vssd1 vssd1 vccd1 vccd1 _5447_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6142__B1 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput430 _8279_/X vssd1 vssd1 vccd1 vccd1 mports_o[35] sky130_fd_sc_hd__buf_12
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput441 _8357_/X vssd1 vssd1 vccd1 vccd1 mports_o[45] sky130_fd_sc_hd__buf_12
XFILLER_0_140_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput452 _8489_/X vssd1 vssd1 vccd1 vccd1 mports_o[55] sky130_fd_sc_hd__buf_12
XANTENNA__5496__A2 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput463 _8565_/X vssd1 vssd1 vccd1 vccd1 mports_o[65] sky130_fd_sc_hd__buf_12
X_5378_ _5385_/A _4868_/A _5386_/A _4870_/A _5377_/X vssd1 vssd1 vccd1 vccd1 _6634_/A
+ sky130_fd_sc_hd__o221a_4
Xoutput474 _8616_/X vssd1 vssd1 vccd1 vccd1 mports_o[75] sky130_fd_sc_hd__buf_12
X_8166_ _8166_/A _8171_/B vssd1 vssd1 vccd1 vccd1 _8166_/Y sky130_fd_sc_hd__nor2_1
Xoutput485 _8650_/X vssd1 vssd1 vccd1 vccd1 mports_o[85] sky130_fd_sc_hd__buf_12
Xoutput496 _8683_/X vssd1 vssd1 vccd1 vccd1 mports_o[95] sky130_fd_sc_hd__buf_12
X_7117_ _5498_/X _7026_/X _7115_/X _7116_/X vssd1 vssd1 vccd1 vccd1 _7117_/X sky130_fd_sc_hd__o22a_1
X_4329_ _4329_/A _8185_/B vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__nand2_1
X_8097_ _8097_/A vssd1 vssd1 vccd1 vccd1 _8097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5190__A _6526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7048_ _7048_/A vssd1 vssd1 vccd1 vccd1 _7048_/X sky130_fd_sc_hd__buf_1
XANTENNA__4518__B _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7829__B _7829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6733__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6748__A2 _5765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7945__B2 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5420__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7158__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8440__S _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7173__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6381__B1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5184__B2 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8658__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8122__A1 _7975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8673__A2 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6684__A1 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6908__B _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6196__A _6234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8615__S _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6924__A _6924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6739__A2 _6549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4680_ _4714_/A _4680_/B vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5175__A1 _5909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6372__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5175__B2 _5997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5275__A _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6350_ _8444_/A _6358_/A1 _8257_/C input13/X vssd1 vssd1 vccd1 vccd1 _6350_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_70_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8113__B2 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5301_ _6711_/S _5301_/B vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6281_ _6278_/Y _6971_/A _6281_/S vssd1 vssd1 vccd1 vccd1 _6322_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5478__A2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5232_ _5227_/X _5228_/X _6689_/S vssd1 vssd1 vccd1 vccd1 _6597_/B sky130_fd_sc_hd__mux2_1
XANTENNA__6675__A1 _5496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8020_ _8015_/Y _6079_/A _8016_/Y _6513_/A _8019_/Y vssd1 vssd1 vccd1 vccd1 _8427_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6818__B _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5163_ _5299_/B _7055_/A _5161_/X _6470_/B vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5094_ _5094_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5094_/Y sky130_fd_sc_hd__nand2_1
X_8922_ _8922_/A hold15/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5650__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8853_ _8857_/A _7761_/A _6264_/X _4611_/A vssd1 vssd1 vccd1 vccd1 _8853_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7927__B2 _6411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7804_ _7803_/Y _7774_/X _7975_/A vssd1 vssd1 vccd1 vccd1 _7804_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5938__B1 _5275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8784_ _8445_/A _8738_/A _8468_/A _8711_/A vssd1 vssd1 vccd1 vccd1 _8784_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5996_ _5995_/X _5942_/X _6711_/S vssd1 vssd1 vccd1 vccd1 _5997_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7735_ _7272_/B _7349_/A _6980_/Y _7753_/B _7749_/S vssd1 vssd1 vccd1 vccd1 _7735_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4947_ _8759_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _5893_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7666_ _7590_/A _7665_/A _7372_/A _6907_/Y vssd1 vssd1 vccd1 vccd1 _7666_/Y sky130_fd_sc_hd__o22ai_1
X_4878_ _6084_/B vssd1 vssd1 vccd1 vccd1 _6284_/A sky130_fd_sc_hd__inv_8
XFILLER_0_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7155__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7384__B _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6617_ _6852_/A _7094_/A vssd1 vssd1 vccd1 vccd1 _6617_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6363__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7597_ _7378_/X _5885_/X _7683_/C vssd1 vssd1 vccd1 vccd1 _7599_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__6902__A2 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5185__A _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6548_ _6547_/A _6545_/X _6854_/A _6547_/Y vssd1 vssd1 vccd1 vccd1 _6548_/X sky130_fd_sc_hd__a211o_1
XANTENNA__8104__B2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6479_ _5028_/X _6429_/S _6478_/X vssd1 vssd1 vccd1 vccd1 _6479_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_112_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5469__A2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7863__B1 _7760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8218_ _5185_/A _8222_/B1 _4312_/B _5682_/B vssd1 vssd1 vccd1 vccd1 _8218_/X sky130_fd_sc_hd__a22o_1
X_8149_ _8145_/Y _7954_/X _8148_/X _7826_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8149_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4529__A _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8812__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6969__A2 _6310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7091__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7918__A1 _7918_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7918__B2 _7835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5929__B1 _5867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8591__A1 _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7575__A _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8343__A1 _8359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8343__B2 _8299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6354__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8646__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7854__B1 hold23/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output435_A _7816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output602_A _5528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7621__A3 _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4840__B1 _7309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5850_ _6266_/A _6818_/A vssd1 vssd1 vccd1 vccd1 _5850_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _4814_/B _4818_/B _8716_/A vssd1 vssd1 vccd1 vccd1 _4801_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5396__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5781_ _5781_/A _6481_/B vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_146_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7520_ _7590_/A _7520_/B vssd1 vssd1 vccd1 vccd1 _7520_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4902__A _5999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4732_ _4732_/A _4732_/B vssd1 vssd1 vccd1 vccd1 _4733_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _8857_/A sky130_fd_sc_hd__inv_2
X_7451_ _7451_/A _7668_/B vssd1 vssd1 vccd1 vccd1 _7451_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4621__B _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5209__S _6386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6402_ _6402_/A _7756_/B vssd1 vssd1 vccd1 vccd1 _6402_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5699__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6896__A1 _6095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4594_ _4552_/A _4552_/B _4837_/A vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__a21oi_1
X_7382_ _7575_/A vssd1 vssd1 vccd1 vccd1 _7694_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6333_ _6333_/A vssd1 vssd1 vccd1 vccd1 _6333_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8637__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6264_ _7398_/A vssd1 vssd1 vccd1 vccd1 _6264_/X sky130_fd_sc_hd__buf_6
X_5215_ input91/X _4935_/A input28/X _4939_/A vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__o22a_1
X_8003_ _8003_/A vssd1 vssd1 vccd1 vccd1 _8003_/Y sky130_fd_sc_hd__inv_2
X_6195_ _6227_/A _5080_/A input4/X _5089_/X _6194_/X vssd1 vssd1 vccd1 vccd1 _6234_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5146_ _5146_/A _6514_/B vssd1 vssd1 vccd1 vccd1 _5146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7073__A1 _6567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5077_ _5077_/A vssd1 vssd1 vccd1 vccd1 _7299_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7612__A3 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5623__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8905_ _4784_/A _4786_/B _8904_/B _8904_/Y vssd1 vssd1 vccd1 vccd1 _8946_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_39_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8836_ _8239_/Y _8803_/B _8240_/Y _8711_/X _8788_/S vssd1 vssd1 vccd1 vccd1 _8836_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5387__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8767_ _8404_/A _8550_/B _8738_/A _7969_/Y _8711_/A vssd1 vssd1 vccd1 vccd1 _8767_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5979_ _6028_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6042_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5908__A _6809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7718_ _7251_/Y _7753_/B _6272_/X _7349_/A _7749_/S vssd1 vssd1 vccd1 vccd1 _7718_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8325__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8698_ _8698_/A _8698_/B vssd1 vssd1 vccd1 vccd1 _8698_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6336__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4531__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7649_ _7532_/A _6074_/A _7348_/A vssd1 vssd1 vccd1 vccd1 _7651_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6887__A1 _6058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7842__B _7858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5362__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A1 _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5311__B2 _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7064__A1 _5159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8800__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7367__A2 _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5378__A1 _5385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5378__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5537__B _6081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7024__B1_N _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8619__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7244__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__A1 _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5003_/A _4913_/X _5004_/A _8516_/B _4999_/X vssd1 vssd1 vccd1 vccd1 _5000_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8252__B1 _8252_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6951_ _6241_/X _6994_/B _7242_/A _6989_/B vssd1 vssd1 vccd1 vccd1 _6951_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_89_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8004__B1 _8011_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5902_ _5902_/A1 _8271_/B input53/X _4917_/A vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6882_ _6882_/A _6882_/B vssd1 vssd1 vccd1 vccd1 _6882_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5369__A1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8621_ _8620_/X _8335_/A _8621_/S vssd1 vssd1 vccd1 vccd1 _8621_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5833_ _6304_/A _7171_/A vssd1 vssd1 vccd1 vccd1 _5833_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6831__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8552_ _4894_/A _8165_/Y _4891_/X _8203_/X _8551_/Y vssd1 vssd1 vccd1 vccd1 _8552_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5764_ _5764_/A1 _5192_/A input48/X _5193_/A vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8307__A1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7503_ _7678_/A _5609_/B _7640_/B vssd1 vssd1 vccd1 vccd1 _7503_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6318__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4715_ _4715_/A _4715_/B vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__nand2_1
X_8483_ _8483_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8483_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4351__B hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5695_ _6284_/A _7524_/A _5762_/A _5684_/X _5694_/X vssd1 vssd1 vccd1 vccd1 _5696_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7434_ _7432_/Y _7433_/Y _7497_/B vssd1 vssd1 vccd1 vccd1 _7434_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4646_ _4818_/B _4927_/A _4823_/B _4931_/A _4645_/X vssd1 vssd1 vccd1 vccd1 _7737_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_115_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5541__A1 _5539_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4577_ _8336_/S hold21/A vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__nand2_8
X_7365_ _5161_/X _7630_/B _6539_/X _7638_/B vssd1 vssd1 vccd1 vccd1 _7365_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6316_ _6314_/Y _6315_/Y _4674_/C vssd1 vssd1 vccd1 vccd1 _6316_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7296_ _7296_/A vssd1 vssd1 vccd1 vccd1 _7296_/X sky130_fd_sc_hd__buf_1
XANTENNA__6097__A2 _5192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6247_ _6247_/A1 _8706_/B input68/X _4940_/X vssd1 vssd1 vccd1 vccd1 _6247_/X sky130_fd_sc_hd__o22a_1
X_6178_ _6103_/X _6177_/X _6870_/S vssd1 vssd1 vccd1 vccd1 _6179_/A sky130_fd_sc_hd__mux2_1
XANTENNA__8243__B1 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ _5129_/A vssd1 vssd1 vccd1 vccd1 _8444_/A sky130_fd_sc_hd__buf_8
XANTENNA__5057__B1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8794__A1 _8081_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7597__A2 _5885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8819_ _8187_/X _8803_/B _8190_/X _8711_/X _8788_/S vssd1 vssd1 vccd1 vccd1 _8819_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6309__B1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7521__A2 _7619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5532__A1 _5575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5532__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6469__A _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7064__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7809__B1 _7814_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5296__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5835__A2 _4871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput330 sports_i[68] vssd1 vssd1 vccd1 vccd1 _4481_/B sky130_fd_sc_hd__clkbuf_4
Xinput341 sports_i[78] vssd1 vssd1 vccd1 vccd1 _7931_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5820__B _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8234__B1 _7875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput352 sports_i[88] vssd1 vssd1 vccd1 vccd1 _8067_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput363 sports_i[98] vssd1 vssd1 vccd1 vccd1 _4312_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4717__A hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5048__B1 _4896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6245__C1 _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8785__A1 _8042_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7588__A2 _5853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5599__B2 _4890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6796__B1 _8151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6260__A2 _8516_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6548__B1 _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7239__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6012__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5220__B1 _6170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5771__A1 _5787_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5771__B2 _4938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4500_ _4613_/B _4658_/A vssd1 vssd1 vccd1 vccd1 _4551_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5480_ _5518_/A _4868_/A _5519_/A _5089_/A _5479_/X vssd1 vssd1 vccd1 vccd1 _7551_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8170__C1 _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8578__B _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4431_ _8977_/Q vssd1 vssd1 vccd1 vccd1 _8578_/B sky130_fd_sc_hd__buf_12
XANTENNA_1 _6770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4362_ hold33/X vssd1 vssd1 vccd1 vccd1 _4681_/B sky130_fd_sc_hd__inv_2
X_7150_ _6732_/A _7138_/X _7148_/X _7149_/X vssd1 vssd1 vccd1 vccd1 _7150_/X sky130_fd_sc_hd__o22a_2
X_6101_ _6075_/A _4909_/A _6076_/A _5191_/A _6100_/X vssd1 vssd1 vccd1 vccd1 _6102_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7081_ _7080_/X _5328_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7082_/A sky130_fd_sc_hd__mux2_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4393_/B vssd1 vssd1 vccd1 vccd1 _4300_/A sky130_fd_sc_hd__inv_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5287__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5826__A2 _4953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6032_ _5965_/A _8335_/B _5966_/A _4913_/A _6031_/X vssd1 vssd1 vccd1 vccd1 _6867_/A
+ sky130_fd_sc_hd__o221a_4
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5730__B _6737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8225__B1 _8857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8776__A1 _8400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7579__A2 _5824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7983_ _7976_/Y _6500_/X _7977_/Y _7769_/X _7982_/Y vssd1 vssd1 vccd1 vccd1 _7983_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7984__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6251__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6934_ _6932_/X _6933_/A _6968_/A _6933_/Y vssd1 vssd1 vccd1 vccd1 _6934_/X sky130_fd_sc_hd__a211o_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8528__A1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6539__B1 _5161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6865_ _6028_/A _6913_/B _7623_/B _6876_/C vssd1 vssd1 vccd1 vccd1 _6865_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_119_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6003__A2 _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8604_ _7837_/X _8685_/B _8686_/B vssd1 vssd1 vccd1 vccd1 _8604_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5816_ _5816_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5816_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6796_ _6788_/B _5197_/X _8151_/B _6801_/B vssd1 vssd1 vccd1 vccd1 _6797_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_107_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7751__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8535_ _8535_/A _8555_/B vssd1 vssd1 vccd1 vccd1 _8535_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5747_ input50/X _5275_/A _5787_/A1 _5274_/X _5746_/X vssd1 vssd1 vccd1 vccd1 _5829_/C
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7673__A _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8466_ _8466_/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8466_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5678_ _5673_/X _5676_/Y _5677_/Y _6170_/A _5628_/A vssd1 vssd1 vccd1 vccd1 _5678_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__8700__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7503__A2 _5609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7417_ _7378_/X _5328_/A _7683_/C vssd1 vssd1 vccd1 vccd1 _7418_/A sky130_fd_sc_hd__o21ai_1
X_4629_ hold7/X vssd1 vssd1 vccd1 vccd1 _8893_/A sky130_fd_sc_hd__inv_2
X_8397_ _7983_/Y _8299_/X _8396_/X _8304_/X _8518_/B vssd1 vssd1 vccd1 vccd1 _8397_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5193__A _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7348_ _7348_/A vssd1 vssd1 vccd1 vccd1 _7640_/B sky130_fd_sc_hd__buf_6
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7267__B2 _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7279_ _6355_/X _7138_/X _7277_/X _7278_/X vssd1 vssd1 vccd1 vccd1 _7279_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5278__B1 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8216__B1 _8163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8767__A1 _8404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7848__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__B1 _5436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7727__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5087__B _5185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5753__A1 _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6702__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6199__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7258__A1 _6310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8845__C _8845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6646__B _6646_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8207__B1 _8206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4447__A _4760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output515_A _6993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput160 mports_i[38] vssd1 vssd1 vccd1 vccd1 _5988_/A sky130_fd_sc_hd__clkbuf_4
Xinput171 mports_i[48] vssd1 vssd1 vccd1 vccd1 _6287_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__8758__A1 _4930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput182 mports_i[58] vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__clkbuf_2
Xinput193 mports_i[68] vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__buf_2
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7758__A _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7430__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8353__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4980_ _4975_/Y _8455_/B _4976_/Y _4891_/X _4979_/X vssd1 vssd1 vccd1 vccd1 _4981_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__7981__A2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7718__C1 _7749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6650_ _6801_/A _7459_/A _6449_/A vssd1 vssd1 vccd1 vccd1 _6650_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5601_ _5601_/A vssd1 vssd1 vccd1 vccd1 _5601_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_144_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5744__A1 _5518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6581_ _6581_/A _6689_/S vssd1 vssd1 vccd1 vccd1 _6581_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5744__B2 _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8320_ _4933_/X _7862_/Y _4940_/X _7807_/X _8319_/X vssd1 vssd1 vccd1 vccd1 _8320_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_42_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5532_ _5575_/A _5080_/A _5576_/A _5089_/X _5531_/X vssd1 vssd1 vccd1 vccd1 _6697_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__4910__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8251_ _7874_/X _8251_/A2 _7875_/X _8251_/B2 vssd1 vssd1 vccd1 vccd1 _8251_/X sky130_fd_sc_hd__a22o_1
X_5463_ input99/X _8368_/A input37/X _4940_/A vssd1 vssd1 vccd1 vccd1 _5463_/X sky130_fd_sc_hd__o22a_1
Xoutput601 _7114_/X vssd1 vssd1 vccd1 vccd1 sports_o[18] sky130_fd_sc_hd__buf_12
XFILLER_0_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput612 _7119_/X vssd1 vssd1 vccd1 vccd1 sports_o[19] sky130_fd_sc_hd__buf_12
X_7202_ _6867_/A _7023_/X _7201_/X vssd1 vssd1 vccd1 vccd1 _7202_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_111_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput623 _6067_/X vssd1 vssd1 vccd1 vccd1 sports_o[209] sky130_fd_sc_hd__buf_12
X_4414_ _4394_/A _4394_/B _4395_/B vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__a21boi_2
Xoutput634 _6291_/X vssd1 vssd1 vccd1 vccd1 sports_o[219] sky130_fd_sc_hd__buf_12
X_8182_ _8179_/Y _8181_/Y hold12/A vssd1 vssd1 vccd1 vccd1 _8182_/X sky130_fd_sc_hd__o21a_1
Xoutput645 _7137_/X vssd1 vssd1 vccd1 vccd1 sports_o[23] sky130_fd_sc_hd__buf_12
XFILLER_0_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5394_ _5394_/A vssd1 vssd1 vccd1 vccd1 _5394_/Y sky130_fd_sc_hd__inv_2
Xoutput656 _7187_/X vssd1 vssd1 vccd1 vccd1 sports_o[33] sky130_fd_sc_hd__buf_12
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7249__A1 _6263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7133_ _7133_/A vssd1 vssd1 vccd1 vccd1 _7133_/X sky130_fd_sc_hd__buf_1
Xoutput667 _7231_/X vssd1 vssd1 vccd1 vccd1 sports_o[43] sky130_fd_sc_hd__buf_12
Xoutput678 _7281_/X vssd1 vssd1 vccd1 vccd1 sports_o[53] sky130_fd_sc_hd__buf_12
X_4345_ hold26/A hold41/A vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__nor2_4
XANTENNA__6837__A _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput689 _6509_/Y vssd1 vssd1 vccd1 vccd1 sports_o[63] sky130_fd_sc_hd__buf_12
XFILLER_0_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5741__A _5741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8755__C _8755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7064_ _7063_/X _5159_/A _7097_/S vssd1 vssd1 vccd1 vccd1 _7065_/A sky130_fd_sc_hd__mux2_1
X_6015_ _5988_/A _4868_/A _5989_/A _4870_/A _6014_/X vssd1 vssd1 vccd1 vccd1 _6016_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8749__A1 _7903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8749__B2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5680__B1 _5678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7957__C1 _7872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7421__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7966_ _7971_/A1 _5146_/A _7971_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _7966_/Y sky130_fd_sc_hd__o22ai_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5432__B1 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7972__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6917_ _6911_/Y _6467_/X _6912_/Y _6913_/Y _6916_/Y vssd1 vssd1 vccd1 vccd1 _6917_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__5983__A1 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7897_ _7897_/A vssd1 vssd1 vccd1 vccd1 _7897_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6848_ _6848_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7724__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8499__A _8499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6779_ _6547_/A _5842_/A _5782_/A vssd1 vssd1 vccd1 vccd1 _6779_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_91_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8518_ _8518_/A _8518_/B vssd1 vssd1 vccd1 vccd1 _8518_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8449_ _8518_/B _8449_/B vssd1 vssd1 vccd1 vccd1 _8449_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5499__B1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6160__B2 _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5370__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6463__A2 _6876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8959__CLK _8978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7412__A1 _5280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7412__B2 _7638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7297__B _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5974__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6151__B2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7100__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5280__B _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6454__A2 _8188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4465__B2 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6206__A2 _8335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7403__A1 _6576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7820_ _7827_/A _4947_/B _7836_/A _5123_/A _7819_/Y vssd1 vssd1 vccd1 vccd1 _7821_/A
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__8600__B1 _8313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7751_ _7749_/X _7332_/A _7750_/Y vssd1 vssd1 vccd1 vccd1 _7751_/Y sky130_fd_sc_hd__a21oi_2
X_4963_ _4956_/A _8516_/B _4957_/A _4913_/X _4962_/X vssd1 vssd1 vccd1 vccd1 _4963_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6702_ _6801_/A _5562_/X _6450_/A vssd1 vssd1 vccd1 vccd1 _6702_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7682_ _6204_/Y _7361_/X _7679_/X _7680_/Y _7681_/Y vssd1 vssd1 vccd1 vccd1 _7682_/X
+ sky130_fd_sc_hd__a221o_1
X_4894_ _4894_/A vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__inv_6
XANTENNA__7706__A2 _7332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5717__A1 _5159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6633_ _6633_/A _6912_/B vssd1 vssd1 vccd1 vccd1 _6633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4640__A _8264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6564_ _6689_/S _5228_/X _6563_/Y vssd1 vssd1 vccd1 vccd1 _6565_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8303_ _4891_/X _7832_/Y _4894_/A _7798_/X _8302_/X vssd1 vssd1 vccd1 vccd1 _8303_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5515_ _5509_/Y _5514_/Y _6081_/S vssd1 vssd1 vccd1 vccd1 _5516_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6495_ _7767_/A _6495_/B _6497_/B vssd1 vssd1 vccd1 vccd1 _6495_/X sky130_fd_sc_hd__or3_1
XANTENNA__8131__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8234_ _7874_/X _8234_/A2 _7875_/X _8234_/B2 vssd1 vssd1 vccd1 vccd1 _8234_/X sky130_fd_sc_hd__a22o_1
Xoutput420 _8155_/X vssd1 vssd1 vccd1 vccd1 mports_o[26] sky130_fd_sc_hd__buf_12
X_5446_ _7450_/A _5445_/X _6166_/B vssd1 vssd1 vccd1 vccd1 _6668_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6142__A1 _6185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6142__B2 _7683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput431 _8283_/X vssd1 vssd1 vccd1 vccd1 mports_o[36] sky130_fd_sc_hd__buf_12
Xoutput442 _8374_/X vssd1 vssd1 vccd1 vccd1 mports_o[46] sky130_fd_sc_hd__buf_12
Xoutput453 _8498_/X vssd1 vssd1 vccd1 vccd1 mports_o[56] sky130_fd_sc_hd__buf_12
Xoutput464 _8569_/Y vssd1 vssd1 vccd1 vccd1 mports_o[66] sky130_fd_sc_hd__buf_12
XANTENNA__6567__A _6567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8165_ _8165_/A vssd1 vssd1 vccd1 vccd1 _8165_/Y sky130_fd_sc_hd__inv_2
X_5377_ input97/X _4871_/A input35/X _5091_/A vssd1 vssd1 vccd1 vccd1 _5377_/X sky130_fd_sc_hd__o22a_1
Xoutput475 _8619_/X vssd1 vssd1 vccd1 vccd1 mports_o[76] sky130_fd_sc_hd__buf_12
XANTENNA__7890__B2 _7769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput486 _8653_/X vssd1 vssd1 vccd1 vccd1 mports_o[86] sky130_fd_sc_hd__buf_12
Xoutput497 _8687_/X vssd1 vssd1 vccd1 vccd1 mports_o[96] sky130_fd_sc_hd__buf_12
X_7116_ _6671_/B _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7116_/X sky130_fd_sc_hd__a21o_1
X_4328_ _4328_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__nand2_1
X_8096_ _7975_/X _8490_/A _8092_/X _8095_/X vssd1 vssd1 vccd1 vccd1 _8096_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5190__B _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7642__A1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7047_ _7046_/Y _7345_/B _7097_/S vssd1 vssd1 vccd1 vccd1 _7048_/A sky130_fd_sc_hd__mux2_1
XANTENNA__7642__B2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7398__A _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7945__A2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A1 _6031_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _7949_/A vssd1 vssd1 vccd1 vccd1 _7949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5956__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8355__C1 _8518_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5708__A1 _6084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5708__B2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6905__B1 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7337__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4550__A hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5184__A2 _5682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6381__B2 _8257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8658__B1 _8469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8122__A2 _8519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7580__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6684__A2 _5544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6196__B _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4709__B _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4428__C _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6940__A _6940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7149__B1 _7012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6372__A1 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5175__A2 _5161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8113__A2 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _7829_/A _7432_/B _5299_/Y vssd1 vssd1 vccd1 vccd1 _5301_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6280_ _6326_/A1 _5080_/A input9/X _5089_/X _6279_/X vssd1 vssd1 vccd1 vccd1 _6971_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5231_ _5313_/A vssd1 vssd1 vccd1 vccd1 _6689_/S sky130_fd_sc_hd__inv_6
XFILLER_0_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6675__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5291__A _6576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5883__A0 _5880_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5162_ _7304_/A vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__buf_8
X_5093_ _5294_/A _4953_/X _5295_/A _5089_/X _5092_/X vssd1 vssd1 vccd1 vccd1 _5094_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__7710__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5635__B1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8921_ _8921_/A vssd1 vssd1 vccd1 vccd1 _8956_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4989__A2 _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8852_ _8855_/A _8851_/Y _4611_/A vssd1 vssd1 vccd1 vccd1 _8852_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7011__A _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7927__A2 _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7803_ _4566_/A _5197_/X _7803_/B1 _5230_/B _7802_/X vssd1 vssd1 vccd1 vccd1 _7803_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5938__A1 _5274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8783_ _8781_/X _8725_/X _8782_/X _8479_/Y _8759_/Y vssd1 vssd1 vccd1 vccd1 _8783_/X
+ sky130_fd_sc_hd__a32o_1
X_5995_ _8140_/A _5992_/Y _7629_/A vssd1 vssd1 vccd1 vccd1 _5995_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7734_ _7732_/Y _7332_/A _7733_/Y vssd1 vssd1 vccd1 vccd1 _7734_/Y sky130_fd_sc_hd__a21oi_2
X_4946_ _4946_/A vssd1 vssd1 vccd1 vccd1 _4947_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_129_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7665__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7665_ _7665_/A _7691_/B vssd1 vssd1 vccd1 vccd1 _7665_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4877_ _6312_/A _7297_/B vssd1 vssd1 vccd1 vccd1 _6084_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6616_ _6616_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6616_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6363__A1 _6368_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6363__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7596_ _6817_/A _7681_/A _6831_/A _7673_/A _7595_/X vssd1 vssd1 vccd1 vccd1 _7596_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5185__B _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4374__B1 _8239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6996__S _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6547_ _6547_/A _6573_/B vssd1 vssd1 vccd1 vccd1 _6547_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8104__A2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7681__A _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6478_ _5000_/X _6467_/X _6468_/X _6477_/X _6450_/X vssd1 vssd1 vccd1 vccd1 _6478_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8217_ _4312_/B _5299_/B _8222_/B1 _5171_/B _8216_/X vssd1 vssd1 vccd1 vccd1 _8217_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5429_ _6133_/B _5423_/X _5427_/X _6233_/B _5428_/X vssd1 vssd1 vccd1 vccd1 _5429_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8148_ _8148_/A1 _6544_/B _8142_/A _4518_/A _8147_/X vssd1 vssd1 vccd1 vccd1 _8148_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4529__B _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8812__B1 _8148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7615__B2 _7361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8079_ _8483_/A _7954_/X _8480_/A _7826_/X _7872_/X vssd1 vssd1 vccd1 vccd1 _8079_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7091__A2 _7023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7379__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7918__A2 _7876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8040__A1 _8036_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5929__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8040__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5929__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8591__A2 _8295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7856__A _7856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6760__A _6760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8343__A2 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6354__A1 _6357_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6354__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6919__B _7678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6657__A2 _6933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output428_A _8254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5093__A1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5093__B2 _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7766__A _8709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4800_/A _4800_/B vssd1 vssd1 vccd1 vccd1 _8875_/A sky130_fd_sc_hd__nand2_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5396__A2 _5094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5780_ _5780_/A vssd1 vssd1 vccd1 vccd1 _5780_/X sky130_fd_sc_hd__buf_8
XFILLER_0_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7790__B1 _7311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _4731_/A _8481_/S vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__nand2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7450_ _7450_/A _7638_/B vssd1 vssd1 vccd1 vccd1 _7450_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4662_ _4662_/A _7737_/B _4662_/C vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__or3_1
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6401_ _6401_/A1 _4930_/X input16/X _4933_/X _6400_/X vssd1 vssd1 vccd1 vccd1 _7756_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6896__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7381_ _7686_/A vssd1 vssd1 vccd1 vccd1 _7542_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4593_ _8845_/A _8759_/A vssd1 vssd1 vccd1 vccd1 _4593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6332_ input73/X _8579_/C _6336_/A1 _8713_/C _6331_/X vssd1 vssd1 vccd1 vccd1 _6333_/A
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7845__A1 _7840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6263_ _6253_/A _8523_/B input6/X _4933_/A _6262_/X vssd1 vssd1 vccd1 vccd1 _6263_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__7845__B2 _7835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4659__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8002_ _8002_/A vssd1 vssd1 vccd1 vccd1 _8002_/Y sky130_fd_sc_hd__inv_2
X_5214_ _5159_/B _5211_/A _5209_/X _6402_/A _5213_/X vssd1 vssd1 vccd1 vccd1 _5214_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6194_ _6229_/A2 _8709_/B input66/X _5091_/X vssd1 vssd1 vccd1 vccd1 _6194_/X sky130_fd_sc_hd__o22a_1
X_5145_ _5145_/A vssd1 vssd1 vccd1 vccd1 _5146_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__7519__A1_N _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _6488_/A _7629_/B _5171_/B _5075_/Y vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5084__A1 _5139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5084__B2 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8904_ _8904_/A _8904_/B vssd1 vssd1 vccd1 vccd1 _8904_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6775__A1_N _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8022__B2 _6500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8835_ _4607_/A _8820_/B _8829_/S vssd1 vssd1 vccd1 vccd1 _8835_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6033__A0 _6030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6580__A _6580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5387__A2 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8766_ _8764_/X _8725_/X _8765_/X _8415_/Y _8759_/Y vssd1 vssd1 vccd1 vccd1 _8766_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5978_ _5965_/A _5080_/A _5966_/A _5089_/X _5977_/X vssd1 vssd1 vccd1 vccd1 _6028_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_149_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7717_ _7717_/A vssd1 vssd1 vccd1 vccd1 _7717_/X sky130_fd_sc_hd__buf_1
X_4929_ _4929_/A vssd1 vssd1 vccd1 vccd1 _8523_/B sky130_fd_sc_hd__buf_12
XFILLER_0_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8697_ _8275_/X _7629_/B hold41/A _8696_/A _8696_/Y vssd1 vssd1 vccd1 vccd1 _8698_/A
+ sky130_fd_sc_hd__a41o_1
XANTENNA__8325__A2 _7878_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5196__A _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6336__A1 _6336_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7648_ _7694_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7648_/X sky130_fd_sc_hd__or2_1
XANTENNA__6336__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7533__B1 _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6887__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7579_ _7378_/X _5824_/X _7683_/C vssd1 vssd1 vccd1 vccd1 _7581_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5924__A _5924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4898__B2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8300__A _8455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8089__B2 _6080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6639__A2 _6467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5847__B1 _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A2 _7413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8446__S _8512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8797__C1 _8788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8955__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6272__B1 _6286_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4822__A1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8013__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5378__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6327__A1 _6326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8721__C1 _8820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5550__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5838__B1 _5805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8252__A1 _8252_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8252__B2 _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6263__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6950_ _8574_/B _6947_/X _6948_/Y _6949_/X vssd1 vssd1 vccd1 vccd1 _6950_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_89_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8004__A1 _8011_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5901_ _5895_/X _5960_/B _6926_/A vssd1 vssd1 vccd1 vccd1 _5901_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6881_ _6881_/A vssd1 vssd1 vccd1 vccd1 _6882_/A sky130_fd_sc_hd__inv_2
XFILLER_0_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6015__B1 _5989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8620_ _8352_/A _8581_/A _7916_/Y _8583_/A vssd1 vssd1 vccd1 vccd1 _8620_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _6780_/A _5832_/B vssd1 vssd1 vccd1 vccd1 _5832_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4913__A _4913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5369__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7763__B1 _4481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8551_ _8551_/A _8755_/B vssd1 vssd1 vccd1 vccd1 _8551_/Y sky130_fd_sc_hd__nand2_1
X_5763_ _6084_/B _7551_/A _5755_/X _5715_/B _5762_/Y vssd1 vssd1 vccd1 vccd1 _5763_/X
+ sky130_fd_sc_hd__a221o_1
X_7502_ _7590_/A _7494_/Y _8759_/A _5645_/Y _7501_/X vssd1 vssd1 vccd1 vccd1 _7502_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4714_ _4714_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6318__A1 _6336_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8482_ _8482_/A _8482_/B vssd1 vssd1 vccd1 vccd1 _8482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6318__B2 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7515__B1 _7385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5694_ _5909_/B _5600_/Y _5693_/X _5997_/B _6234_/B vssd1 vssd1 vccd1 vccd1 _5694_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7433_ _5094_/Y _8578_/B _8919_/A vssd1 vssd1 vccd1 vccd1 _7433_/Y sky130_fd_sc_hd__a21oi_1
X_4645_ _4800_/B _4934_/A _4810_/B _4937_/A vssd1 vssd1 vccd1 vccd1 _4645_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7364_ _7364_/A vssd1 vssd1 vccd1 vccd1 _7638_/B sky130_fd_sc_hd__inv_6
X_4576_ _8584_/A vssd1 vssd1 vccd1 vccd1 _5193_/A sky130_fd_sc_hd__clkinv_8
XANTENNA__5541__A2 _7629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6315_ hold26/A _6315_/B vssd1 vssd1 vccd1 vccd1 _6315_/Y sky130_fd_sc_hd__nand2_1
X_7295_ _7294_/Y _7756_/B _7295_/S vssd1 vssd1 vccd1 vccd1 _7296_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_97_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6246_ _6128_/B _7707_/D _6245_/X vssd1 vssd1 vccd1 vccd1 _6246_/X sky130_fd_sc_hd__o21a_1
XANTENNA__8266__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6575__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6177_ _6173_/Y _6176_/Y _8150_/A vssd1 vssd1 vccd1 vccd1 _6177_/X sky130_fd_sc_hd__mux2_1
X_5128_ _5128_/A vssd1 vssd1 vccd1 vccd1 _5128_/Y sky130_fd_sc_hd__inv_2
XANTENNA__8243__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8243__B2 _8252_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5057__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _7037_/B sky130_fd_sc_hd__inv_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8546__A2 _8175_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8818_ _8157_/X _8725_/X _8815_/Y _8817_/X vssd1 vssd1 vccd1 vccd1 _8818_/X sky130_fd_sc_hd__o22a_2
XFILLER_0_67_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8749_ _7903_/Y _8711_/X _8362_/X _8803_/B _8820_/B vssd1 vssd1 vccd1 vccd1 _8749_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6309__A1 _6309_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6309__B2 _4917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8703__C1 _8621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7853__B _7859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5654__A _6743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5532__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7809__A1 _7814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7809__B2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5296__A1 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5296__B2 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput320 sports_i[59] vssd1 vssd1 vccd1 vccd1 _8124_/A sky130_fd_sc_hd__clkbuf_1
Xinput331 sports_i[69] vssd1 vssd1 vccd1 vccd1 _7790_/B2 sky130_fd_sc_hd__buf_2
Xinput342 sports_i[79] vssd1 vssd1 vccd1 vccd1 _7944_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__8234__A1 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput353 sports_i[89] vssd1 vssd1 vccd1 vccd1 _8080_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__8234__B2 _8234_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5048__A1 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput364 sports_i[99] vssd1 vssd1 vccd1 vccd1 _8235_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4717__B hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5048__B2 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6245__B1 _7242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5599__A2 _4885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6796__A1 _6788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7993__B1 _7998_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6796__B2 _6801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8537__A2 _8820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5829__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6548__A1 _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5771__A2 _4934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7255__S _7295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8170__B1 _8169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4430_ _4430_/A vssd1 vssd1 vccd1 vccd1 _4430_/Y sky130_fd_sc_hd__inv_2
XANTENNA_2 _6285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4361_ _8938_/S vssd1 vssd1 vccd1 vccd1 _8936_/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6100_ _6136_/A1 _5192_/A input62/X _5193_/A vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__o22a_1
XANTENNA__8473__A1 _8068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7080_ _5323_/A _7023_/X _7079_/X vssd1 vssd1 vccd1 vccd1 _7080_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_120_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4292_ _7683_/B _4658_/A vssd1 vssd1 vccd1 vccd1 _4393_/B sky130_fd_sc_hd__nand2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5287__A1 _6284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6031_ _6031_/A1 _8271_/B input58/X _4917_/A vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__o22a_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7028__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8225__A1 _7761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8225__B2 _8234_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5039__A1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5039__B2 _4917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8776__A2 _8806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7982_ _7985_/A1 _5780_/X _7985_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7982_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__7984__B1 _7983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6933_ _6933_/A _7686_/B vssd1 vssd1 vccd1 vccd1 _6933_/Y sky130_fd_sc_hd__nor2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6539__A1 _7383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6864_ _7630_/A _6475_/X _5975_/X _6851_/B vssd1 vssd1 vccd1 vccd1 _6864_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6539__B2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8603_ _7825_/X _8583_/X _7832_/Y _8581_/X _8685_/B vssd1 vssd1 vccd1 vccd1 _8603_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5815_ _5751_/X _5814_/X _6780_/A vssd1 vssd1 vccd1 vccd1 _5816_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6795_ _6792_/X _6933_/A _6968_/A _6794_/X vssd1 vssd1 vccd1 vccd1 _6795_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_123_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8534_ _8157_/X _8323_/X _8532_/X _8533_/Y vssd1 vssd1 vccd1 vccd1 _8534_/X sky130_fd_sc_hd__a22o_2
X_5746_ _5129_/A _5788_/A1 _5130_/A _5788_/B1 vssd1 vssd1 vccd1 vccd1 _5746_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4970__B1 _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8465_ _8445_/Y _8464_/Y hold26/A vssd1 vssd1 vccd1 vccd1 _8466_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5677_ _5660_/A _5845_/B _6386_/S vssd1 vssd1 vccd1 vccd1 _5677_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7416_ _5247_/X _7361_/X _7414_/X _7754_/A _7415_/Y vssd1 vssd1 vccd1 vccd1 _7416_/X
+ sky130_fd_sc_hd__a221o_1
X_4628_ _8953_/D hold7/X vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8396_ _8755_/B _8395_/X _8713_/C _8359_/A vssd1 vssd1 vccd1 vccd1 _8396_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7347_ _7347_/A vssd1 vssd1 vccd1 vccd1 _7348_/A sky130_fd_sc_hd__inv_6
X_4559_ _8181_/A hold12/A vssd1 vssd1 vccd1 vccd1 _5229_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7267__A2 _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7278_ _7278_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7278_/X sky130_fd_sc_hd__and2_1
XANTENNA__5278__A1 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6229_ _8713_/C _6229_/A2 _8579_/C input66/X vssd1 vssd1 vccd1 vccd1 _6229_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__8216__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8216__B2 _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4537__B _8716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8767__A2 _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6778__A1 _5772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6778__B2 _6512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7848__B _7859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5986__C1 _5985_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5450__A1 _5435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5450__B2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6950__A1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5384__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6702__A1 _6801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6199__B _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8970__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7258__A2 _7026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5269__A1 _6304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8207__A1 _8203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8207__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput150 mports_i[29] vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__clkbuf_4
Xinput161 mports_i[39] vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__clkbuf_4
Xinput172 mports_i[49] vssd1 vssd1 vccd1 vccd1 _6299_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__8758__A2 _8345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput183 mports_i[59] vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output410_A _8027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput194 mports_i[69] vssd1 vssd1 vccd1 vccd1 _5326_/B1 sky130_fd_sc_hd__clkbuf_2
XANTENNA_output508_A _6964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7966__B1 _7971_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7758__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7430__A2 _7681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6662__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4463__A _5780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7194__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7774__A _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ _5666_/C vssd1 vssd1 vccd1 vccd1 _5600_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_156_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6580_ _6580_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6580_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5744__A2 _5111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5531_ _5587_/A1 _8709_/B input41/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_143_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5294__A _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8250_ _8247_/Y _7826_/A _8249_/X _7768_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8250_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5462_ _5462_/A vssd1 vssd1 vccd1 vccd1 _5462_/X sky130_fd_sc_hd__buf_1
XANTENNA__8694__A1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8694__B2 _8590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput602 _5528_/X vssd1 vssd1 vccd1 vccd1 sports_o[190] sky130_fd_sc_hd__buf_12
X_7201_ _6028_/A _7004_/X _7630_/A _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7201_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput613 _7025_/X vssd1 vssd1 vccd1 vccd1 sports_o[1] sky130_fd_sc_hd__buf_12
X_4413_ _4413_/A _6434_/B vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__nand2_1
Xoutput624 _7125_/X vssd1 vssd1 vccd1 vccd1 sports_o[20] sky130_fd_sc_hd__buf_12
X_8181_ _8181_/A _8194_/B vssd1 vssd1 vccd1 vccd1 _8181_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__8809__S _8824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5393_ _6166_/B _5301_/B _5392_/X vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__o21ai_1
Xoutput635 _7129_/X vssd1 vssd1 vccd1 vccd1 sports_o[21] sky130_fd_sc_hd__buf_12
Xoutput646 _7143_/X vssd1 vssd1 vccd1 vccd1 sports_o[24] sky130_fd_sc_hd__buf_12
XFILLER_0_10_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput657 _7191_/X vssd1 vssd1 vccd1 vccd1 sports_o[34] sky130_fd_sc_hd__buf_12
X_7132_ _7131_/X _5645_/A _7175_/S vssd1 vssd1 vccd1 vccd1 _7133_/A sky130_fd_sc_hd__mux2_1
Xoutput668 _7236_/X vssd1 vssd1 vccd1 vccd1 sports_o[44] sky130_fd_sc_hd__buf_12
X_4344_ _5130_/A _4823_/B vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__nand2_1
Xoutput679 _7286_/X vssd1 vssd1 vccd1 vccd1 sports_o[54] sky130_fd_sc_hd__buf_12
XANTENNA__6837__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7063_ _5196_/A _7023_/X _7062_/X vssd1 vssd1 vccd1 vccd1 _7063_/X sky130_fd_sc_hd__o21a_1
X_6014_ _6061_/A1 _5090_/A input59/X _4874_/A vssd1 vssd1 vccd1 vccd1 _6014_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5680__A1 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8749__A2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5680__B2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7957__B1 _7956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7421__A2 _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7668__B _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7965_ _7962_/Y _7013_/A _7963_/Y _5117_/A _7964_/Y vssd1 vssd1 vccd1 vccd1 _8375_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5432__A1 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _6102_/A _6801_/A _6924_/A _6915_/Y _6450_/A vssd1 vssd1 vccd1 vccd1 _6916_/Y
+ sky130_fd_sc_hd__o221ai_4
X_7896_ _7896_/A vssd1 vssd1 vccd1 vccd1 _7896_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_134_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7185__A1 _6828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6847_ _6847_/A vssd1 vssd1 vccd1 vccd1 _6848_/A sky130_fd_sc_hd__inv_2
XFILLER_0_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8382__B1 _8349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6778_ _5772_/X _6908_/B _5778_/A _6512_/X _6777_/X vssd1 vssd1 vccd1 vccd1 _6778_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8499__B _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6932__B2 _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8517_ _8515_/Y _8516_/Y _8904_/A vssd1 vssd1 vccd1 vccd1 _8518_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ _6780_/B _5692_/X _6837_/A vssd1 vssd1 vccd1 vccd1 _6755_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8448_ _8039_/A _8259_/A _8429_/Y _8447_/X vssd1 vssd1 vccd1 vccd1 _8449_/B sky130_fd_sc_hd__o22a_1
XANTENNA__5499__A1 _5557_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5499__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6696__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8379_ _8441_/B _7912_/Y _8435_/A _8759_/B vssd1 vssd1 vccd1 vccd1 _8379_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6160__A2 _4891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5932__A _5932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6999__B2 _6989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__A1 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7859__A _8194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7412__A2 _7668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8125__B1 _8132_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8676__A1 _8523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6151__A2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7100__A1 _6634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6454__A3 _6544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6483__A1_N _6854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4465__A2 _4318_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7769__A _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7939__B1 _7944_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8600__A1 _8309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7488__B _7680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7403__A2 _7532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8600__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5414__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4962_ input81/X _8716_/B input18/X _4917_/X vssd1 vssd1 vccd1 vccd1 _4962_/X sky130_fd_sc_hd__o22a_1
X_7750_ _7756_/A _7750_/B vssd1 vssd1 vccd1 vccd1 _7750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6701_ _6924_/A _6701_/B vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7681_ _7681_/A _7681_/B vssd1 vssd1 vccd1 vccd1 _7681_/Y sky130_fd_sc_hd__nor2_1
X_4893_ _4893_/A vssd1 vssd1 vccd1 vccd1 _8713_/C sky130_fd_sc_hd__buf_8
XFILLER_0_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6632_ _6632_/A _6933_/A vssd1 vssd1 vccd1 vccd1 _6632_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4921__A _6181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5717__A2 _6743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6563_ _6563_/A _6689_/S vssd1 vssd1 vccd1 vccd1 _6563_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__8116__B1 _8119_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6390__A2 _6402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8302_ _7765_/X hold26/A _8513_/B vssd1 vssd1 vccd1 vccd1 _8302_/X sky130_fd_sc_hd__a21o_1
X_5514_ _6080_/A _7120_/A vssd1 vssd1 vccd1 vccd1 _5514_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8667__A1 _8490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6494_ _6513_/A vssd1 vssd1 vccd1 vccd1 _6495_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8233_ _7772_/X _8230_/Y _8232_/X _7768_/X _7872_/A vssd1 vssd1 vccd1 vccd1 _8233_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6678__B1 _6436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5445_ _5537_/A _5444_/Y _6081_/S vssd1 vssd1 vccd1 vccd1 _5445_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput410 _8027_/X vssd1 vssd1 vccd1 vccd1 mports_o[17] sky130_fd_sc_hd__buf_12
XANTENNA__6142__A2 _8924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput421 _8177_/X vssd1 vssd1 vccd1 vccd1 mports_o[27] sky130_fd_sc_hd__buf_12
Xoutput432 _8288_/X vssd1 vssd1 vccd1 vccd1 mports_o[37] sky130_fd_sc_hd__buf_12
XANTENNA__5752__A _6166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput443 _8389_/X vssd1 vssd1 vccd1 vccd1 mports_o[47] sky130_fd_sc_hd__buf_12
XFILLER_0_100_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8164_ _8175_/A1 _6456_/B _8159_/Y _8161_/Y _8163_/Y vssd1 vssd1 vccd1 vccd1 _8165_/A
+ sky130_fd_sc_hd__o221ai_2
Xoutput454 _8509_/X vssd1 vssd1 vccd1 vccd1 mports_o[57] sky130_fd_sc_hd__buf_12
XANTENNA__7890__A2 _6500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5376_ _5348_/Y _6402_/A _5355_/Y _5356_/X _5375_/X vssd1 vssd1 vccd1 vccd1 _5376_/X
+ sky130_fd_sc_hd__a41o_2
Xoutput465 _8573_/X vssd1 vssd1 vccd1 vccd1 mports_o[67] sky130_fd_sc_hd__buf_12
XANTENNA__6567__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput476 _8623_/X vssd1 vssd1 vccd1 vccd1 mports_o[77] sky130_fd_sc_hd__buf_12
Xoutput487 _8657_/X vssd1 vssd1 vccd1 vccd1 mports_o[87] sky130_fd_sc_hd__buf_12
X_7115_ _7115_/A _7246_/B vssd1 vssd1 vccd1 vccd1 _7115_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput498 _8691_/X vssd1 vssd1 vccd1 vccd1 mports_o[97] sky130_fd_sc_hd__buf_12
X_4327_ _4337_/A _7818_/A vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__nand2_1
X_8095_ _7777_/A _8516_/A _7792_/A vssd1 vssd1 vccd1 vccd1 _8095_/X sky130_fd_sc_hd__o21ba_1
X_7046_ _7046_/A vssd1 vssd1 vccd1 vccd1 _7046_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7642__A2 _7389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8782__B _8782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5653__A1 _5661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _7948_/A vssd1 vssd1 vccd1 vccd1 _7948_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5956__A2 _8368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7158__A1 _7551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7879_ _7777_/X _7878_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _7879_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__7158__B2 _7088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5708__A2 _6727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6905__A1 _6058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6905__B2 _6095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6381__A2 _8444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8658__A1 _8464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8658__B2 _8583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6758__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6477__B _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5892__A1 _6906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4709__C _7272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7633__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7397__A1 _6566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7397__B2 _7326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7149__A1 _6727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8897__A1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8649__A1 _8433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7857__C1 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7321__A1 _4963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5230_ _7874_/A _5230_/B vssd1 vssd1 vccd1 vccd1 _5313_/A sky130_fd_sc_hd__nor2_2
XANTENNA__5883__A1 _6801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5161_ input26/X _4896_/A input88/X _4893_/A _5160_/X vssd1 vssd1 vccd1 vccd1 _5161_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7624__A2 _7660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5092_ input95/X _8709_/B input32/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5635__A1 _5635_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold10_A hold10/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5635__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6832__B1 _6824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8920_ _4761_/A hold36/X _8922_/A vssd1 vssd1 vccd1 vccd1 _8921_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4916__A _5193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8851_ _8861_/A _8856_/B vssd1 vssd1 vccd1 vccd1 _8851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7388__A1 _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7388__B2 _7694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7802_ _7874_/A _7802_/A2 _8174_/A _4326_/B vssd1 vssd1 vccd1 vccd1 _7802_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5938__A2 _5962_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5994_ _5994_/A vssd1 vssd1 vccd1 vccd1 _7629_/A sky130_fd_sc_hd__inv_2
X_8782_ _8782_/A _8782_/B vssd1 vssd1 vccd1 vccd1 _8782_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6060__A1 _8842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7733_ _7756_/A _7733_/B vssd1 vssd1 vccd1 vccd1 _7733_/Y sky130_fd_sc_hd__nor2_1
X_4945_ _5741_/B vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__inv_2
XFILLER_0_115_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4651__A hold44/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4876_ input1/X _5080_/A _4888_/A _4870_/X _4875_/X vssd1 vssd1 vccd1 vccd1 _4876_/X
+ sky130_fd_sc_hd__o221a_2
X_7664_ _7701_/A _6094_/X _6264_/X vssd1 vssd1 vccd1 vccd1 _7665_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6615_ _6608_/X _6609_/Y _6610_/X _6614_/X vssd1 vssd1 vccd1 vccd1 _6615_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_28_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4370__B _4800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7595_ _7592_/Y _7593_/X _5864_/A _7680_/B _7594_/Y vssd1 vssd1 vccd1 vccd1 _7595_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6363__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8949__CLK _8979_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6546_ _6550_/A _6017_/A _7299_/A _6526_/A vssd1 vssd1 vccd1 vccd1 _6573_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6477_ _6477_/A _6899_/B vssd1 vssd1 vccd1 vccd1 _6477_/X sky130_fd_sc_hd__and2_1
XANTENNA__6578__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5482__A _6481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8216_ _6965_/A _8221_/A2 _8163_/A _4478_/B vssd1 vssd1 vccd1 vccd1 _8216_/X sky130_fd_sc_hd__a22o_1
X_5428_ _6634_/A _5845_/B _6386_/S vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5874__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5359_ _5359_/A _5359_/B vssd1 vssd1 vccd1 vccd1 _6926_/A sky130_fd_sc_hd__nor2_4
X_8147_ _8151_/A _8188_/S _8189_/B _8146_/Y vssd1 vssd1 vccd1 vccd1 _8147_/X sky130_fd_sc_hd__a211o_1
XANTENNA__8812__A1 _8145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8078_ _8071_/Y _7769_/A _8072_/Y _6500_/A _8077_/Y vssd1 vssd1 vccd1 vccd1 _8480_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7615__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8812__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5626__A1 _5640_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5626__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7029_ _4992_/X _7026_/X _7027_/X _7028_/X vssd1 vssd1 vccd1 vccd1 _7029_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6823__B1 _8574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__B _8150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7379__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8040__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5929__A2 _8271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6760__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8328__B1 _8323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4561__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6354__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7872__A _7872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5314__B1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6814__B1 _7707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5093__A2 _4953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7766__B _8480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8319__B1 _8759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7790__A1 _7874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7790__B2 _7790_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4730_ _4759_/A _4759_/B _4760_/A vssd1 vssd1 vccd1 vccd1 _4750_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__4471__A _7852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ _4661_/A vssd1 vssd1 vccd1 vccd1 _4662_/C sky130_fd_sc_hd__clkinv_4
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6400_ _6400_/A1 _8706_/B input79/X _4940_/X vssd1 vssd1 vccd1 vccd1 _6400_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7380_ _7380_/A _7619_/B vssd1 vssd1 vccd1 vccd1 _7380_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5553__B1 _6281_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4592_ hold20/X vssd1 vssd1 vccd1 vccd1 _8759_/A sky130_fd_sc_hd__inv_12
XFILLER_0_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6331_ _8444_/A _6337_/B1 _8257_/C input10/X vssd1 vssd1 vccd1 vccd1 _6331_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6262_ _6262_/A1 _8368_/A input69/X _4940_/A vssd1 vssd1 vccd1 vccd1 _6262_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_40_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7845__A2 _7876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8402__A1_N _8555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8001_ _7975_/X _8400_/A _7997_/X _8000_/X vssd1 vssd1 vccd1 vccd1 _8001_/X sky130_fd_sc_hd__a22o_4
X_5213_ _6535_/A _8574_/B _5359_/B vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__and3_2
X_6193_ _6115_/Y _6152_/Y _6281_/S vssd1 vssd1 vccd1 vccd1 _7680_/A sky130_fd_sc_hd__mux2_1
X_5144_ _5999_/B vssd1 vssd1 vccd1 vccd1 _5909_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5075_ _6304_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _5075_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__7022__A _7089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5084__A2 _5080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6281__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8903_ _8903_/A _8903_/B vssd1 vssd1 vccd1 vccd1 _8975_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8834_ _8226_/X _8725_/X _8831_/Y _8833_/X vssd1 vssd1 vccd1 vccd1 _8834_/X sky130_fd_sc_hd__o22a_2
XANTENNA__8022__A2 _7769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6033__A1 _6867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7230__A0 _7229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8765_ _8782_/A _8765_/B vssd1 vssd1 vccd1 vccd1 _8765_/X sky130_fd_sc_hd__or2_1
XANTENNA__6580__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5977_ _6031_/A1 _8709_/B input58/X _5091_/X vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__o22a_1
XANTENNA__7781__A1 _7777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7716_ _7715_/X _6263_/X _7741_/S vssd1 vssd1 vccd1 vccd1 _7717_/A sky130_fd_sc_hd__mux2_1
X_4928_ _5111_/A vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__buf_8
X_8696_ _8696_/A _8696_/B vssd1 vssd1 vccd1 vccd1 _8696_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7688__A1_N _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7647_ _6905_/X _7619_/B _7643_/X _7645_/Y _7646_/Y vssd1 vssd1 vccd1 vccd1 _7647_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6336__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4859_ _4859_/A _8933_/B vssd1 vssd1 vccd1 vccd1 _4860_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7692__A _7701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5544__B1 _5511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7578_ _6788_/B _7696_/B _7576_/X _7326_/A _7577_/Y vssd1 vssd1 vccd1 vccd1 _7578_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4898__A2 _8550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5924__B _6626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8089__A2 _6513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6529_ _6882_/B vssd1 vssd1 vccd1 vccd1 _6871_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5847__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5940__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7049__B1 _7138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6755__B _6851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8797__B1 _8091_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8028__A _8028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6272__A1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6272__B2 _8713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8549__B1 _4870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8013__A2 _8012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6771__A _6771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7221__A0 _7220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4291__A _7510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8721__B1 _8313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5550__A3 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5838__A1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5838__B2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output440_A _8350_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8252__A2 _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output705_A _6692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6263__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5996__S _6711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5900_ _8842_/B _5898_/Y _7607_/B vssd1 vssd1 vccd1 vccd1 _5960_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6880_ _6867_/A _5197_/X _7707_/B _6063_/A vssd1 vssd1 vccd1 vccd1 _6881_/A sky130_fd_sc_hd__a22o_1
XANTENNA__6015__A1 _5988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7212__A0 _7211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6015__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5831_ _6470_/B _5813_/Y _5830_/Y vssd1 vssd1 vccd1 vccd1 _5832_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__7763__A1 _4318_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7763__B2 _7316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8550_ _8550_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8551_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5762_ _5762_/A _5762_/B vssd1 vssd1 vccd1 vccd1 _5762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7501_ _5566_/Y _7361_/X _7499_/X _7723_/B _7500_/X vssd1 vssd1 vccd1 vccd1 _7501_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4713_ _4713_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__nor2_1
XANTENNA__6318__A2 _8310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8481_ _8480_/Y _8458_/Y _8481_/S vssd1 vssd1 vccd1 vccd1 _8482_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5693_ _5608_/X _5692_/X _6166_/B vssd1 vssd1 vccd1 vccd1 _5693_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7716__S _7741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4644_ _8574_/A vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__inv_2
X_7432_ _7532_/A _7432_/B vssd1 vssd1 vccd1 vccd1 _7432_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_142_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4575_ _8336_/S _4788_/C vssd1 vssd1 vccd1 vccd1 _8584_/A sky130_fd_sc_hd__nor2_4
X_7363_ _7363_/A vssd1 vssd1 vccd1 vccd1 _7680_/B sky130_fd_sc_hd__buf_6
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5541__A3 _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6314_ _8512_/S _6314_/B vssd1 vssd1 vccd1 vccd1 _6314_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7294_ _7294_/A vssd1 vssd1 vccd1 vccd1 _7294_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6245_ _6241_/X _6234_/B _7242_/A _5128_/A _6356_/S vssd1 vssd1 vccd1 vccd1 _6245_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6856__A _6856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6176_ _6212_/B _6868_/B vssd1 vssd1 vccd1 vccd1 _6176_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6575__B _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5127_ _5100_/X _6402_/A _5108_/X _5109_/X _5126_/X vssd1 vssd1 vccd1 vccd1 _5127_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__4376__A _5827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5058_ _5051_/X _7629_/B _5171_/B _5057_/Y vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__a31o_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8282__S _8572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6591__A _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8817_ _8817_/A _8833_/B vssd1 vssd1 vccd1 vccd1 _8817_/X sky130_fd_sc_hd__and2_1
XANTENNA__5214__C1 _5213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4823__B _4823_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5765__B1 _5519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8748_ _8748_/A vssd1 vssd1 vccd1 vccd1 _8748_/X sky130_fd_sc_hd__buf_1
XANTENNA__4568__B2 _4601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6309__A2 _8716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8679_ _8538_/X _8685_/B _8686_/B vssd1 vssd1 vccd1 vccd1 _8679_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__7506__A1 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8703__B1 _8249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5935__A _6024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8311__A _8311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6714__C1 _7000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7809__A2 _5171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7565__A1_N _7700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5670__A _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5296__A2 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6493__A1 _7345_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7690__B1 _7683_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput310 sports_i[4] vssd1 vssd1 vccd1 vccd1 _7829_/B sky130_fd_sc_hd__buf_2
Xinput321 sports_i[5] vssd1 vssd1 vccd1 vccd1 _7858_/B sky130_fd_sc_hd__buf_2
Xinput332 sports_i[6] vssd1 vssd1 vccd1 vccd1 _7864_/A sky130_fd_sc_hd__buf_1
Xinput343 sports_i[7] vssd1 vssd1 vccd1 vccd1 _7883_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__8234__A2 _8234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput354 sports_i[8] vssd1 vssd1 vccd1 vccd1 _7896_/A sky130_fd_sc_hd__buf_1
Xinput365 sports_i[9] vssd1 vssd1 vccd1 vccd1 _7909_/A sky130_fd_sc_hd__buf_1
XANTENNA__5048__A2 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6245__A1 _6241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6245__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7442__B1 _7440_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7993__A1 _7998_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6796__A2 _5197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7993__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6705__S _6837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5829__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6006__A _6006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5220__A2 _6233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8170__A1 _7768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8170__B2 _7826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _7729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ _4406_/A _4360_/B vssd1 vssd1 vccd1 vccd1 _8938_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8875__B _8875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8367__S _8496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8473__A2 _8567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6676__A _7767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4291_ _7510_/B vssd1 vssd1 vccd1 vccd1 _7683_/B sky130_fd_sc_hd__clkinv_4
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7130__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _5096_/A _7637_/B _6027_/X _5715_/B _6029_/Y vssd1 vssd1 vccd1 vccd1 _6030_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6484__A1 _6899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5287__A2 _6578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6395__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8225__A2 _8234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5039__A2 _8271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7433__B1 _8919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7981_ _7976_/Y _6513_/A _7977_/Y _6080_/A _7980_/Y vssd1 vssd1 vccd1 vccd1 _8394_/A
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__7984__A1 _8394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7984__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6932_ _6931_/Y _6475_/X _6161_/Y _6851_/B vssd1 vssd1 vccd1 vccd1 _6932_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4924__A _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7300__A _7686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6863_ _6856_/Y _6450_/X _6859_/Y _6861_/Y _6862_/X vssd1 vssd1 vccd1 vccd1 _6863_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__7197__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6539__A2 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7736__A1 _4793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8602_ _8320_/X _8577_/X _8600_/X _8601_/X vssd1 vssd1 vccd1 vccd1 _8602_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5747__B1 _5787_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5814_ _5904_/A _5813_/Y _6081_/S vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_146_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6794_ _6854_/A _7575_/B _5879_/A _6913_/B vssd1 vssd1 vccd1 vccd1 _6794_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8533_ _8175_/Y _8518_/B _8572_/S vssd1 vssd1 vccd1 vccd1 _8533_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5745_ _5745_/A vssd1 vssd1 vccd1 vccd1 _5745_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4970__A1 _4975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8464_ _8464_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8464_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4970__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5676_ _8189_/A _5675_/Y _6133_/B vssd1 vssd1 vccd1 vccd1 _5676_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7415_ _7681_/A _7415_/B vssd1 vssd1 vccd1 vccd1 _7415_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_142_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4627_ _4627_/A _4662_/A vssd1 vssd1 vccd1 vccd1 _8953_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_142_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8395_ _8394_/Y _8358_/Y _8512_/S vssd1 vssd1 vccd1 vccd1 _8395_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4558_ _4611_/B vssd1 vssd1 vccd1 vccd1 _7778_/B sky130_fd_sc_hd__inv_2
X_7346_ _7344_/Y _7332_/A _7345_/Y vssd1 vssd1 vccd1 vccd1 _7346_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_130_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7277_ _6349_/X _7059_/X _7061_/X vssd1 vssd1 vccd1 vccd1 _7277_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ hold36/A hold15/A vssd1 vssd1 vccd1 vccd1 _4871_/A sky130_fd_sc_hd__nand2_8
XANTENNA__5490__A _5490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7181__S _7249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5278__A2 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6228_ input4/X vssd1 vssd1 vccd1 vccd1 _6228_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4818__B _4818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6159_ _4893_/A _6174_/A1 _4896_/A input64/X vssd1 vssd1 vccd1 vccd1 _6159_/Y sky130_fd_sc_hd__a22oi_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6778__A2 _6908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5986__B1 _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__A2 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7727__A1 _6317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7188__C1 _7089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7727__B2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5202__A2 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5665__A _6079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4961__A1 _6440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4961__B2 _5128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8152__B2 _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6163__B1 _6182_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6702__A2 _5562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6199__C _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5269__A2 _6576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8207__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput140 mports_i[225] vssd1 vssd1 vccd1 vccd1 _6368_/A1 sky130_fd_sc_hd__buf_4
Xinput151 mports_i[2] vssd1 vssd1 vccd1 vccd1 _4975_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6218__A1 _6628_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput162 mports_i[3] vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__buf_2
Xinput173 mports_i[4] vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__buf_2
XANTENNA__8758__A3 _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput184 mports_i[5] vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__buf_2
Xinput195 mports_i[6] vssd1 vssd1 vccd1 vccd1 _5131_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__7966__A1 _7971_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6769__A2 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7966__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7120__A _7120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7718__B2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7194__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5575__A _5575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5530_ _5510_/A _4930_/X _5511_/A _4933_/X _5529_/X vssd1 vssd1 vccd1 vccd1 _5530_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5461_ _5458_/X _5460_/X _6224_/S vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7200_ _7200_/A vssd1 vssd1 vccd1 vccd1 _7200_/X sky130_fd_sc_hd__buf_1
X_4412_ _8239_/A _6411_/A _4412_/C vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput603 _5546_/X vssd1 vssd1 vccd1 vccd1 sports_o[191] sky130_fd_sc_hd__buf_12
Xoutput614 _5802_/X vssd1 vssd1 vccd1 vccd1 sports_o[200] sky130_fd_sc_hd__buf_12
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8180_ _8180_/A vssd1 vssd1 vccd1 vccd1 _8194_/B sky130_fd_sc_hd__inv_2
X_5392_ _8140_/A _5389_/Y _6711_/S _5391_/Y vssd1 vssd1 vccd1 vccd1 _5392_/X sky130_fd_sc_hd__a211o_1
Xoutput625 _6092_/X vssd1 vssd1 vccd1 vccd1 sports_o[210] sky130_fd_sc_hd__buf_12
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput636 _6313_/X vssd1 vssd1 vccd1 vccd1 sports_o[220] sky130_fd_sc_hd__buf_12
Xoutput647 _7147_/X vssd1 vssd1 vccd1 vccd1 sports_o[25] sky130_fd_sc_hd__buf_12
XFILLER_0_111_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7131_ _5562_/X _7023_/X _7130_/X vssd1 vssd1 vccd1 vccd1 _7131_/X sky130_fd_sc_hd__o21a_1
X_4343_ hold41/A _4349_/A vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput658 _7196_/X vssd1 vssd1 vccd1 vccd1 sports_o[35] sky130_fd_sc_hd__buf_12
Xoutput669 _7240_/X vssd1 vssd1 vccd1 vccd1 sports_o[45] sky130_fd_sc_hd__buf_12
XFILLER_0_10_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7062_ _6526_/A _7059_/X _5161_/X _7246_/B _7061_/X vssd1 vssd1 vccd1 vccd1 _7062_/X
+ sky130_fd_sc_hd__a221o_1
X_6013_ _6891_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8825__S _8829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7957__A1 _8358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7957__B2 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4654__A hold44/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7964_ _7971_/A1 _4947_/B _7971_/B1 _5123_/A vssd1 vssd1 vccd1 vccd1 _7964_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5432__A2 _6635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6915_ _8150_/A _6102_/Y _6914_/X vssd1 vssd1 vccd1 vccd1 _6915_/Y sky130_fd_sc_hd__o21ai_2
X_7895_ _7760_/X _7886_/Y _7891_/X _7894_/Y vssd1 vssd1 vccd1 vccd1 _7895_/X sky130_fd_sc_hd__a22o_2
XANTENNA__7709__A1 _7707_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6846_ _7604_/B _6871_/B vssd1 vssd1 vccd1 vccd1 _6846_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__7185__A2 _7138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8382__A1 _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6393__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6777_ _6772_/Y _6924_/A _6773_/X _6776_/X vssd1 vssd1 vccd1 vccd1 _6777_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_80_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6932__A2 _6475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8516_ _8516_/A _8516_/B vssd1 vssd1 vccd1 vccd1 _8516_/Y sky130_fd_sc_hd__nand2_1
X_5728_ _6470_/B _5749_/A _5727_/Y vssd1 vssd1 vccd1 vccd1 _6780_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8447_ _8446_/X _8395_/X _8755_/B vssd1 vssd1 vccd1 vccd1 _8447_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5659_ _5659_/A _5827_/B vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5499__A2 _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6696__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8378_ _8378_/A vssd1 vssd1 vccd1 vccd1 _8435_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7329_ _7741_/S vssd1 vssd1 vccd1 vccd1 _7330_/A sky130_fd_sc_hd__inv_2
XANTENNA__6999__A2 _6994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5120__A1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5120__B2 _4939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7859__B _7859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5423__A2 _6875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7875__A _8174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8373__A1 _8372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6384__B1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7086__S _7097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8125__A1 _8132_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8125__B2 _5123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6136__B1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6687__A1 _5500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6687__B2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5842__B _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4739__A _6342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7636__B1 _8759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7100__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output520_A _7333_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7939__A1 _7944_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7939__B2 _7431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8600__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5414__A2 _5367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _6440_/A _6234_/B _6456_/A _5128_/A vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_98_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6700_ _5558_/X _7536_/B _7707_/B _5562_/X vssd1 vssd1 vccd1 vccd1 _6701_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7680_ _7680_/A _7680_/B vssd1 vssd1 vccd1 vccd1 _7680_/Y sky130_fd_sc_hd__nand2_1
X_4892_ _5274_/A vssd1 vssd1 vccd1 vccd1 _4893_/A sky130_fd_sc_hd__buf_8
XFILLER_0_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5178__A1 _5208_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6631_ _7451_/A _6475_/X _5394_/Y _6851_/B vssd1 vssd1 vccd1 vccd1 _6632_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5178__B2 _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6562_ _6562_/A _6958_/B vssd1 vssd1 vccd1 vccd1 _6562_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8116__A1 _8119_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8116__B2 _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8301_ _8755_/B vssd1 vssd1 vccd1 vccd1 _8513_/B sky130_fd_sc_hd__inv_2
X_5513_ _5510_/Y _4886_/A _5511_/Y _4891_/A _5512_/Y vssd1 vssd1 vccd1 vccd1 _7120_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6127__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8667__A2 _8577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6493_ _7345_/B _6429_/S _6491_/Y _6492_/X vssd1 vssd1 vccd1 vccd1 _6493_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6678__A1 _6432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8232_ _8235_/A1 _5299_/B _8235_/B1 _5171_/B _8231_/X vssd1 vssd1 vccd1 vccd1 _8232_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_124_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput400 _8822_/X vssd1 vssd1 vccd1 vccd1 mports_o[130] sky130_fd_sc_hd__buf_12
XFILLER_0_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5444_ _6079_/A _6653_/A vssd1 vssd1 vccd1 vccd1 _5444_/Y sky130_fd_sc_hd__nor2_1
Xoutput411 _8044_/X vssd1 vssd1 vccd1 vccd1 mports_o[18] sky130_fd_sc_hd__buf_12
XFILLER_0_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6848__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput422 _8197_/X vssd1 vssd1 vccd1 vccd1 mports_o[28] sky130_fd_sc_hd__buf_12
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput433 _8307_/X vssd1 vssd1 vccd1 vccd1 mports_o[38] sky130_fd_sc_hd__buf_12
XANTENNA__5350__A1 _5337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput444 _8399_/X vssd1 vssd1 vccd1 vccd1 mports_o[48] sky130_fd_sc_hd__buf_12
X_8163_ _8163_/A _8174_/B vssd1 vssd1 vccd1 vccd1 _8163_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5350__B2 _5191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput455 _8522_/X vssd1 vssd1 vccd1 vccd1 mports_o[58] sky130_fd_sc_hd__buf_12
X_5375_ _5159_/B _5362_/A _5374_/Y _5125_/X vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_100_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput466 _8592_/X vssd1 vssd1 vccd1 vccd1 mports_o[68] sky130_fd_sc_hd__buf_12
XFILLER_0_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7114_ _7114_/A vssd1 vssd1 vccd1 vccd1 _7114_/X sky130_fd_sc_hd__buf_1
Xoutput477 _8626_/X vssd1 vssd1 vccd1 vccd1 mports_o[78] sky130_fd_sc_hd__buf_12
Xoutput488 _8660_/X vssd1 vssd1 vccd1 vccd1 mports_o[88] sky130_fd_sc_hd__buf_12
X_4326_ _7847_/A _4326_/B vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__nand2_1
Xoutput499 _8694_/X vssd1 vssd1 vccd1 vccd1 mports_o[98] sky130_fd_sc_hd__buf_12
X_8094_ _8084_/Y _8174_/A _8085_/Y _7874_/A _8093_/Y vssd1 vssd1 vccd1 vccd1 _8094_/Y
+ sky130_fd_sc_hd__a221oi_1
XANTENNA__4368__B _4810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7045_ _5109_/B _7138_/A _7044_/X vssd1 vssd1 vccd1 vccd1 _7046_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__6583__B _6871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4384__A _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6602__A1 _7422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6602__B2 _6912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7947_ _7760_/X _8376_/A _7943_/X _7946_/X vssd1 vssd1 vccd1 vccd1 _7947_/X sky130_fd_sc_hd__a22o_4
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8355__A1 _7942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7878_ _7864_/Y _7874_/X _7865_/Y _7875_/X _7877_/Y vssd1 vssd1 vccd1 vccd1 _7878_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7158__A2 _7004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8355__B2 _8304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6366__B1 _6368_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6829_ _6827_/Y _6828_/Y _8150_/A vssd1 vssd1 vccd1 vccd1 _6829_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6905__A2 _6059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8107__B2 _7874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8658__A2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8949__RESET_B fanout732/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7866__B1 _7877_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6758__B _6758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4559__A _8181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7618__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4993__S _6356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8465__S hold26/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7589__B _7691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4294__A _8968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8594__A1 _8272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7397__A2 _7696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7149__A2 _7019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7857__B1 _7772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6668__B _6694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7609__B1 _7398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _8444_/A _5195_/A1 _8257_/C _5195_/B1 vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7085__A1 _5356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5091_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__buf_6
XANTENNA__5635__A2 _4935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6832__A1 _6827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8034__B1 _6411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8850_ _8893_/A _8850_/B vssd1 vssd1 vccd1 vccd1 _8856_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7388__A2 _7542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7801_ _7798_/X _7768_/X _7800_/X _7772_/X _7774_/X vssd1 vssd1 vccd1 vccd1 _7801_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5399__A1 _5031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8781_ _8423_/A _8711_/A _8486_/Y _8770_/B _8788_/S vssd1 vssd1 vccd1 vccd1 _8781_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6596__B1 _6968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5993_ _8160_/A _6231_/C _5993_/C vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__or3_1
XFILLER_0_91_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7732_ _6337_/X _7723_/B _7731_/X vssd1 vssd1 vccd1 vccd1 _7732_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8404__A _8404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ _6312_/A _7372_/B vssd1 vssd1 vccd1 vccd1 _5741_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_87_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6348__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7663_ _7661_/X _7723_/B _7662_/X vssd1 vssd1 vccd1 vccd1 _7663_/X sky130_fd_sc_hd__a21o_1
X_4875_ input80/X _8310_/B input17/X _4874_/X vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6614_ _6611_/A _6908_/B _6613_/X _6512_/X vssd1 vssd1 vccd1 vccd1 _6614_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7594_ _7542_/A _6811_/B _7326_/A vssd1 vssd1 vccd1 vccd1 _7594_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5571__A1 _5640_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6545_ _6543_/Y _6544_/Y _8188_/S vssd1 vssd1 vccd1 vccd1 _6545_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5571__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6476_ _6469_/X _6472_/X _6694_/B _7032_/A _6475_/X vssd1 vssd1 vccd1 vccd1 _6477_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6578__B _6578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8215_ _4312_/B _7316_/A _8222_/B1 _5359_/B _8214_/X vssd1 vssd1 vccd1 vccd1 _8215_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5427_ _5909_/B _7451_/A _5426_/Y _7629_/B vssd1 vssd1 vccd1 vccd1 _5427_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5874__A2 _4886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8146_ _8188_/S _8146_/B vssd1 vssd1 vccd1 vccd1 _8146_/Y sky130_fd_sc_hd__nor2_1
X_5358_ _5272_/A _4929_/A _5273_/A _4932_/A _5357_/X vssd1 vssd1 vccd1 vccd1 _5362_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7076__A1 _5248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8273__B1 _8364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4309_ _8954_/Q vssd1 vssd1 vccd1 vccd1 _4337_/A sky130_fd_sc_hd__buf_6
XANTENNA__8812__A2 _8803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8077_ _8080_/A1 _5780_/A _8080_/B1 _5079_/A vssd1 vssd1 vccd1 vccd1 _8077_/Y sky130_fd_sc_hd__o22ai_2
X_5289_ _5108_/A _5247_/X _5136_/A _5249_/Y _5288_/Y vssd1 vssd1 vccd1 vccd1 _5289_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5626__A2 _5192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6823__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7028_ _6461_/A _7019_/X _7012_/S vssd1 vssd1 vccd1 vccd1 _7028_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4834__B1 _4760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7379__A2 _5211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8979_ _8979_/CLK hold14/X input229/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8328__A1 _8333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6339__B1 _6264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4561__B hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5562__A1 _5575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5562__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5314__A1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5314__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7067__A1 _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6814__A1 _6801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6814__B2 _6828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7775__C1 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8319__A1 _7784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5250__B1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7790__A2 _7790_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4471__B _8189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4660_ _7778_/B _5359_/A _4560_/Y _5359_/B _4659_/Y vssd1 vssd1 vccd1 vccd1 _4661_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6679__A _6841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5553__A1 _6697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4591_ _4591_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _8845_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5553__B2 _5552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5583__A _6697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6330_ _6224_/S _7729_/B _6327_/X _6329_/Y vssd1 vssd1 vccd1 vccd1 _6330_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6261_ _6261_/A _6261_/B vssd1 vssd1 vccd1 vccd1 _6261_/X sky130_fd_sc_hd__or2_1
X_8000_ _7777_/X _7999_/Y _7792_/X vssd1 vssd1 vccd1 vccd1 _8000_/X sky130_fd_sc_hd__o21ba_1
X_5212_ _7013_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _6535_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6192_ _6192_/A vssd1 vssd1 vccd1 vccd1 _7686_/B sky130_fd_sc_hd__inv_2
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8255__B1 _8295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5143_ _6514_/B vssd1 vssd1 vccd1 vccd1 _7055_/A sky130_fd_sc_hd__inv_2
XANTENNA__4927__A _4927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5608__A2 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7303__A _7630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6805__A1 _5853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5074_ _5075_/B vssd1 vssd1 vccd1 vccd1 _6488_/A sky130_fd_sc_hd__inv_2
X_8902_ _4824_/B _8901_/Y _4800_/A vssd1 vssd1 vccd1 vccd1 _8903_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8833_ _8833_/A _8833_/B vssd1 vssd1 vccd1 vccd1 _8833_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6861__B _6925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7230__A1 _6185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8764_ _7956_/Y _8711_/A _8419_/X _8770_/B _8788_/S vssd1 vssd1 vccd1 vccd1 _8764_/X
+ sky130_fd_sc_hd__a221o_1
X_5976_ _5909_/B _7611_/A _5975_/X _5174_/A vssd1 vssd1 vccd1 vccd1 _5976_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7781__A2 _8295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7715_ _7714_/X _6261_/B _7715_/S vssd1 vssd1 vccd1 vccd1 _7715_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5792__A1 _5792_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4927_ _4927_/A vssd1 vssd1 vccd1 vccd1 _5111_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8695_ _8716_/A _4788_/C _8273_/X _8590_/A vssd1 vssd1 vccd1 vccd1 _8695_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5792__B2 _5193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7646_ _7701_/A _7646_/B vssd1 vssd1 vccd1 vccd1 _7646_/Y sky130_fd_sc_hd__nor2_1
X_4858_ _4858_/A vssd1 vssd1 vccd1 vccd1 _8933_/B sky130_fd_sc_hd__inv_2
XANTENNA__8191__C1 _7774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8730__A1 _7796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7533__A2 _8578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5544__A1 _5510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5544__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7577_ _7673_/A _7577_/B vssd1 vssd1 vccd1 vccd1 _7577_/Y sky130_fd_sc_hd__nor2_1
X_4789_ _4789_/A _4789_/B vssd1 vssd1 vccd1 vccd1 _4790_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6528_ _6528_/A vssd1 vssd1 vccd1 vccd1 _6882_/B sky130_fd_sc_hd__inv_2
XFILLER_0_31_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6459_ _6457_/Y _4986_/Y _6473_/A _7027_/A _6475_/A vssd1 vssd1 vccd1 vccd1 _6459_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5847__A2 _6788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5940__B _6231_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8246__B1 _8252_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8129_ _8132_/A1 _5780_/X _8132_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _8129_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__8797__A1 _8511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7213__A _7213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8797__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6272__A2 _8579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8549__A1 _4874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5480__B1 _5519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8549__B2 _8206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6771__B _7536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7221__A1 _6908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7883__A _7883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8964__RESET_B fanout733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8698__B _8698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8721__A1 _8309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8721__B2 _8711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6499__A _6499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5838__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8788__A1 _8055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6263__A2 _8523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7460__A1 _7673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6681__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6015__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7212__A1 _6095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5830_ _5830_/A vssd1 vssd1 vccd1 vccd1 _5830_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5223__B1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7763__A2 _5359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5761_ _6593_/A _5482_/B _5760_/Y vssd1 vssd1 vccd1 vccd1 _5762_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7500_ _5562_/X _7681_/A _7700_/B _7494_/Y vssd1 vssd1 vccd1 vccd1 _7500_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4712_ _4771_/A _4771_/B _4810_/B vssd1 vssd1 vccd1 vccd1 _4732_/B sky130_fd_sc_hd__nand3_1
X_8480_ _8480_/A _8480_/B vssd1 vssd1 vccd1 vccd1 _8480_/Y sky130_fd_sc_hd__nand2_1
X_5692_ _8140_/A _5689_/Y _7531_/A vssd1 vssd1 vccd1 vccd1 _5692_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7515__A2 _7297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7431_ _7767_/A _7431_/B _7432_/B vssd1 vssd1 vccd1 vccd1 _7431_/X sky130_fd_sc_hd__or3_1
X_4643_ hold31/A _4643_/B vssd1 vssd1 vccd1 vccd1 _8574_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_126_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7362_ _7575_/A vssd1 vssd1 vccd1 vccd1 _7363_/A sky130_fd_sc_hd__inv_2
X_4574_ hold21/X vssd1 vssd1 vccd1 vccd1 _4788_/C sky130_fd_sc_hd__inv_2
XFILLER_0_114_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6313_ _5125_/X _6298_/X _6307_/X _6311_/X _6312_/Y vssd1 vssd1 vccd1 vccd1 _6313_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7293_ _7754_/B _7138_/A _7292_/X vssd1 vssd1 vccd1 vccd1 _7294_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6244_ _6244_/A vssd1 vssd1 vccd1 vccd1 _7242_/A sky130_fd_sc_hd__inv_2
XANTENNA__6856__B _6958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8228__B1 _8234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5760__B _6593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6175_ input2/X _5191_/A _6158_/A _5102_/A _6174_/X vssd1 vssd1 vccd1 vccd1 _6212_/B
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6575__C _8185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7050__A_N _6497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5126_ _5159_/B _7345_/B _5124_/X _5125_/X vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4376__B _4591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5057_ _6304_/A _5050_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5057_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7203__A1 _6059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8816_ _8165_/Y _8738_/A _8169_/Y _8711_/A vssd1 vssd1 vccd1 vccd1 _8817_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5765__A1 _5518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8747_ _8746_/X _7886_/Y _8829_/S vssd1 vssd1 vccd1 vccd1 _8748_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4568__A2 _4478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5765__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5959_ _5958_/Y _5923_/Y _8842_/B vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8678_ _8148_/X _8583_/A _8803_/A _8581_/X _8621_/S vssd1 vssd1 vccd1 vccd1 _8678_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8703__A1 _8247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7506__A2 _5634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8703__B2 _8581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5935__B _6852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5517__A1 _6780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7629_ _7629_/A _7629_/B vssd1 vssd1 vccd1 vccd1 _7629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7208__A _7208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6112__A _6212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6190__B2 _5125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__8467__B1 _8304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5536__A1_N _6133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6478__C1 _6450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6493__A2 _6429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7690__A1 _7378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput300 sports_i[40] vssd1 vssd1 vccd1 vccd1 _7865_/A sky130_fd_sc_hd__buf_1
Xinput311 sports_i[50] vssd1 vssd1 vccd1 vccd1 _8003_/A sky130_fd_sc_hd__clkbuf_1
Xinput322 sports_i[60] vssd1 vssd1 vccd1 vccd1 _8142_/A sky130_fd_sc_hd__buf_2
Xinput333 sports_i[70] vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__buf_4
Xinput344 sports_i[80] vssd1 vssd1 vccd1 vccd1 _7958_/B1 sky130_fd_sc_hd__buf_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput355 sports_i[90] vssd1 vssd1 vccd1 vccd1 _8093_/B1 sky130_fd_sc_hd__buf_2
XANTENNA__6245__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7442__B2 _7754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6782__A _6852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7993__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5829__C _5829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5756__A1 _5787_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5756__B2 _4874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6006__B _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5845__B _5845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5508__B2 _4891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8170__A2 _8165_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 _6740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4290_ _8970_/Q vssd1 vssd1 vccd1 vccd1 _7510_/B sky130_fd_sc_hd__buf_12
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6676__B _7829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4477__A _6440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6236__A2 _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8630__B1 _7956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7980_ _7985_/A1 _5146_/A _7985_/B1 _7431_/B vssd1 vssd1 vccd1 vccd1 _7980_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__7984__A2 _7954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6931_ _6931_/A vssd1 vssd1 vccd1 vccd1 _6931_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5995__A1 _8140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4924__B _5108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7300__B _7575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6862_ _5923_/A _6510_/A _7610_/A _6512_/A vssd1 vssd1 vccd1 vccd1 _6862_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5101__A _5136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7736__A2 _7723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8601_ _8698_/B _8317_/X _8590_/X vssd1 vssd1 vccd1 vccd1 _8601_/X sky130_fd_sc_hd__o21a_1
X_5813_ _6079_/A _7171_/A vssd1 vssd1 vccd1 vccd1 _5813_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5747__B2 _5274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6793_ _5760_/A _5856_/A _6793_/S vssd1 vssd1 vccd1 vccd1 _7575_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8532_ _8165_/Y _8304_/X _8169_/Y _8299_/X _8496_/S vssd1 vssd1 vccd1 vccd1 _8532_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4940__A _4940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5744_ _5518_/A _5111_/A _5519_/A _4931_/A _5743_/X vssd1 vssd1 vccd1 vccd1 _5744_/X
+ sky130_fd_sc_hd__o221a_4
XANTENNA__8412__A _8412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8463_ _8323_/X _8453_/Y _8454_/Y _8462_/X vssd1 vssd1 vccd1 vccd1 _8463_/X sky130_fd_sc_hd__a31o_2
XFILLER_0_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4970__A2 _4868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5675_ _6875_/B _5573_/X _5674_/X vssd1 vssd1 vccd1 vccd1 _5675_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5247__S _6689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7414_ _5264_/Y _7680_/B _7412_/X _7640_/B _7413_/X vssd1 vssd1 vccd1 vccd1 _7414_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6172__A1 _6183_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4626_ _4626_/A vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__inv_2
X_8394_ _8394_/A _8550_/B vssd1 vssd1 vccd1 vccd1 _8394_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6172__B2 _5191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7345_ _7756_/A _7345_/B vssd1 vssd1 vccd1 vccd1 _7345_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4557_ _4557_/A _4557_/B vssd1 vssd1 vccd1 vccd1 _4590_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6867__A _6867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7276_ _7276_/A vssd1 vssd1 vccd1 vccd1 _7276_/X sky130_fd_sc_hd__buf_1
X_4488_ _8481_/S hold15/A vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__nand2_8
XANTENNA__5490__B _6202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6227_ _6227_/A vssd1 vssd1 vccd1 vccd1 _6227_/Y sky130_fd_sc_hd__inv_2
X_6158_ _6158_/A vssd1 vssd1 vccd1 vccd1 _6158_/Y sky130_fd_sc_hd__inv_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5109_ _6212_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__or2_1
X_6089_ _6089_/A1 _4934_/A input60/X _4938_/A vssd1 vssd1 vccd1 vccd1 _6089_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5710__S _8160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5986__A1 _6128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8306__B _8564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7188__B1 _5930_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6107__A _6107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7727__A2 _7349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6935__B1 _6450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5665__B _7532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8688__B1 _8206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4961__A2 _6234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6163__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6163__B2 _4893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5910__A1 _5962_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5910__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5681__A _5738_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4297__A _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput130 mports_i[216] vssd1 vssd1 vccd1 vccd1 _6229_/A2 sky130_fd_sc_hd__buf_2
Xinput141 mports_i[226] vssd1 vssd1 vccd1 vccd1 _6387_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput152 mports_i[30] vssd1 vssd1 vccd1 vccd1 _5788_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput163 mports_i[40] vssd1 vssd1 vccd1 vccd1 _6047_/A sky130_fd_sc_hd__clkbuf_4
Xinput174 mports_i[50] vssd1 vssd1 vccd1 vccd1 _6326_/A1 sky130_fd_sc_hd__buf_2
Xinput185 mports_i[60] vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5620__S _6547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput196 mports_i[70] vssd1 vssd1 vccd1 vccd1 _5273_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__7966__A2 _5146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7401__A _7590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5977__A1 _6031_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5977__B2 _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4744__B _7266_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6017__A _6017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7718__A2 _7753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8915__A1 _6470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4760__A _4760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8043__B1_N _7792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8679__B1 _8686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5460_ _5401_/A _4930_/X _5402_/A _4933_/A _5459_/X vssd1 vssd1 vccd1 vccd1 _5460_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4411_ _8185_/B _7847_/A vssd1 vssd1 vccd1 vccd1 _6411_/A sky130_fd_sc_hd__nor2_4
Xoutput604 _5570_/X vssd1 vssd1 vccd1 vccd1 sports_o[192] sky130_fd_sc_hd__buf_12
Xoutput615 _5822_/X vssd1 vssd1 vccd1 vccd1 sports_o[201] sky130_fd_sc_hd__buf_12
X_5391_ _5391_/A vssd1 vssd1 vccd1 vccd1 _5391_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5591__A _5591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput626 _6130_/X vssd1 vssd1 vccd1 vccd1 sports_o[211] sky130_fd_sc_hd__buf_12
XFILLER_0_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput637 _6330_/X vssd1 vssd1 vccd1 vccd1 sports_o[221] sky130_fd_sc_hd__buf_12
X_7130_ _6697_/B _7004_/X _5581_/Y _7088_/X _7089_/X vssd1 vssd1 vccd1 vccd1 _7130_/X
+ sky130_fd_sc_hd__a221o_2
Xoutput648 _7152_/X vssd1 vssd1 vccd1 vccd1 sports_o[26] sky130_fd_sc_hd__buf_12
XFILLER_0_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7103__A0 _7101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ hold26/A vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__inv_4
Xoutput659 _7200_/X vssd1 vssd1 vccd1 vccd1 sports_o[36] sky130_fd_sc_hd__buf_12
XFILLER_0_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7061_ _7089_/A vssd1 vssd1 vccd1 vccd1 _7061_/X sky130_fd_sc_hd__buf_8
X_6012_ _6020_/A _5080_/A _6021_/A _5089_/X _6011_/X vssd1 vssd1 vccd1 vccd1 _6891_/A
+ sky130_fd_sc_hd__o221a_2
.ends

