magic
tech sky130A
magscale 1 2
timestamp 1763066510
<< obsli1 >>
rect 1104 2159 158884 157777
<< obsm1 >>
rect 1104 76 159330 157808
<< metal2 >>
rect 12530 0 12586 800
rect 12990 0 13046 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17590 0 17646 800
rect 18050 0 18106 800
rect 18510 0 18566 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19890 0 19946 800
rect 20350 0 20406 800
rect 20810 0 20866 800
rect 21270 0 21326 800
rect 21730 0 21786 800
rect 22190 0 22246 800
rect 22650 0 22706 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24490 0 24546 800
rect 24950 0 25006 800
rect 25410 0 25466 800
rect 25870 0 25926 800
rect 26330 0 26386 800
rect 26790 0 26846 800
rect 27250 0 27306 800
rect 27710 0 27766 800
rect 28170 0 28226 800
rect 28630 0 28686 800
rect 29090 0 29146 800
rect 29550 0 29606 800
rect 30010 0 30066 800
rect 30470 0 30526 800
rect 30930 0 30986 800
rect 31390 0 31446 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32770 0 32826 800
rect 33230 0 33286 800
rect 33690 0 33746 800
rect 34150 0 34206 800
rect 34610 0 34666 800
rect 35070 0 35126 800
rect 35530 0 35586 800
rect 35990 0 36046 800
rect 36450 0 36506 800
rect 36910 0 36966 800
rect 37370 0 37426 800
rect 37830 0 37886 800
rect 38290 0 38346 800
rect 38750 0 38806 800
rect 39210 0 39266 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 41050 0 41106 800
rect 41510 0 41566 800
rect 41970 0 42026 800
rect 42430 0 42486 800
rect 42890 0 42946 800
rect 43350 0 43406 800
rect 43810 0 43866 800
rect 44270 0 44326 800
rect 44730 0 44786 800
rect 45190 0 45246 800
rect 45650 0 45706 800
rect 46110 0 46166 800
rect 46570 0 46626 800
rect 47030 0 47086 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48870 0 48926 800
rect 49330 0 49386 800
rect 49790 0 49846 800
rect 50250 0 50306 800
rect 50710 0 50766 800
rect 51170 0 51226 800
rect 51630 0 51686 800
rect 52090 0 52146 800
rect 52550 0 52606 800
rect 53010 0 53066 800
rect 53470 0 53526 800
rect 53930 0 53986 800
rect 54390 0 54446 800
rect 54850 0 54906 800
rect 55310 0 55366 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57150 0 57206 800
rect 57610 0 57666 800
rect 58070 0 58126 800
rect 58530 0 58586 800
rect 58990 0 59046 800
rect 59450 0 59506 800
rect 59910 0 59966 800
rect 60370 0 60426 800
rect 60830 0 60886 800
rect 61290 0 61346 800
rect 61750 0 61806 800
rect 62210 0 62266 800
rect 62670 0 62726 800
rect 63130 0 63186 800
rect 63590 0 63646 800
rect 64050 0 64106 800
rect 64510 0 64566 800
rect 64970 0 65026 800
rect 65430 0 65486 800
rect 65890 0 65946 800
rect 66350 0 66406 800
rect 66810 0 66866 800
rect 67270 0 67326 800
rect 67730 0 67786 800
rect 68190 0 68246 800
rect 68650 0 68706 800
rect 69110 0 69166 800
rect 69570 0 69626 800
rect 70030 0 70086 800
rect 70490 0 70546 800
rect 70950 0 71006 800
rect 71410 0 71466 800
rect 71870 0 71926 800
rect 72330 0 72386 800
rect 72790 0 72846 800
rect 73250 0 73306 800
rect 73710 0 73766 800
rect 74170 0 74226 800
rect 74630 0 74686 800
rect 75090 0 75146 800
rect 75550 0 75606 800
rect 76010 0 76066 800
rect 76470 0 76526 800
rect 76930 0 76986 800
rect 77390 0 77446 800
rect 77850 0 77906 800
rect 78310 0 78366 800
rect 78770 0 78826 800
rect 79230 0 79286 800
rect 79690 0 79746 800
rect 80150 0 80206 800
rect 80610 0 80666 800
rect 81070 0 81126 800
rect 81530 0 81586 800
rect 81990 0 82046 800
rect 82450 0 82506 800
rect 82910 0 82966 800
rect 83370 0 83426 800
rect 83830 0 83886 800
rect 84290 0 84346 800
rect 84750 0 84806 800
rect 85210 0 85266 800
rect 85670 0 85726 800
rect 86130 0 86186 800
rect 86590 0 86646 800
rect 87050 0 87106 800
rect 87510 0 87566 800
rect 87970 0 88026 800
rect 88430 0 88486 800
rect 88890 0 88946 800
rect 89350 0 89406 800
rect 89810 0 89866 800
rect 90270 0 90326 800
rect 90730 0 90786 800
rect 91190 0 91246 800
rect 91650 0 91706 800
rect 92110 0 92166 800
rect 92570 0 92626 800
rect 93030 0 93086 800
rect 93490 0 93546 800
rect 93950 0 94006 800
rect 94410 0 94466 800
rect 94870 0 94926 800
rect 95330 0 95386 800
rect 95790 0 95846 800
rect 96250 0 96306 800
rect 96710 0 96766 800
rect 97170 0 97226 800
rect 97630 0 97686 800
rect 98090 0 98146 800
rect 98550 0 98606 800
rect 99010 0 99066 800
rect 99470 0 99526 800
rect 99930 0 99986 800
rect 100390 0 100446 800
rect 100850 0 100906 800
rect 101310 0 101366 800
rect 101770 0 101826 800
rect 102230 0 102286 800
rect 102690 0 102746 800
rect 103150 0 103206 800
rect 103610 0 103666 800
rect 104070 0 104126 800
rect 104530 0 104586 800
rect 104990 0 105046 800
rect 105450 0 105506 800
rect 105910 0 105966 800
rect 106370 0 106426 800
rect 106830 0 106886 800
rect 107290 0 107346 800
rect 107750 0 107806 800
rect 108210 0 108266 800
rect 108670 0 108726 800
rect 109130 0 109186 800
rect 109590 0 109646 800
rect 110050 0 110106 800
rect 110510 0 110566 800
rect 110970 0 111026 800
rect 111430 0 111486 800
rect 111890 0 111946 800
rect 112350 0 112406 800
rect 112810 0 112866 800
rect 113270 0 113326 800
rect 113730 0 113786 800
rect 114190 0 114246 800
rect 114650 0 114706 800
rect 115110 0 115166 800
rect 115570 0 115626 800
rect 116030 0 116086 800
rect 116490 0 116546 800
rect 116950 0 117006 800
rect 117410 0 117466 800
rect 117870 0 117926 800
rect 118330 0 118386 800
rect 118790 0 118846 800
rect 119250 0 119306 800
rect 119710 0 119766 800
rect 120170 0 120226 800
rect 120630 0 120686 800
rect 121090 0 121146 800
rect 121550 0 121606 800
rect 122010 0 122066 800
rect 122470 0 122526 800
rect 122930 0 122986 800
rect 123390 0 123446 800
rect 123850 0 123906 800
rect 124310 0 124366 800
rect 124770 0 124826 800
rect 125230 0 125286 800
rect 125690 0 125746 800
rect 126150 0 126206 800
rect 126610 0 126666 800
rect 127070 0 127126 800
rect 127530 0 127586 800
rect 127990 0 128046 800
rect 128450 0 128506 800
rect 128910 0 128966 800
rect 129370 0 129426 800
rect 129830 0 129886 800
rect 130290 0 130346 800
rect 130750 0 130806 800
rect 131210 0 131266 800
rect 131670 0 131726 800
rect 132130 0 132186 800
rect 132590 0 132646 800
rect 133050 0 133106 800
rect 133510 0 133566 800
rect 133970 0 134026 800
rect 134430 0 134486 800
rect 134890 0 134946 800
rect 135350 0 135406 800
rect 135810 0 135866 800
rect 136270 0 136326 800
rect 136730 0 136786 800
rect 137190 0 137246 800
rect 137650 0 137706 800
rect 138110 0 138166 800
rect 138570 0 138626 800
rect 139030 0 139086 800
rect 139490 0 139546 800
rect 139950 0 140006 800
rect 140410 0 140466 800
rect 140870 0 140926 800
rect 141330 0 141386 800
rect 141790 0 141846 800
rect 142250 0 142306 800
rect 142710 0 142766 800
rect 143170 0 143226 800
rect 143630 0 143686 800
rect 144090 0 144146 800
rect 144550 0 144606 800
rect 145010 0 145066 800
rect 145470 0 145526 800
rect 145930 0 145986 800
rect 146390 0 146446 800
rect 146850 0 146906 800
rect 147310 0 147366 800
<< obsm2 >>
rect 3422 856 159324 158681
rect 3422 31 12474 856
rect 12642 31 12934 856
rect 13102 31 13394 856
rect 13562 31 13854 856
rect 14022 31 14314 856
rect 14482 31 14774 856
rect 14942 31 15234 856
rect 15402 31 15694 856
rect 15862 31 16154 856
rect 16322 31 16614 856
rect 16782 31 17074 856
rect 17242 31 17534 856
rect 17702 31 17994 856
rect 18162 31 18454 856
rect 18622 31 18914 856
rect 19082 31 19374 856
rect 19542 31 19834 856
rect 20002 31 20294 856
rect 20462 31 20754 856
rect 20922 31 21214 856
rect 21382 31 21674 856
rect 21842 31 22134 856
rect 22302 31 22594 856
rect 22762 31 23054 856
rect 23222 31 23514 856
rect 23682 31 23974 856
rect 24142 31 24434 856
rect 24602 31 24894 856
rect 25062 31 25354 856
rect 25522 31 25814 856
rect 25982 31 26274 856
rect 26442 31 26734 856
rect 26902 31 27194 856
rect 27362 31 27654 856
rect 27822 31 28114 856
rect 28282 31 28574 856
rect 28742 31 29034 856
rect 29202 31 29494 856
rect 29662 31 29954 856
rect 30122 31 30414 856
rect 30582 31 30874 856
rect 31042 31 31334 856
rect 31502 31 31794 856
rect 31962 31 32254 856
rect 32422 31 32714 856
rect 32882 31 33174 856
rect 33342 31 33634 856
rect 33802 31 34094 856
rect 34262 31 34554 856
rect 34722 31 35014 856
rect 35182 31 35474 856
rect 35642 31 35934 856
rect 36102 31 36394 856
rect 36562 31 36854 856
rect 37022 31 37314 856
rect 37482 31 37774 856
rect 37942 31 38234 856
rect 38402 31 38694 856
rect 38862 31 39154 856
rect 39322 31 39614 856
rect 39782 31 40074 856
rect 40242 31 40534 856
rect 40702 31 40994 856
rect 41162 31 41454 856
rect 41622 31 41914 856
rect 42082 31 42374 856
rect 42542 31 42834 856
rect 43002 31 43294 856
rect 43462 31 43754 856
rect 43922 31 44214 856
rect 44382 31 44674 856
rect 44842 31 45134 856
rect 45302 31 45594 856
rect 45762 31 46054 856
rect 46222 31 46514 856
rect 46682 31 46974 856
rect 47142 31 47434 856
rect 47602 31 47894 856
rect 48062 31 48354 856
rect 48522 31 48814 856
rect 48982 31 49274 856
rect 49442 31 49734 856
rect 49902 31 50194 856
rect 50362 31 50654 856
rect 50822 31 51114 856
rect 51282 31 51574 856
rect 51742 31 52034 856
rect 52202 31 52494 856
rect 52662 31 52954 856
rect 53122 31 53414 856
rect 53582 31 53874 856
rect 54042 31 54334 856
rect 54502 31 54794 856
rect 54962 31 55254 856
rect 55422 31 55714 856
rect 55882 31 56174 856
rect 56342 31 56634 856
rect 56802 31 57094 856
rect 57262 31 57554 856
rect 57722 31 58014 856
rect 58182 31 58474 856
rect 58642 31 58934 856
rect 59102 31 59394 856
rect 59562 31 59854 856
rect 60022 31 60314 856
rect 60482 31 60774 856
rect 60942 31 61234 856
rect 61402 31 61694 856
rect 61862 31 62154 856
rect 62322 31 62614 856
rect 62782 31 63074 856
rect 63242 31 63534 856
rect 63702 31 63994 856
rect 64162 31 64454 856
rect 64622 31 64914 856
rect 65082 31 65374 856
rect 65542 31 65834 856
rect 66002 31 66294 856
rect 66462 31 66754 856
rect 66922 31 67214 856
rect 67382 31 67674 856
rect 67842 31 68134 856
rect 68302 31 68594 856
rect 68762 31 69054 856
rect 69222 31 69514 856
rect 69682 31 69974 856
rect 70142 31 70434 856
rect 70602 31 70894 856
rect 71062 31 71354 856
rect 71522 31 71814 856
rect 71982 31 72274 856
rect 72442 31 72734 856
rect 72902 31 73194 856
rect 73362 31 73654 856
rect 73822 31 74114 856
rect 74282 31 74574 856
rect 74742 31 75034 856
rect 75202 31 75494 856
rect 75662 31 75954 856
rect 76122 31 76414 856
rect 76582 31 76874 856
rect 77042 31 77334 856
rect 77502 31 77794 856
rect 77962 31 78254 856
rect 78422 31 78714 856
rect 78882 31 79174 856
rect 79342 31 79634 856
rect 79802 31 80094 856
rect 80262 31 80554 856
rect 80722 31 81014 856
rect 81182 31 81474 856
rect 81642 31 81934 856
rect 82102 31 82394 856
rect 82562 31 82854 856
rect 83022 31 83314 856
rect 83482 31 83774 856
rect 83942 31 84234 856
rect 84402 31 84694 856
rect 84862 31 85154 856
rect 85322 31 85614 856
rect 85782 31 86074 856
rect 86242 31 86534 856
rect 86702 31 86994 856
rect 87162 31 87454 856
rect 87622 31 87914 856
rect 88082 31 88374 856
rect 88542 31 88834 856
rect 89002 31 89294 856
rect 89462 31 89754 856
rect 89922 31 90214 856
rect 90382 31 90674 856
rect 90842 31 91134 856
rect 91302 31 91594 856
rect 91762 31 92054 856
rect 92222 31 92514 856
rect 92682 31 92974 856
rect 93142 31 93434 856
rect 93602 31 93894 856
rect 94062 31 94354 856
rect 94522 31 94814 856
rect 94982 31 95274 856
rect 95442 31 95734 856
rect 95902 31 96194 856
rect 96362 31 96654 856
rect 96822 31 97114 856
rect 97282 31 97574 856
rect 97742 31 98034 856
rect 98202 31 98494 856
rect 98662 31 98954 856
rect 99122 31 99414 856
rect 99582 31 99874 856
rect 100042 31 100334 856
rect 100502 31 100794 856
rect 100962 31 101254 856
rect 101422 31 101714 856
rect 101882 31 102174 856
rect 102342 31 102634 856
rect 102802 31 103094 856
rect 103262 31 103554 856
rect 103722 31 104014 856
rect 104182 31 104474 856
rect 104642 31 104934 856
rect 105102 31 105394 856
rect 105562 31 105854 856
rect 106022 31 106314 856
rect 106482 31 106774 856
rect 106942 31 107234 856
rect 107402 31 107694 856
rect 107862 31 108154 856
rect 108322 31 108614 856
rect 108782 31 109074 856
rect 109242 31 109534 856
rect 109702 31 109994 856
rect 110162 31 110454 856
rect 110622 31 110914 856
rect 111082 31 111374 856
rect 111542 31 111834 856
rect 112002 31 112294 856
rect 112462 31 112754 856
rect 112922 31 113214 856
rect 113382 31 113674 856
rect 113842 31 114134 856
rect 114302 31 114594 856
rect 114762 31 115054 856
rect 115222 31 115514 856
rect 115682 31 115974 856
rect 116142 31 116434 856
rect 116602 31 116894 856
rect 117062 31 117354 856
rect 117522 31 117814 856
rect 117982 31 118274 856
rect 118442 31 118734 856
rect 118902 31 119194 856
rect 119362 31 119654 856
rect 119822 31 120114 856
rect 120282 31 120574 856
rect 120742 31 121034 856
rect 121202 31 121494 856
rect 121662 31 121954 856
rect 122122 31 122414 856
rect 122582 31 122874 856
rect 123042 31 123334 856
rect 123502 31 123794 856
rect 123962 31 124254 856
rect 124422 31 124714 856
rect 124882 31 125174 856
rect 125342 31 125634 856
rect 125802 31 126094 856
rect 126262 31 126554 856
rect 126722 31 127014 856
rect 127182 31 127474 856
rect 127642 31 127934 856
rect 128102 31 128394 856
rect 128562 31 128854 856
rect 129022 31 129314 856
rect 129482 31 129774 856
rect 129942 31 130234 856
rect 130402 31 130694 856
rect 130862 31 131154 856
rect 131322 31 131614 856
rect 131782 31 132074 856
rect 132242 31 132534 856
rect 132702 31 132994 856
rect 133162 31 133454 856
rect 133622 31 133914 856
rect 134082 31 134374 856
rect 134542 31 134834 856
rect 135002 31 135294 856
rect 135462 31 135754 856
rect 135922 31 136214 856
rect 136382 31 136674 856
rect 136842 31 137134 856
rect 137302 31 137594 856
rect 137762 31 138054 856
rect 138222 31 138514 856
rect 138682 31 138974 856
rect 139142 31 139434 856
rect 139602 31 139894 856
rect 140062 31 140354 856
rect 140522 31 140814 856
rect 140982 31 141274 856
rect 141442 31 141734 856
rect 141902 31 142194 856
rect 142362 31 142654 856
rect 142822 31 143114 856
rect 143282 31 143574 856
rect 143742 31 144034 856
rect 144202 31 144494 856
rect 144662 31 144954 856
rect 145122 31 145414 856
rect 145582 31 145874 856
rect 146042 31 146334 856
rect 146502 31 146794 856
rect 146962 31 147254 856
rect 147422 31 159324 856
<< metal3 >>
rect 159200 158584 160000 158704
rect 159200 157224 160000 157344
rect 0 155864 800 155984
rect 159200 155864 160000 155984
rect 159200 154504 160000 154624
rect 159200 153144 160000 153264
rect 159200 151784 160000 151904
rect 159200 150424 160000 150544
rect 159200 149064 160000 149184
rect 0 148248 800 148368
rect 159200 147704 160000 147824
rect 159200 146344 160000 146464
rect 159200 144984 160000 145104
rect 159200 143624 160000 143744
rect 159200 142264 160000 142384
rect 159200 140904 160000 141024
rect 0 140632 800 140752
rect 159200 139544 160000 139664
rect 159200 138184 160000 138304
rect 159200 136824 160000 136944
rect 159200 135464 160000 135584
rect 159200 134104 160000 134224
rect 0 133016 800 133136
rect 159200 132744 160000 132864
rect 159200 131384 160000 131504
rect 159200 130024 160000 130144
rect 159200 128664 160000 128784
rect 159200 127304 160000 127424
rect 159200 125944 160000 126064
rect 0 125400 800 125520
rect 159200 124584 160000 124704
rect 159200 123224 160000 123344
rect 159200 121864 160000 121984
rect 159200 120504 160000 120624
rect 159200 119144 160000 119264
rect 0 117784 800 117904
rect 159200 117784 160000 117904
rect 159200 116424 160000 116544
rect 159200 115064 160000 115184
rect 159200 113704 160000 113824
rect 159200 112344 160000 112464
rect 159200 110984 160000 111104
rect 0 110168 800 110288
rect 159200 109624 160000 109744
rect 159200 108264 160000 108384
rect 159200 106904 160000 107024
rect 159200 105544 160000 105664
rect 159200 104184 160000 104304
rect 159200 102824 160000 102944
rect 0 102552 800 102672
rect 159200 101464 160000 101584
rect 159200 100104 160000 100224
rect 159200 98744 160000 98864
rect 159200 97384 160000 97504
rect 159200 96024 160000 96144
rect 0 94936 800 95056
rect 159200 94664 160000 94784
rect 159200 93304 160000 93424
rect 159200 91944 160000 92064
rect 159200 90584 160000 90704
rect 159200 89224 160000 89344
rect 159200 87864 160000 87984
rect 0 87320 800 87440
rect 159200 86504 160000 86624
rect 159200 85144 160000 85264
rect 159200 83784 160000 83904
rect 159200 82424 160000 82544
rect 159200 81064 160000 81184
rect 0 79704 800 79824
rect 159200 79704 160000 79824
rect 159200 78344 160000 78464
rect 159200 76984 160000 77104
rect 159200 75624 160000 75744
rect 159200 74264 160000 74384
rect 159200 72904 160000 73024
rect 0 72088 800 72208
rect 159200 71544 160000 71664
rect 159200 70184 160000 70304
rect 159200 68824 160000 68944
rect 159200 67464 160000 67584
rect 159200 66104 160000 66224
rect 159200 64744 160000 64864
rect 0 64472 800 64592
rect 159200 63384 160000 63504
rect 159200 62024 160000 62144
rect 159200 60664 160000 60784
rect 159200 59304 160000 59424
rect 159200 57944 160000 58064
rect 0 56856 800 56976
rect 159200 56584 160000 56704
rect 159200 55224 160000 55344
rect 159200 53864 160000 53984
rect 159200 52504 160000 52624
rect 159200 51144 160000 51264
rect 159200 49784 160000 49904
rect 0 49240 800 49360
rect 159200 48424 160000 48544
rect 159200 47064 160000 47184
rect 159200 45704 160000 45824
rect 159200 44344 160000 44464
rect 159200 42984 160000 43104
rect 0 41624 800 41744
rect 159200 41624 160000 41744
rect 159200 40264 160000 40384
rect 159200 38904 160000 39024
rect 159200 37544 160000 37664
rect 159200 36184 160000 36304
rect 159200 34824 160000 34944
rect 0 34008 800 34128
rect 159200 33464 160000 33584
rect 159200 32104 160000 32224
rect 159200 30744 160000 30864
rect 159200 29384 160000 29504
rect 159200 28024 160000 28144
rect 159200 26664 160000 26784
rect 0 26392 800 26512
rect 159200 25304 160000 25424
rect 159200 23944 160000 24064
rect 159200 22584 160000 22704
rect 159200 21224 160000 21344
rect 159200 19864 160000 19984
rect 0 18776 800 18896
rect 159200 18504 160000 18624
rect 159200 17144 160000 17264
rect 159200 15784 160000 15904
rect 159200 14424 160000 14544
rect 159200 13064 160000 13184
rect 159200 11704 160000 11824
rect 0 11160 800 11280
rect 159200 10344 160000 10464
rect 159200 8984 160000 9104
rect 159200 7624 160000 7744
rect 159200 6264 160000 6384
rect 159200 4904 160000 5024
rect 0 3544 800 3664
rect 159200 3544 160000 3664
rect 159200 2184 160000 2304
rect 159200 824 160000 944
<< obsm3 >>
rect 800 158504 159120 158677
rect 800 157424 159200 158504
rect 800 157144 159120 157424
rect 800 156064 159200 157144
rect 880 155784 159120 156064
rect 800 154704 159200 155784
rect 800 154424 159120 154704
rect 800 153344 159200 154424
rect 800 153064 159120 153344
rect 800 151984 159200 153064
rect 800 151704 159120 151984
rect 800 150624 159200 151704
rect 800 150344 159120 150624
rect 800 149264 159200 150344
rect 800 148984 159120 149264
rect 800 148448 159200 148984
rect 880 148168 159200 148448
rect 800 147904 159200 148168
rect 800 147624 159120 147904
rect 800 146544 159200 147624
rect 800 146264 159120 146544
rect 800 145184 159200 146264
rect 800 144904 159120 145184
rect 800 143824 159200 144904
rect 800 143544 159120 143824
rect 800 142464 159200 143544
rect 800 142184 159120 142464
rect 800 141104 159200 142184
rect 800 140832 159120 141104
rect 880 140824 159120 140832
rect 880 140552 159200 140824
rect 800 139744 159200 140552
rect 800 139464 159120 139744
rect 800 138384 159200 139464
rect 800 138104 159120 138384
rect 800 137024 159200 138104
rect 800 136744 159120 137024
rect 800 135664 159200 136744
rect 800 135384 159120 135664
rect 800 134304 159200 135384
rect 800 134024 159120 134304
rect 800 133216 159200 134024
rect 880 132944 159200 133216
rect 880 132936 159120 132944
rect 800 132664 159120 132936
rect 800 131584 159200 132664
rect 800 131304 159120 131584
rect 800 130224 159200 131304
rect 800 129944 159120 130224
rect 800 128864 159200 129944
rect 800 128584 159120 128864
rect 800 127504 159200 128584
rect 800 127224 159120 127504
rect 800 126144 159200 127224
rect 800 125864 159120 126144
rect 800 125600 159200 125864
rect 880 125320 159200 125600
rect 800 124784 159200 125320
rect 800 124504 159120 124784
rect 800 123424 159200 124504
rect 800 123144 159120 123424
rect 800 122064 159200 123144
rect 800 121784 159120 122064
rect 800 120704 159200 121784
rect 800 120424 159120 120704
rect 800 119344 159200 120424
rect 800 119064 159120 119344
rect 800 117984 159200 119064
rect 880 117704 159120 117984
rect 800 116624 159200 117704
rect 800 116344 159120 116624
rect 800 115264 159200 116344
rect 800 114984 159120 115264
rect 800 113904 159200 114984
rect 800 113624 159120 113904
rect 800 112544 159200 113624
rect 800 112264 159120 112544
rect 800 111184 159200 112264
rect 800 110904 159120 111184
rect 800 110368 159200 110904
rect 880 110088 159200 110368
rect 800 109824 159200 110088
rect 800 109544 159120 109824
rect 800 108464 159200 109544
rect 800 108184 159120 108464
rect 800 107104 159200 108184
rect 800 106824 159120 107104
rect 800 105744 159200 106824
rect 800 105464 159120 105744
rect 800 104384 159200 105464
rect 800 104104 159120 104384
rect 800 103024 159200 104104
rect 800 102752 159120 103024
rect 880 102744 159120 102752
rect 880 102472 159200 102744
rect 800 101664 159200 102472
rect 800 101384 159120 101664
rect 800 100304 159200 101384
rect 800 100024 159120 100304
rect 800 98944 159200 100024
rect 800 98664 159120 98944
rect 800 97584 159200 98664
rect 800 97304 159120 97584
rect 800 96224 159200 97304
rect 800 95944 159120 96224
rect 800 95136 159200 95944
rect 880 94864 159200 95136
rect 880 94856 159120 94864
rect 800 94584 159120 94856
rect 800 93504 159200 94584
rect 800 93224 159120 93504
rect 800 92144 159200 93224
rect 800 91864 159120 92144
rect 800 90784 159200 91864
rect 800 90504 159120 90784
rect 800 89424 159200 90504
rect 800 89144 159120 89424
rect 800 88064 159200 89144
rect 800 87784 159120 88064
rect 800 87520 159200 87784
rect 880 87240 159200 87520
rect 800 86704 159200 87240
rect 800 86424 159120 86704
rect 800 85344 159200 86424
rect 800 85064 159120 85344
rect 800 83984 159200 85064
rect 800 83704 159120 83984
rect 800 82624 159200 83704
rect 800 82344 159120 82624
rect 800 81264 159200 82344
rect 800 80984 159120 81264
rect 800 79904 159200 80984
rect 880 79624 159120 79904
rect 800 78544 159200 79624
rect 800 78264 159120 78544
rect 800 77184 159200 78264
rect 800 76904 159120 77184
rect 800 75824 159200 76904
rect 800 75544 159120 75824
rect 800 74464 159200 75544
rect 800 74184 159120 74464
rect 800 73104 159200 74184
rect 800 72824 159120 73104
rect 800 72288 159200 72824
rect 880 72008 159200 72288
rect 800 71744 159200 72008
rect 800 71464 159120 71744
rect 800 70384 159200 71464
rect 800 70104 159120 70384
rect 800 69024 159200 70104
rect 800 68744 159120 69024
rect 800 67664 159200 68744
rect 800 67384 159120 67664
rect 800 66304 159200 67384
rect 800 66024 159120 66304
rect 800 64944 159200 66024
rect 800 64672 159120 64944
rect 880 64664 159120 64672
rect 880 64392 159200 64664
rect 800 63584 159200 64392
rect 800 63304 159120 63584
rect 800 62224 159200 63304
rect 800 61944 159120 62224
rect 800 60864 159200 61944
rect 800 60584 159120 60864
rect 800 59504 159200 60584
rect 800 59224 159120 59504
rect 800 58144 159200 59224
rect 800 57864 159120 58144
rect 800 57056 159200 57864
rect 880 56784 159200 57056
rect 880 56776 159120 56784
rect 800 56504 159120 56776
rect 800 55424 159200 56504
rect 800 55144 159120 55424
rect 800 54064 159200 55144
rect 800 53784 159120 54064
rect 800 52704 159200 53784
rect 800 52424 159120 52704
rect 800 51344 159200 52424
rect 800 51064 159120 51344
rect 800 49984 159200 51064
rect 800 49704 159120 49984
rect 800 49440 159200 49704
rect 880 49160 159200 49440
rect 800 48624 159200 49160
rect 800 48344 159120 48624
rect 800 47264 159200 48344
rect 800 46984 159120 47264
rect 800 45904 159200 46984
rect 800 45624 159120 45904
rect 800 44544 159200 45624
rect 800 44264 159120 44544
rect 800 43184 159200 44264
rect 800 42904 159120 43184
rect 800 41824 159200 42904
rect 880 41544 159120 41824
rect 800 40464 159200 41544
rect 800 40184 159120 40464
rect 800 39104 159200 40184
rect 800 38824 159120 39104
rect 800 37744 159200 38824
rect 800 37464 159120 37744
rect 800 36384 159200 37464
rect 800 36104 159120 36384
rect 800 35024 159200 36104
rect 800 34744 159120 35024
rect 800 34208 159200 34744
rect 880 33928 159200 34208
rect 800 33664 159200 33928
rect 800 33384 159120 33664
rect 800 32304 159200 33384
rect 800 32024 159120 32304
rect 800 30944 159200 32024
rect 800 30664 159120 30944
rect 800 29584 159200 30664
rect 800 29304 159120 29584
rect 800 28224 159200 29304
rect 800 27944 159120 28224
rect 800 26864 159200 27944
rect 800 26592 159120 26864
rect 880 26584 159120 26592
rect 880 26312 159200 26584
rect 800 25504 159200 26312
rect 800 25224 159120 25504
rect 800 24144 159200 25224
rect 800 23864 159120 24144
rect 800 22784 159200 23864
rect 800 22504 159120 22784
rect 800 21424 159200 22504
rect 800 21144 159120 21424
rect 800 20064 159200 21144
rect 800 19784 159120 20064
rect 800 18976 159200 19784
rect 880 18704 159200 18976
rect 880 18696 159120 18704
rect 800 18424 159120 18696
rect 800 17344 159200 18424
rect 800 17064 159120 17344
rect 800 15984 159200 17064
rect 800 15704 159120 15984
rect 800 14624 159200 15704
rect 800 14344 159120 14624
rect 800 13264 159200 14344
rect 800 12984 159120 13264
rect 800 11904 159200 12984
rect 800 11624 159120 11904
rect 800 11360 159200 11624
rect 880 11080 159200 11360
rect 800 10544 159200 11080
rect 800 10264 159120 10544
rect 800 9184 159200 10264
rect 800 8904 159120 9184
rect 800 7824 159200 8904
rect 800 7544 159120 7824
rect 800 6464 159200 7544
rect 800 6184 159120 6464
rect 800 5104 159200 6184
rect 800 4824 159120 5104
rect 800 3744 159200 4824
rect 880 3464 159120 3744
rect 800 2384 159200 3464
rect 800 2104 159120 2384
rect 800 1024 159200 2104
rect 800 744 159120 1024
rect 800 35 159200 744
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
rect 157808 2128 158128 157808
<< obsm4 >>
rect 35571 2048 50208 157045
rect 50688 2048 65568 157045
rect 66048 2048 80928 157045
rect 81408 2048 96288 157045
rect 96768 2048 111648 157045
rect 112128 2048 127008 157045
rect 127488 2048 142368 157045
rect 142848 2048 155973 157045
rect 35571 171 155973 2048
<< labels >>
rlabel metal2 s 14830 0 14886 800 6 busy_o
port 1 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 clk_i
port 2 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 discard_o
port 3 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 init_o
port 4 nsew signal output
rlabel metal3 s 159200 824 160000 944 6 mstream_i
port 5 nsew signal input
rlabel metal3 s 159200 2184 160000 2304 6 mstream_o[0]
port 6 nsew signal output
rlabel metal3 s 159200 138184 160000 138304 6 mstream_o[100]
port 7 nsew signal output
rlabel metal3 s 159200 139544 160000 139664 6 mstream_o[101]
port 8 nsew signal output
rlabel metal3 s 159200 140904 160000 141024 6 mstream_o[102]
port 9 nsew signal output
rlabel metal3 s 159200 142264 160000 142384 6 mstream_o[103]
port 10 nsew signal output
rlabel metal3 s 159200 143624 160000 143744 6 mstream_o[104]
port 11 nsew signal output
rlabel metal3 s 159200 144984 160000 145104 6 mstream_o[105]
port 12 nsew signal output
rlabel metal3 s 159200 146344 160000 146464 6 mstream_o[106]
port 13 nsew signal output
rlabel metal3 s 159200 147704 160000 147824 6 mstream_o[107]
port 14 nsew signal output
rlabel metal3 s 159200 149064 160000 149184 6 mstream_o[108]
port 15 nsew signal output
rlabel metal3 s 159200 150424 160000 150544 6 mstream_o[109]
port 16 nsew signal output
rlabel metal3 s 159200 15784 160000 15904 6 mstream_o[10]
port 17 nsew signal output
rlabel metal3 s 159200 151784 160000 151904 6 mstream_o[110]
port 18 nsew signal output
rlabel metal3 s 159200 153144 160000 153264 6 mstream_o[111]
port 19 nsew signal output
rlabel metal3 s 159200 154504 160000 154624 6 mstream_o[112]
port 20 nsew signal output
rlabel metal3 s 159200 155864 160000 155984 6 mstream_o[113]
port 21 nsew signal output
rlabel metal3 s 159200 157224 160000 157344 6 mstream_o[114]
port 22 nsew signal output
rlabel metal3 s 159200 158584 160000 158704 6 mstream_o[115]
port 23 nsew signal output
rlabel metal3 s 159200 17144 160000 17264 6 mstream_o[11]
port 24 nsew signal output
rlabel metal3 s 159200 18504 160000 18624 6 mstream_o[12]
port 25 nsew signal output
rlabel metal3 s 159200 19864 160000 19984 6 mstream_o[13]
port 26 nsew signal output
rlabel metal3 s 159200 21224 160000 21344 6 mstream_o[14]
port 27 nsew signal output
rlabel metal3 s 159200 22584 160000 22704 6 mstream_o[15]
port 28 nsew signal output
rlabel metal3 s 159200 23944 160000 24064 6 mstream_o[16]
port 29 nsew signal output
rlabel metal3 s 159200 25304 160000 25424 6 mstream_o[17]
port 30 nsew signal output
rlabel metal3 s 159200 26664 160000 26784 6 mstream_o[18]
port 31 nsew signal output
rlabel metal3 s 159200 28024 160000 28144 6 mstream_o[19]
port 32 nsew signal output
rlabel metal3 s 159200 3544 160000 3664 6 mstream_o[1]
port 33 nsew signal output
rlabel metal3 s 159200 29384 160000 29504 6 mstream_o[20]
port 34 nsew signal output
rlabel metal3 s 159200 30744 160000 30864 6 mstream_o[21]
port 35 nsew signal output
rlabel metal3 s 159200 32104 160000 32224 6 mstream_o[22]
port 36 nsew signal output
rlabel metal3 s 159200 33464 160000 33584 6 mstream_o[23]
port 37 nsew signal output
rlabel metal3 s 159200 34824 160000 34944 6 mstream_o[24]
port 38 nsew signal output
rlabel metal3 s 159200 36184 160000 36304 6 mstream_o[25]
port 39 nsew signal output
rlabel metal3 s 159200 37544 160000 37664 6 mstream_o[26]
port 40 nsew signal output
rlabel metal3 s 159200 38904 160000 39024 6 mstream_o[27]
port 41 nsew signal output
rlabel metal3 s 159200 40264 160000 40384 6 mstream_o[28]
port 42 nsew signal output
rlabel metal3 s 159200 41624 160000 41744 6 mstream_o[29]
port 43 nsew signal output
rlabel metal3 s 159200 4904 160000 5024 6 mstream_o[2]
port 44 nsew signal output
rlabel metal3 s 159200 42984 160000 43104 6 mstream_o[30]
port 45 nsew signal output
rlabel metal3 s 159200 44344 160000 44464 6 mstream_o[31]
port 46 nsew signal output
rlabel metal3 s 159200 45704 160000 45824 6 mstream_o[32]
port 47 nsew signal output
rlabel metal3 s 159200 47064 160000 47184 6 mstream_o[33]
port 48 nsew signal output
rlabel metal3 s 159200 48424 160000 48544 6 mstream_o[34]
port 49 nsew signal output
rlabel metal3 s 159200 49784 160000 49904 6 mstream_o[35]
port 50 nsew signal output
rlabel metal3 s 159200 51144 160000 51264 6 mstream_o[36]
port 51 nsew signal output
rlabel metal3 s 159200 52504 160000 52624 6 mstream_o[37]
port 52 nsew signal output
rlabel metal3 s 159200 53864 160000 53984 6 mstream_o[38]
port 53 nsew signal output
rlabel metal3 s 159200 55224 160000 55344 6 mstream_o[39]
port 54 nsew signal output
rlabel metal3 s 159200 6264 160000 6384 6 mstream_o[3]
port 55 nsew signal output
rlabel metal3 s 159200 56584 160000 56704 6 mstream_o[40]
port 56 nsew signal output
rlabel metal3 s 159200 57944 160000 58064 6 mstream_o[41]
port 57 nsew signal output
rlabel metal3 s 159200 59304 160000 59424 6 mstream_o[42]
port 58 nsew signal output
rlabel metal3 s 159200 60664 160000 60784 6 mstream_o[43]
port 59 nsew signal output
rlabel metal3 s 159200 62024 160000 62144 6 mstream_o[44]
port 60 nsew signal output
rlabel metal3 s 159200 63384 160000 63504 6 mstream_o[45]
port 61 nsew signal output
rlabel metal3 s 159200 64744 160000 64864 6 mstream_o[46]
port 62 nsew signal output
rlabel metal3 s 159200 66104 160000 66224 6 mstream_o[47]
port 63 nsew signal output
rlabel metal3 s 159200 67464 160000 67584 6 mstream_o[48]
port 64 nsew signal output
rlabel metal3 s 159200 68824 160000 68944 6 mstream_o[49]
port 65 nsew signal output
rlabel metal3 s 159200 7624 160000 7744 6 mstream_o[4]
port 66 nsew signal output
rlabel metal3 s 159200 70184 160000 70304 6 mstream_o[50]
port 67 nsew signal output
rlabel metal3 s 159200 71544 160000 71664 6 mstream_o[51]
port 68 nsew signal output
rlabel metal3 s 159200 72904 160000 73024 6 mstream_o[52]
port 69 nsew signal output
rlabel metal3 s 159200 74264 160000 74384 6 mstream_o[53]
port 70 nsew signal output
rlabel metal3 s 159200 75624 160000 75744 6 mstream_o[54]
port 71 nsew signal output
rlabel metal3 s 159200 76984 160000 77104 6 mstream_o[55]
port 72 nsew signal output
rlabel metal3 s 159200 78344 160000 78464 6 mstream_o[56]
port 73 nsew signal output
rlabel metal3 s 159200 79704 160000 79824 6 mstream_o[57]
port 74 nsew signal output
rlabel metal3 s 159200 81064 160000 81184 6 mstream_o[58]
port 75 nsew signal output
rlabel metal3 s 159200 82424 160000 82544 6 mstream_o[59]
port 76 nsew signal output
rlabel metal3 s 159200 8984 160000 9104 6 mstream_o[5]
port 77 nsew signal output
rlabel metal3 s 159200 83784 160000 83904 6 mstream_o[60]
port 78 nsew signal output
rlabel metal3 s 159200 85144 160000 85264 6 mstream_o[61]
port 79 nsew signal output
rlabel metal3 s 159200 86504 160000 86624 6 mstream_o[62]
port 80 nsew signal output
rlabel metal3 s 159200 87864 160000 87984 6 mstream_o[63]
port 81 nsew signal output
rlabel metal3 s 159200 89224 160000 89344 6 mstream_o[64]
port 82 nsew signal output
rlabel metal3 s 159200 90584 160000 90704 6 mstream_o[65]
port 83 nsew signal output
rlabel metal3 s 159200 91944 160000 92064 6 mstream_o[66]
port 84 nsew signal output
rlabel metal3 s 159200 93304 160000 93424 6 mstream_o[67]
port 85 nsew signal output
rlabel metal3 s 159200 94664 160000 94784 6 mstream_o[68]
port 86 nsew signal output
rlabel metal3 s 159200 96024 160000 96144 6 mstream_o[69]
port 87 nsew signal output
rlabel metal3 s 159200 10344 160000 10464 6 mstream_o[6]
port 88 nsew signal output
rlabel metal3 s 159200 97384 160000 97504 6 mstream_o[70]
port 89 nsew signal output
rlabel metal3 s 159200 98744 160000 98864 6 mstream_o[71]
port 90 nsew signal output
rlabel metal3 s 159200 100104 160000 100224 6 mstream_o[72]
port 91 nsew signal output
rlabel metal3 s 159200 101464 160000 101584 6 mstream_o[73]
port 92 nsew signal output
rlabel metal3 s 159200 102824 160000 102944 6 mstream_o[74]
port 93 nsew signal output
rlabel metal3 s 159200 104184 160000 104304 6 mstream_o[75]
port 94 nsew signal output
rlabel metal3 s 159200 105544 160000 105664 6 mstream_o[76]
port 95 nsew signal output
rlabel metal3 s 159200 106904 160000 107024 6 mstream_o[77]
port 96 nsew signal output
rlabel metal3 s 159200 108264 160000 108384 6 mstream_o[78]
port 97 nsew signal output
rlabel metal3 s 159200 109624 160000 109744 6 mstream_o[79]
port 98 nsew signal output
rlabel metal3 s 159200 11704 160000 11824 6 mstream_o[7]
port 99 nsew signal output
rlabel metal3 s 159200 110984 160000 111104 6 mstream_o[80]
port 100 nsew signal output
rlabel metal3 s 159200 112344 160000 112464 6 mstream_o[81]
port 101 nsew signal output
rlabel metal3 s 159200 113704 160000 113824 6 mstream_o[82]
port 102 nsew signal output
rlabel metal3 s 159200 115064 160000 115184 6 mstream_o[83]
port 103 nsew signal output
rlabel metal3 s 159200 116424 160000 116544 6 mstream_o[84]
port 104 nsew signal output
rlabel metal3 s 159200 117784 160000 117904 6 mstream_o[85]
port 105 nsew signal output
rlabel metal3 s 159200 119144 160000 119264 6 mstream_o[86]
port 106 nsew signal output
rlabel metal3 s 159200 120504 160000 120624 6 mstream_o[87]
port 107 nsew signal output
rlabel metal3 s 159200 121864 160000 121984 6 mstream_o[88]
port 108 nsew signal output
rlabel metal3 s 159200 123224 160000 123344 6 mstream_o[89]
port 109 nsew signal output
rlabel metal3 s 159200 13064 160000 13184 6 mstream_o[8]
port 110 nsew signal output
rlabel metal3 s 159200 124584 160000 124704 6 mstream_o[90]
port 111 nsew signal output
rlabel metal3 s 159200 125944 160000 126064 6 mstream_o[91]
port 112 nsew signal output
rlabel metal3 s 159200 127304 160000 127424 6 mstream_o[92]
port 113 nsew signal output
rlabel metal3 s 159200 128664 160000 128784 6 mstream_o[93]
port 114 nsew signal output
rlabel metal3 s 159200 130024 160000 130144 6 mstream_o[94]
port 115 nsew signal output
rlabel metal3 s 159200 131384 160000 131504 6 mstream_o[95]
port 116 nsew signal output
rlabel metal3 s 159200 132744 160000 132864 6 mstream_o[96]
port 117 nsew signal output
rlabel metal3 s 159200 134104 160000 134224 6 mstream_o[97]
port 118 nsew signal output
rlabel metal3 s 159200 135464 160000 135584 6 mstream_o[98]
port 119 nsew signal output
rlabel metal3 s 159200 136824 160000 136944 6 mstream_o[99]
port 120 nsew signal output
rlabel metal3 s 159200 14424 160000 14544 6 mstream_o[9]
port 121 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 nrst_i
port 122 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 run_i
port 123 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 sstream_i[0]
port 124 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 sstream_i[10]
port 125 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 sstream_i[11]
port 126 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 sstream_i[12]
port 127 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 sstream_i[13]
port 128 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 sstream_i[14]
port 129 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 sstream_i[15]
port 130 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 sstream_i[16]
port 131 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 sstream_i[17]
port 132 nsew signal input
rlabel metal3 s 0 140632 800 140752 6 sstream_i[18]
port 133 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 sstream_i[19]
port 134 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 sstream_i[1]
port 135 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 sstream_i[2]
port 136 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 sstream_i[3]
port 137 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 sstream_i[4]
port 138 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 sstream_i[5]
port 139 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 sstream_i[6]
port 140 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 sstream_i[7]
port 141 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 sstream_i[8]
port 142 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 sstream_i[9]
port 143 nsew signal input
rlabel metal3 s 0 155864 800 155984 6 sstream_o
port 144 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 v0x[0]
port 145 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 v0x[10]
port 146 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 v0x[11]
port 147 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 v0x[12]
port 148 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 v0x[13]
port 149 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 v0x[14]
port 150 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 v0x[15]
port 151 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 v0x[16]
port 152 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 v0x[17]
port 153 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 v0x[18]
port 154 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 v0x[19]
port 155 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 v0x[1]
port 156 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 v0x[20]
port 157 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 v0x[21]
port 158 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 v0x[22]
port 159 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 v0x[23]
port 160 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 v0x[24]
port 161 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 v0x[25]
port 162 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 v0x[26]
port 163 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 v0x[27]
port 164 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 v0x[28]
port 165 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 v0x[29]
port 166 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 v0x[2]
port 167 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 v0x[30]
port 168 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 v0x[31]
port 169 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 v0x[3]
port 170 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 v0x[4]
port 171 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 v0x[5]
port 172 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 v0x[6]
port 173 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 v0x[7]
port 174 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 v0x[8]
port 175 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 v0x[9]
port 176 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 v0y[0]
port 177 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 v0y[10]
port 178 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 v0y[11]
port 179 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 v0y[12]
port 180 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 v0y[13]
port 181 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 v0y[14]
port 182 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 v0y[15]
port 183 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 v0y[16]
port 184 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 v0y[17]
port 185 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 v0y[18]
port 186 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 v0y[19]
port 187 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 v0y[1]
port 188 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 v0y[20]
port 189 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 v0y[21]
port 190 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 v0y[22]
port 191 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 v0y[23]
port 192 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 v0y[24]
port 193 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 v0y[25]
port 194 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 v0y[26]
port 195 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 v0y[27]
port 196 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 v0y[28]
port 197 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 v0y[29]
port 198 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 v0y[2]
port 199 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 v0y[30]
port 200 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 v0y[31]
port 201 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 v0y[3]
port 202 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 v0y[4]
port 203 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 v0y[5]
port 204 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 v0y[6]
port 205 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 v0y[7]
port 206 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 v0y[8]
port 207 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 v0y[9]
port 208 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 v0z[0]
port 209 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 v0z[10]
port 210 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 v0z[11]
port 211 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 v0z[12]
port 212 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 v0z[13]
port 213 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 v0z[14]
port 214 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 v0z[15]
port 215 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 v0z[16]
port 216 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 v0z[17]
port 217 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 v0z[18]
port 218 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 v0z[19]
port 219 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 v0z[1]
port 220 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 v0z[20]
port 221 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 v0z[21]
port 222 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 v0z[22]
port 223 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 v0z[23]
port 224 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 v0z[24]
port 225 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 v0z[25]
port 226 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 v0z[26]
port 227 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 v0z[27]
port 228 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 v0z[28]
port 229 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 v0z[29]
port 230 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 v0z[2]
port 231 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 v0z[30]
port 232 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 v0z[31]
port 233 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 v0z[3]
port 234 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 v0z[4]
port 235 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 v0z[5]
port 236 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 v0z[6]
port 237 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 v0z[7]
port 238 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 v0z[8]
port 239 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 v0z[9]
port 240 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 v1x[0]
port 241 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 v1x[10]
port 242 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 v1x[11]
port 243 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 v1x[12]
port 244 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 v1x[13]
port 245 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 v1x[14]
port 246 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 v1x[15]
port 247 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 v1x[16]
port 248 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 v1x[17]
port 249 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 v1x[18]
port 250 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 v1x[19]
port 251 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 v1x[1]
port 252 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 v1x[20]
port 253 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 v1x[21]
port 254 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 v1x[22]
port 255 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 v1x[23]
port 256 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 v1x[24]
port 257 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 v1x[25]
port 258 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 v1x[26]
port 259 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 v1x[27]
port 260 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 v1x[28]
port 261 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 v1x[29]
port 262 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 v1x[2]
port 263 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 v1x[30]
port 264 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 v1x[31]
port 265 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 v1x[3]
port 266 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 v1x[4]
port 267 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 v1x[5]
port 268 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 v1x[6]
port 269 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 v1x[7]
port 270 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 v1x[8]
port 271 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 v1x[9]
port 272 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 v1y[0]
port 273 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 v1y[10]
port 274 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 v1y[11]
port 275 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 v1y[12]
port 276 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 v1y[13]
port 277 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 v1y[14]
port 278 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 v1y[15]
port 279 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 v1y[16]
port 280 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 v1y[17]
port 281 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 v1y[18]
port 282 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 v1y[19]
port 283 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 v1y[1]
port 284 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 v1y[20]
port 285 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 v1y[21]
port 286 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 v1y[22]
port 287 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 v1y[23]
port 288 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 v1y[24]
port 289 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 v1y[25]
port 290 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 v1y[26]
port 291 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 v1y[27]
port 292 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 v1y[28]
port 293 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 v1y[29]
port 294 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 v1y[2]
port 295 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 v1y[30]
port 296 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 v1y[31]
port 297 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 v1y[3]
port 298 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 v1y[4]
port 299 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 v1y[5]
port 300 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 v1y[6]
port 301 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 v1y[7]
port 302 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 v1y[8]
port 303 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 v1y[9]
port 304 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 v1z[0]
port 305 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 v1z[10]
port 306 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 v1z[11]
port 307 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 v1z[12]
port 308 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 v1z[13]
port 309 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 v1z[14]
port 310 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 v1z[15]
port 311 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 v1z[16]
port 312 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 v1z[17]
port 313 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 v1z[18]
port 314 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 v1z[19]
port 315 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 v1z[1]
port 316 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 v1z[20]
port 317 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 v1z[21]
port 318 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 v1z[22]
port 319 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 v1z[23]
port 320 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 v1z[24]
port 321 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 v1z[25]
port 322 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 v1z[26]
port 323 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 v1z[27]
port 324 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 v1z[28]
port 325 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 v1z[29]
port 326 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 v1z[2]
port 327 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 v1z[30]
port 328 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 v1z[31]
port 329 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 v1z[3]
port 330 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 v1z[4]
port 331 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 v1z[5]
port 332 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 v1z[6]
port 333 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 v1z[7]
port 334 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 v1z[8]
port 335 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 v1z[9]
port 336 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 v2x[0]
port 337 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 v2x[10]
port 338 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 v2x[11]
port 339 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 v2x[12]
port 340 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 v2x[13]
port 341 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 v2x[14]
port 342 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 v2x[15]
port 343 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 v2x[16]
port 344 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 v2x[17]
port 345 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 v2x[18]
port 346 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 v2x[19]
port 347 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 v2x[1]
port 348 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 v2x[20]
port 349 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 v2x[21]
port 350 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 v2x[22]
port 351 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 v2x[23]
port 352 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 v2x[24]
port 353 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 v2x[25]
port 354 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 v2x[26]
port 355 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 v2x[27]
port 356 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 v2x[28]
port 357 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 v2x[29]
port 358 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 v2x[2]
port 359 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 v2x[30]
port 360 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 v2x[31]
port 361 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 v2x[3]
port 362 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 v2x[4]
port 363 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 v2x[5]
port 364 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 v2x[6]
port 365 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 v2x[7]
port 366 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 v2x[8]
port 367 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 v2x[9]
port 368 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 v2y[0]
port 369 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 v2y[10]
port 370 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 v2y[11]
port 371 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 v2y[12]
port 372 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 v2y[13]
port 373 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 v2y[14]
port 374 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 v2y[15]
port 375 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 v2y[16]
port 376 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 v2y[17]
port 377 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 v2y[18]
port 378 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 v2y[19]
port 379 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 v2y[1]
port 380 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 v2y[20]
port 381 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 v2y[21]
port 382 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 v2y[22]
port 383 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 v2y[23]
port 384 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 v2y[24]
port 385 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 v2y[25]
port 386 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 v2y[26]
port 387 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 v2y[27]
port 388 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 v2y[28]
port 389 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 v2y[29]
port 390 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 v2y[2]
port 391 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 v2y[30]
port 392 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 v2y[31]
port 393 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 v2y[3]
port 394 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 v2y[4]
port 395 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 v2y[5]
port 396 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 v2y[6]
port 397 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 v2y[7]
port 398 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 v2y[8]
port 399 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 v2y[9]
port 400 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 v2z[0]
port 401 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 v2z[10]
port 402 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 v2z[11]
port 403 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 v2z[12]
port 404 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 v2z[13]
port 405 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 v2z[14]
port 406 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 v2z[15]
port 407 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 v2z[16]
port 408 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 v2z[17]
port 409 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 v2z[18]
port 410 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 v2z[19]
port 411 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 v2z[1]
port 412 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 v2z[20]
port 413 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 v2z[21]
port 414 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 v2z[22]
port 415 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 v2z[23]
port 416 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 v2z[24]
port 417 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 v2z[25]
port 418 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 v2z[26]
port 419 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 v2z[27]
port 420 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 v2z[28]
port 421 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 v2z[29]
port 422 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 v2z[2]
port 423 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 v2z[30]
port 424 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 v2z[31]
port 425 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 v2z[3]
port 426 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 v2z[4]
port 427 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 v2z[5]
port 428 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 v2z[6]
port 429 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 v2z[7]
port 430 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 v2z[8]
port 431 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 v2z[9]
port 432 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 434 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 160000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 50198744
string GDS_FILE /home/sforde22/Caravel/sdmay26-24/openlane/bary_pipe/runs/25_11_13_14_18/results/signoff/bary_pipe_m.magic.gds
string GDS_START 1752488
<< end >>

