magic
tech sky130A
magscale 1 2
timestamp 1761083769
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 934 1844 119586 117632
<< metal2 >>
rect 29918 119200 29974 120000
rect 89902 119200 89958 120000
rect 6090 0 6146 800
rect 18050 0 18106 800
rect 30010 0 30066 800
rect 41970 0 42026 800
rect 53930 0 53986 800
rect 65890 0 65946 800
rect 77850 0 77906 800
rect 89810 0 89866 800
rect 101770 0 101826 800
rect 113730 0 113786 800
<< obsm2 >>
rect 938 119144 29862 119200
rect 30030 119144 89846 119200
rect 90014 119144 119580 119200
rect 938 856 119580 119144
rect 938 734 6034 856
rect 6202 734 17994 856
rect 18162 734 29954 856
rect 30122 734 41914 856
rect 42082 734 53874 856
rect 54042 734 65834 856
rect 66002 734 77794 856
rect 77962 734 89754 856
rect 89922 734 101714 856
rect 101882 734 113674 856
rect 113842 734 119580 856
<< metal3 >>
rect 119200 118328 120000 118448
rect 119200 115608 120000 115728
rect 0 115336 800 115456
rect 0 113704 800 113824
rect 119200 112888 120000 113008
rect 0 112072 800 112192
rect 0 110440 800 110560
rect 119200 110168 120000 110288
rect 0 108808 800 108928
rect 119200 107448 120000 107568
rect 0 107176 800 107296
rect 0 105544 800 105664
rect 119200 104728 120000 104848
rect 0 103912 800 104032
rect 0 102280 800 102400
rect 119200 102008 120000 102128
rect 0 100648 800 100768
rect 119200 99288 120000 99408
rect 0 99016 800 99136
rect 0 97384 800 97504
rect 119200 96568 120000 96688
rect 0 95752 800 95872
rect 0 94120 800 94240
rect 119200 93848 120000 93968
rect 0 92488 800 92608
rect 119200 91128 120000 91248
rect 0 90856 800 90976
rect 0 89224 800 89344
rect 119200 88408 120000 88528
rect 0 87592 800 87712
rect 0 85960 800 86080
rect 119200 85688 120000 85808
rect 0 84328 800 84448
rect 119200 82968 120000 83088
rect 0 82696 800 82816
rect 0 81064 800 81184
rect 119200 80248 120000 80368
rect 0 79432 800 79552
rect 0 77800 800 77920
rect 119200 77528 120000 77648
rect 0 76168 800 76288
rect 119200 74808 120000 74928
rect 0 74536 800 74656
rect 0 72904 800 73024
rect 119200 72088 120000 72208
rect 0 71272 800 71392
rect 0 69640 800 69760
rect 119200 69368 120000 69488
rect 0 68008 800 68128
rect 119200 66648 120000 66768
rect 0 66376 800 66496
rect 0 64744 800 64864
rect 119200 63928 120000 64048
rect 0 63112 800 63232
rect 0 61480 800 61600
rect 119200 61208 120000 61328
rect 0 59848 800 59968
rect 119200 58488 120000 58608
rect 0 58216 800 58336
rect 0 56584 800 56704
rect 119200 55768 120000 55888
rect 0 54952 800 55072
rect 0 53320 800 53440
rect 119200 53048 120000 53168
rect 0 51688 800 51808
rect 119200 50328 120000 50448
rect 0 50056 800 50176
rect 0 48424 800 48544
rect 119200 47608 120000 47728
rect 0 46792 800 46912
rect 0 45160 800 45280
rect 119200 44888 120000 45008
rect 0 43528 800 43648
rect 119200 42168 120000 42288
rect 0 41896 800 42016
rect 0 40264 800 40384
rect 119200 39448 120000 39568
rect 0 38632 800 38752
rect 0 37000 800 37120
rect 119200 36728 120000 36848
rect 0 35368 800 35488
rect 119200 34008 120000 34128
rect 0 33736 800 33856
rect 0 32104 800 32224
rect 119200 31288 120000 31408
rect 0 30472 800 30592
rect 0 28840 800 28960
rect 119200 28568 120000 28688
rect 0 27208 800 27328
rect 119200 25848 120000 25968
rect 0 25576 800 25696
rect 0 23944 800 24064
rect 119200 23128 120000 23248
rect 0 22312 800 22432
rect 0 20680 800 20800
rect 119200 20408 120000 20528
rect 0 19048 800 19168
rect 119200 17688 120000 17808
rect 0 17416 800 17536
rect 0 15784 800 15904
rect 119200 14968 120000 15088
rect 0 14152 800 14272
rect 0 12520 800 12640
rect 119200 12248 120000 12368
rect 0 10888 800 11008
rect 119200 9528 120000 9648
rect 0 9256 800 9376
rect 0 7624 800 7744
rect 119200 6808 120000 6928
rect 0 5992 800 6112
rect 0 4360 800 4480
rect 119200 4088 120000 4208
rect 119200 1368 120000 1488
<< obsm3 >>
rect 798 115808 119219 117537
rect 798 115536 119120 115808
rect 880 115528 119120 115536
rect 880 115256 119219 115528
rect 798 113904 119219 115256
rect 880 113624 119219 113904
rect 798 113088 119219 113624
rect 798 112808 119120 113088
rect 798 112272 119219 112808
rect 880 111992 119219 112272
rect 798 110640 119219 111992
rect 880 110368 119219 110640
rect 880 110360 119120 110368
rect 798 110088 119120 110360
rect 798 109008 119219 110088
rect 880 108728 119219 109008
rect 798 107648 119219 108728
rect 798 107376 119120 107648
rect 880 107368 119120 107376
rect 880 107096 119219 107368
rect 798 105744 119219 107096
rect 880 105464 119219 105744
rect 798 104928 119219 105464
rect 798 104648 119120 104928
rect 798 104112 119219 104648
rect 880 103832 119219 104112
rect 798 102480 119219 103832
rect 880 102208 119219 102480
rect 880 102200 119120 102208
rect 798 101928 119120 102200
rect 798 100848 119219 101928
rect 880 100568 119219 100848
rect 798 99488 119219 100568
rect 798 99216 119120 99488
rect 880 99208 119120 99216
rect 880 98936 119219 99208
rect 798 97584 119219 98936
rect 880 97304 119219 97584
rect 798 96768 119219 97304
rect 798 96488 119120 96768
rect 798 95952 119219 96488
rect 880 95672 119219 95952
rect 798 94320 119219 95672
rect 880 94048 119219 94320
rect 880 94040 119120 94048
rect 798 93768 119120 94040
rect 798 92688 119219 93768
rect 880 92408 119219 92688
rect 798 91328 119219 92408
rect 798 91056 119120 91328
rect 880 91048 119120 91056
rect 880 90776 119219 91048
rect 798 89424 119219 90776
rect 880 89144 119219 89424
rect 798 88608 119219 89144
rect 798 88328 119120 88608
rect 798 87792 119219 88328
rect 880 87512 119219 87792
rect 798 86160 119219 87512
rect 880 85888 119219 86160
rect 880 85880 119120 85888
rect 798 85608 119120 85880
rect 798 84528 119219 85608
rect 880 84248 119219 84528
rect 798 83168 119219 84248
rect 798 82896 119120 83168
rect 880 82888 119120 82896
rect 880 82616 119219 82888
rect 798 81264 119219 82616
rect 880 80984 119219 81264
rect 798 80448 119219 80984
rect 798 80168 119120 80448
rect 798 79632 119219 80168
rect 880 79352 119219 79632
rect 798 78000 119219 79352
rect 880 77728 119219 78000
rect 880 77720 119120 77728
rect 798 77448 119120 77720
rect 798 76368 119219 77448
rect 880 76088 119219 76368
rect 798 75008 119219 76088
rect 798 74736 119120 75008
rect 880 74728 119120 74736
rect 880 74456 119219 74728
rect 798 73104 119219 74456
rect 880 72824 119219 73104
rect 798 72288 119219 72824
rect 798 72008 119120 72288
rect 798 71472 119219 72008
rect 880 71192 119219 71472
rect 798 69840 119219 71192
rect 880 69568 119219 69840
rect 880 69560 119120 69568
rect 798 69288 119120 69560
rect 798 68208 119219 69288
rect 880 67928 119219 68208
rect 798 66848 119219 67928
rect 798 66576 119120 66848
rect 880 66568 119120 66576
rect 880 66296 119219 66568
rect 798 64944 119219 66296
rect 880 64664 119219 64944
rect 798 64128 119219 64664
rect 798 63848 119120 64128
rect 798 63312 119219 63848
rect 880 63032 119219 63312
rect 798 61680 119219 63032
rect 880 61408 119219 61680
rect 880 61400 119120 61408
rect 798 61128 119120 61400
rect 798 60048 119219 61128
rect 880 59768 119219 60048
rect 798 58688 119219 59768
rect 798 58416 119120 58688
rect 880 58408 119120 58416
rect 880 58136 119219 58408
rect 798 56784 119219 58136
rect 880 56504 119219 56784
rect 798 55968 119219 56504
rect 798 55688 119120 55968
rect 798 55152 119219 55688
rect 880 54872 119219 55152
rect 798 53520 119219 54872
rect 880 53248 119219 53520
rect 880 53240 119120 53248
rect 798 52968 119120 53240
rect 798 51888 119219 52968
rect 880 51608 119219 51888
rect 798 50528 119219 51608
rect 798 50256 119120 50528
rect 880 50248 119120 50256
rect 880 49976 119219 50248
rect 798 48624 119219 49976
rect 880 48344 119219 48624
rect 798 47808 119219 48344
rect 798 47528 119120 47808
rect 798 46992 119219 47528
rect 880 46712 119219 46992
rect 798 45360 119219 46712
rect 880 45088 119219 45360
rect 880 45080 119120 45088
rect 798 44808 119120 45080
rect 798 43728 119219 44808
rect 880 43448 119219 43728
rect 798 42368 119219 43448
rect 798 42096 119120 42368
rect 880 42088 119120 42096
rect 880 41816 119219 42088
rect 798 40464 119219 41816
rect 880 40184 119219 40464
rect 798 39648 119219 40184
rect 798 39368 119120 39648
rect 798 38832 119219 39368
rect 880 38552 119219 38832
rect 798 37200 119219 38552
rect 880 36928 119219 37200
rect 880 36920 119120 36928
rect 798 36648 119120 36920
rect 798 35568 119219 36648
rect 880 35288 119219 35568
rect 798 34208 119219 35288
rect 798 33936 119120 34208
rect 880 33928 119120 33936
rect 880 33656 119219 33928
rect 798 32304 119219 33656
rect 880 32024 119219 32304
rect 798 31488 119219 32024
rect 798 31208 119120 31488
rect 798 30672 119219 31208
rect 880 30392 119219 30672
rect 798 29040 119219 30392
rect 880 28768 119219 29040
rect 880 28760 119120 28768
rect 798 28488 119120 28760
rect 798 27408 119219 28488
rect 880 27128 119219 27408
rect 798 26048 119219 27128
rect 798 25776 119120 26048
rect 880 25768 119120 25776
rect 880 25496 119219 25768
rect 798 24144 119219 25496
rect 880 23864 119219 24144
rect 798 23328 119219 23864
rect 798 23048 119120 23328
rect 798 22512 119219 23048
rect 880 22232 119219 22512
rect 798 20880 119219 22232
rect 880 20608 119219 20880
rect 880 20600 119120 20608
rect 798 20328 119120 20600
rect 798 19248 119219 20328
rect 880 18968 119219 19248
rect 798 17888 119219 18968
rect 798 17616 119120 17888
rect 880 17608 119120 17616
rect 880 17336 119219 17608
rect 798 15984 119219 17336
rect 880 15704 119219 15984
rect 798 15168 119219 15704
rect 798 14888 119120 15168
rect 798 14352 119219 14888
rect 880 14072 119219 14352
rect 798 12720 119219 14072
rect 880 12448 119219 12720
rect 880 12440 119120 12448
rect 798 12168 119120 12440
rect 798 11088 119219 12168
rect 880 10808 119219 11088
rect 798 9728 119219 10808
rect 798 9456 119120 9728
rect 880 9448 119120 9456
rect 880 9176 119219 9448
rect 798 7824 119219 9176
rect 880 7544 119219 7824
rect 798 7008 119219 7544
rect 798 6728 119120 7008
rect 798 6192 119219 6728
rect 880 5912 119219 6192
rect 798 4560 119219 5912
rect 880 4288 119219 4560
rect 880 4280 119120 4288
rect 798 4008 119120 4280
rect 798 1568 119219 4008
rect 798 1395 119120 1568
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 3187 3027 4128 117197
rect 4608 3027 19488 117197
rect 19968 3027 34848 117197
rect 35328 3027 50208 117197
rect 50688 3027 65568 117197
rect 66048 3027 80928 117197
rect 81408 3027 96288 117197
rect 96768 3027 111648 117197
rect 112128 3027 117149 117197
<< labels >>
rlabel metal2 s 29918 119200 29974 120000 6 clk_i
port 1 nsew signal input
rlabel metal3 s 119200 93848 120000 93968 6 enable_i
port 2 nsew signal input
rlabel metal3 s 119200 118328 120000 118448 6 fb_i
port 3 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 hsync_o
port 4 nsew signal output
rlabel metal3 s 119200 1368 120000 1488 6 mport_i[0]
port 5 nsew signal input
rlabel metal3 s 119200 28568 120000 28688 6 mport_i[10]
port 6 nsew signal input
rlabel metal3 s 119200 31288 120000 31408 6 mport_i[11]
port 7 nsew signal input
rlabel metal3 s 119200 34008 120000 34128 6 mport_i[12]
port 8 nsew signal input
rlabel metal3 s 119200 36728 120000 36848 6 mport_i[13]
port 9 nsew signal input
rlabel metal3 s 119200 39448 120000 39568 6 mport_i[14]
port 10 nsew signal input
rlabel metal3 s 119200 42168 120000 42288 6 mport_i[15]
port 11 nsew signal input
rlabel metal3 s 119200 44888 120000 45008 6 mport_i[16]
port 12 nsew signal input
rlabel metal3 s 119200 47608 120000 47728 6 mport_i[17]
port 13 nsew signal input
rlabel metal3 s 119200 50328 120000 50448 6 mport_i[18]
port 14 nsew signal input
rlabel metal3 s 119200 53048 120000 53168 6 mport_i[19]
port 15 nsew signal input
rlabel metal3 s 119200 4088 120000 4208 6 mport_i[1]
port 16 nsew signal input
rlabel metal3 s 119200 55768 120000 55888 6 mport_i[20]
port 17 nsew signal input
rlabel metal3 s 119200 58488 120000 58608 6 mport_i[21]
port 18 nsew signal input
rlabel metal3 s 119200 61208 120000 61328 6 mport_i[22]
port 19 nsew signal input
rlabel metal3 s 119200 63928 120000 64048 6 mport_i[23]
port 20 nsew signal input
rlabel metal3 s 119200 66648 120000 66768 6 mport_i[24]
port 21 nsew signal input
rlabel metal3 s 119200 69368 120000 69488 6 mport_i[25]
port 22 nsew signal input
rlabel metal3 s 119200 72088 120000 72208 6 mport_i[26]
port 23 nsew signal input
rlabel metal3 s 119200 74808 120000 74928 6 mport_i[27]
port 24 nsew signal input
rlabel metal3 s 119200 77528 120000 77648 6 mport_i[28]
port 25 nsew signal input
rlabel metal3 s 119200 80248 120000 80368 6 mport_i[29]
port 26 nsew signal input
rlabel metal3 s 119200 6808 120000 6928 6 mport_i[2]
port 27 nsew signal input
rlabel metal3 s 119200 82968 120000 83088 6 mport_i[30]
port 28 nsew signal input
rlabel metal3 s 119200 85688 120000 85808 6 mport_i[31]
port 29 nsew signal input
rlabel metal3 s 119200 88408 120000 88528 6 mport_i[32]
port 30 nsew signal input
rlabel metal3 s 119200 91128 120000 91248 6 mport_i[33]
port 31 nsew signal input
rlabel metal3 s 119200 9528 120000 9648 6 mport_i[3]
port 32 nsew signal input
rlabel metal3 s 119200 12248 120000 12368 6 mport_i[4]
port 33 nsew signal input
rlabel metal3 s 119200 14968 120000 15088 6 mport_i[5]
port 34 nsew signal input
rlabel metal3 s 119200 17688 120000 17808 6 mport_i[6]
port 35 nsew signal input
rlabel metal3 s 119200 20408 120000 20528 6 mport_i[7]
port 36 nsew signal input
rlabel metal3 s 119200 23128 120000 23248 6 mport_i[8]
port 37 nsew signal input
rlabel metal3 s 119200 25848 120000 25968 6 mport_i[9]
port 38 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 mport_o[0]
port 39 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 mport_o[10]
port 40 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 mport_o[11]
port 41 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 mport_o[12]
port 42 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 mport_o[13]
port 43 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 mport_o[14]
port 44 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 mport_o[15]
port 45 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 mport_o[16]
port 46 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 mport_o[17]
port 47 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 mport_o[18]
port 48 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 mport_o[19]
port 49 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 mport_o[1]
port 50 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 mport_o[20]
port 51 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 mport_o[21]
port 52 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 mport_o[22]
port 53 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 mport_o[23]
port 54 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 mport_o[24]
port 55 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 mport_o[25]
port 56 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 mport_o[26]
port 57 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 mport_o[27]
port 58 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 mport_o[28]
port 59 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 mport_o[29]
port 60 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 mport_o[2]
port 61 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 mport_o[30]
port 62 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 mport_o[31]
port 63 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 mport_o[32]
port 64 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 mport_o[33]
port 65 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 mport_o[34]
port 66 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 mport_o[35]
port 67 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 mport_o[36]
port 68 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 mport_o[37]
port 69 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 mport_o[38]
port 70 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 mport_o[39]
port 71 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 mport_o[3]
port 72 nsew signal output
rlabel metal3 s 0 69640 800 69760 6 mport_o[40]
port 73 nsew signal output
rlabel metal3 s 0 71272 800 71392 6 mport_o[41]
port 74 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 mport_o[42]
port 75 nsew signal output
rlabel metal3 s 0 74536 800 74656 6 mport_o[43]
port 76 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 mport_o[44]
port 77 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 mport_o[45]
port 78 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 mport_o[46]
port 79 nsew signal output
rlabel metal3 s 0 81064 800 81184 6 mport_o[47]
port 80 nsew signal output
rlabel metal3 s 0 82696 800 82816 6 mport_o[48]
port 81 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 mport_o[49]
port 82 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 mport_o[4]
port 83 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 mport_o[50]
port 84 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 mport_o[51]
port 85 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 mport_o[52]
port 86 nsew signal output
rlabel metal3 s 0 90856 800 90976 6 mport_o[53]
port 87 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 mport_o[54]
port 88 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 mport_o[55]
port 89 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 mport_o[56]
port 90 nsew signal output
rlabel metal3 s 0 97384 800 97504 6 mport_o[57]
port 91 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 mport_o[58]
port 92 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 mport_o[59]
port 93 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 mport_o[5]
port 94 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 mport_o[60]
port 95 nsew signal output
rlabel metal3 s 0 103912 800 104032 6 mport_o[61]
port 96 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 mport_o[62]
port 97 nsew signal output
rlabel metal3 s 0 107176 800 107296 6 mport_o[63]
port 98 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 mport_o[64]
port 99 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 mport_o[65]
port 100 nsew signal output
rlabel metal3 s 0 112072 800 112192 6 mport_o[66]
port 101 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 mport_o[67]
port 102 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 mport_o[68]
port 103 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 mport_o[6]
port 104 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 mport_o[7]
port 105 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 mport_o[8]
port 106 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 mport_o[9]
port 107 nsew signal output
rlabel metal2 s 89902 119200 89958 120000 6 nrst_i
port 108 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 pixel_o[0]
port 109 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 pixel_o[1]
port 110 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 pixel_o[2]
port 111 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 pixel_o[3]
port 112 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 pixel_o[4]
port 113 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 pixel_o[5]
port 114 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 pixel_o[6]
port 115 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 pixel_o[7]
port 116 nsew signal output
rlabel metal3 s 119200 96568 120000 96688 6 prescaler_i[0]
port 117 nsew signal input
rlabel metal3 s 119200 99288 120000 99408 6 prescaler_i[1]
port 118 nsew signal input
rlabel metal3 s 119200 102008 120000 102128 6 prescaler_i[2]
port 119 nsew signal input
rlabel metal3 s 119200 104728 120000 104848 6 prescaler_i[3]
port 120 nsew signal input
rlabel metal3 s 119200 107448 120000 107568 6 resolution_i[0]
port 121 nsew signal input
rlabel metal3 s 119200 110168 120000 110288 6 resolution_i[1]
port 122 nsew signal input
rlabel metal3 s 119200 112888 120000 113008 6 resolution_i[2]
port 123 nsew signal input
rlabel metal3 s 119200 115608 120000 115728 6 resolution_i[3]
port 124 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 125 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 125 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 125 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 125 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 126 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 126 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 126 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 126 nsew ground bidirectional
rlabel metal2 s 113730 0 113786 800 6 vsync_o
port 127 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 55442140
string GDS_FILE /home/mdrobot7/sdmay26-24/openlane/vga/runs/25_10_21_16_39/results/signoff/vga.magic.gds
string GDS_START 994976
<< end >>

