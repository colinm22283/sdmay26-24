VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bary_pipe_m
  CLASS BLOCK ;
  FOREIGN bary_pipe_m ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN busy_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END busy_o
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END clk_i
  PIN discard_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END discard_o
  PIN init_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END init_o
  PIN mstream_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 4.120 800.000 4.720 ;
    END
  END mstream_i
  PIN mstream_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 10.920 800.000 11.520 ;
    END
  END mstream_o[0]
  PIN mstream_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 690.920 800.000 691.520 ;
    END
  END mstream_o[100]
  PIN mstream_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 697.720 800.000 698.320 ;
    END
  END mstream_o[101]
  PIN mstream_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 704.520 800.000 705.120 ;
    END
  END mstream_o[102]
  PIN mstream_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 711.320 800.000 711.920 ;
    END
  END mstream_o[103]
  PIN mstream_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 718.120 800.000 718.720 ;
    END
  END mstream_o[104]
  PIN mstream_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 724.920 800.000 725.520 ;
    END
  END mstream_o[105]
  PIN mstream_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 731.720 800.000 732.320 ;
    END
  END mstream_o[106]
  PIN mstream_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 738.520 800.000 739.120 ;
    END
  END mstream_o[107]
  PIN mstream_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 745.320 800.000 745.920 ;
    END
  END mstream_o[108]
  PIN mstream_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 752.120 800.000 752.720 ;
    END
  END mstream_o[109]
  PIN mstream_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 78.920 800.000 79.520 ;
    END
  END mstream_o[10]
  PIN mstream_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 758.920 800.000 759.520 ;
    END
  END mstream_o[110]
  PIN mstream_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 765.720 800.000 766.320 ;
    END
  END mstream_o[111]
  PIN mstream_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 772.520 800.000 773.120 ;
    END
  END mstream_o[112]
  PIN mstream_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 779.320 800.000 779.920 ;
    END
  END mstream_o[113]
  PIN mstream_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 6.976800 ;
    PORT
      LAYER met3 ;
        RECT 796.000 786.120 800.000 786.720 ;
    END
  END mstream_o[114]
  PIN mstream_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 792.920 800.000 793.520 ;
    END
  END mstream_o[115]
  PIN mstream_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 85.720 800.000 86.320 ;
    END
  END mstream_o[11]
  PIN mstream_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 92.520 800.000 93.120 ;
    END
  END mstream_o[12]
  PIN mstream_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 99.320 800.000 99.920 ;
    END
  END mstream_o[13]
  PIN mstream_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 106.120 800.000 106.720 ;
    END
  END mstream_o[14]
  PIN mstream_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 112.920 800.000 113.520 ;
    END
  END mstream_o[15]
  PIN mstream_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 119.720 800.000 120.320 ;
    END
  END mstream_o[16]
  PIN mstream_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 126.520 800.000 127.120 ;
    END
  END mstream_o[17]
  PIN mstream_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 133.320 800.000 133.920 ;
    END
  END mstream_o[18]
  PIN mstream_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 140.120 800.000 140.720 ;
    END
  END mstream_o[19]
  PIN mstream_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 17.720 800.000 18.320 ;
    END
  END mstream_o[1]
  PIN mstream_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 146.920 800.000 147.520 ;
    END
  END mstream_o[20]
  PIN mstream_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 153.720 800.000 154.320 ;
    END
  END mstream_o[21]
  PIN mstream_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 160.520 800.000 161.120 ;
    END
  END mstream_o[22]
  PIN mstream_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 167.320 800.000 167.920 ;
    END
  END mstream_o[23]
  PIN mstream_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 174.120 800.000 174.720 ;
    END
  END mstream_o[24]
  PIN mstream_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 180.920 800.000 181.520 ;
    END
  END mstream_o[25]
  PIN mstream_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 187.720 800.000 188.320 ;
    END
  END mstream_o[26]
  PIN mstream_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 194.520 800.000 195.120 ;
    END
  END mstream_o[27]
  PIN mstream_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 201.320 800.000 201.920 ;
    END
  END mstream_o[28]
  PIN mstream_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 208.120 800.000 208.720 ;
    END
  END mstream_o[29]
  PIN mstream_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 24.520 800.000 25.120 ;
    END
  END mstream_o[2]
  PIN mstream_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 214.920 800.000 215.520 ;
    END
  END mstream_o[30]
  PIN mstream_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 221.720 800.000 222.320 ;
    END
  END mstream_o[31]
  PIN mstream_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 228.520 800.000 229.120 ;
    END
  END mstream_o[32]
  PIN mstream_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 235.320 800.000 235.920 ;
    END
  END mstream_o[33]
  PIN mstream_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 242.120 800.000 242.720 ;
    END
  END mstream_o[34]
  PIN mstream_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 248.920 800.000 249.520 ;
    END
  END mstream_o[35]
  PIN mstream_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 255.720 800.000 256.320 ;
    END
  END mstream_o[36]
  PIN mstream_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 262.520 800.000 263.120 ;
    END
  END mstream_o[37]
  PIN mstream_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 269.320 800.000 269.920 ;
    END
  END mstream_o[38]
  PIN mstream_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 276.120 800.000 276.720 ;
    END
  END mstream_o[39]
  PIN mstream_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 31.320 800.000 31.920 ;
    END
  END mstream_o[3]
  PIN mstream_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 282.920 800.000 283.520 ;
    END
  END mstream_o[40]
  PIN mstream_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 289.720 800.000 290.320 ;
    END
  END mstream_o[41]
  PIN mstream_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 296.520 800.000 297.120 ;
    END
  END mstream_o[42]
  PIN mstream_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 303.320 800.000 303.920 ;
    END
  END mstream_o[43]
  PIN mstream_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 310.120 800.000 310.720 ;
    END
  END mstream_o[44]
  PIN mstream_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 316.920 800.000 317.520 ;
    END
  END mstream_o[45]
  PIN mstream_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 323.720 800.000 324.320 ;
    END
  END mstream_o[46]
  PIN mstream_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 330.520 800.000 331.120 ;
    END
  END mstream_o[47]
  PIN mstream_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 337.320 800.000 337.920 ;
    END
  END mstream_o[48]
  PIN mstream_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 344.120 800.000 344.720 ;
    END
  END mstream_o[49]
  PIN mstream_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 38.120 800.000 38.720 ;
    END
  END mstream_o[4]
  PIN mstream_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 350.920 800.000 351.520 ;
    END
  END mstream_o[50]
  PIN mstream_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 357.720 800.000 358.320 ;
    END
  END mstream_o[51]
  PIN mstream_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 364.520 800.000 365.120 ;
    END
  END mstream_o[52]
  PIN mstream_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 371.320 800.000 371.920 ;
    END
  END mstream_o[53]
  PIN mstream_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 378.120 800.000 378.720 ;
    END
  END mstream_o[54]
  PIN mstream_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 384.920 800.000 385.520 ;
    END
  END mstream_o[55]
  PIN mstream_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 391.720 800.000 392.320 ;
    END
  END mstream_o[56]
  PIN mstream_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 398.520 800.000 399.120 ;
    END
  END mstream_o[57]
  PIN mstream_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 405.320 800.000 405.920 ;
    END
  END mstream_o[58]
  PIN mstream_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 412.120 800.000 412.720 ;
    END
  END mstream_o[59]
  PIN mstream_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 44.920 800.000 45.520 ;
    END
  END mstream_o[5]
  PIN mstream_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 418.920 800.000 419.520 ;
    END
  END mstream_o[60]
  PIN mstream_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 425.720 800.000 426.320 ;
    END
  END mstream_o[61]
  PIN mstream_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 432.520 800.000 433.120 ;
    END
  END mstream_o[62]
  PIN mstream_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 439.320 800.000 439.920 ;
    END
  END mstream_o[63]
  PIN mstream_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 446.120 800.000 446.720 ;
    END
  END mstream_o[64]
  PIN mstream_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 452.920 800.000 453.520 ;
    END
  END mstream_o[65]
  PIN mstream_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 459.720 800.000 460.320 ;
    END
  END mstream_o[66]
  PIN mstream_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 466.520 800.000 467.120 ;
    END
  END mstream_o[67]
  PIN mstream_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 473.320 800.000 473.920 ;
    END
  END mstream_o[68]
  PIN mstream_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 480.120 800.000 480.720 ;
    END
  END mstream_o[69]
  PIN mstream_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 51.720 800.000 52.320 ;
    END
  END mstream_o[6]
  PIN mstream_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 486.920 800.000 487.520 ;
    END
  END mstream_o[70]
  PIN mstream_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 493.720 800.000 494.320 ;
    END
  END mstream_o[71]
  PIN mstream_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 500.520 800.000 501.120 ;
    END
  END mstream_o[72]
  PIN mstream_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 507.320 800.000 507.920 ;
    END
  END mstream_o[73]
  PIN mstream_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 514.120 800.000 514.720 ;
    END
  END mstream_o[74]
  PIN mstream_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 520.920 800.000 521.520 ;
    END
  END mstream_o[75]
  PIN mstream_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 527.720 800.000 528.320 ;
    END
  END mstream_o[76]
  PIN mstream_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 534.520 800.000 535.120 ;
    END
  END mstream_o[77]
  PIN mstream_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 541.320 800.000 541.920 ;
    END
  END mstream_o[78]
  PIN mstream_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 548.120 800.000 548.720 ;
    END
  END mstream_o[79]
  PIN mstream_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 58.520 800.000 59.120 ;
    END
  END mstream_o[7]
  PIN mstream_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 554.920 800.000 555.520 ;
    END
  END mstream_o[80]
  PIN mstream_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 561.720 800.000 562.320 ;
    END
  END mstream_o[81]
  PIN mstream_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 568.520 800.000 569.120 ;
    END
  END mstream_o[82]
  PIN mstream_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 575.320 800.000 575.920 ;
    END
  END mstream_o[83]
  PIN mstream_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 582.120 800.000 582.720 ;
    END
  END mstream_o[84]
  PIN mstream_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 588.920 800.000 589.520 ;
    END
  END mstream_o[85]
  PIN mstream_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 595.720 800.000 596.320 ;
    END
  END mstream_o[86]
  PIN mstream_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 602.520 800.000 603.120 ;
    END
  END mstream_o[87]
  PIN mstream_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 609.320 800.000 609.920 ;
    END
  END mstream_o[88]
  PIN mstream_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 616.120 800.000 616.720 ;
    END
  END mstream_o[89]
  PIN mstream_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 65.320 800.000 65.920 ;
    END
  END mstream_o[8]
  PIN mstream_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 622.920 800.000 623.520 ;
    END
  END mstream_o[90]
  PIN mstream_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 629.720 800.000 630.320 ;
    END
  END mstream_o[91]
  PIN mstream_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 636.520 800.000 637.120 ;
    END
  END mstream_o[92]
  PIN mstream_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 643.320 800.000 643.920 ;
    END
  END mstream_o[93]
  PIN mstream_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 13.062600 ;
    PORT
      LAYER met3 ;
        RECT 796.000 650.120 800.000 650.720 ;
    END
  END mstream_o[94]
  PIN mstream_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 656.920 800.000 657.520 ;
    END
  END mstream_o[95]
  PIN mstream_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 663.720 800.000 664.320 ;
    END
  END mstream_o[96]
  PIN mstream_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 670.520 800.000 671.120 ;
    END
  END mstream_o[97]
  PIN mstream_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 677.320 800.000 677.920 ;
    END
  END mstream_o[98]
  PIN mstream_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 684.120 800.000 684.720 ;
    END
  END mstream_o[99]
  PIN mstream_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 72.120 800.000 72.720 ;
    END
  END mstream_o[9]
  PIN nrst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END nrst_i
  PIN run_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END run_i
  PIN sstream_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END sstream_i[0]
  PIN sstream_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 10.432799 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END sstream_i[10]
  PIN sstream_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END sstream_i[11]
  PIN sstream_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END sstream_i[12]
  PIN sstream_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END sstream_i[13]
  PIN sstream_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END sstream_i[14]
  PIN sstream_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END sstream_i[15]
  PIN sstream_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END sstream_i[16]
  PIN sstream_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END sstream_i[17]
  PIN sstream_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END sstream_i[18]
  PIN sstream_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END sstream_i[19]
  PIN sstream_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END sstream_i[1]
  PIN sstream_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END sstream_i[2]
  PIN sstream_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END sstream_i[3]
  PIN sstream_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 6.520500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END sstream_i[4]
  PIN sstream_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END sstream_i[5]
  PIN sstream_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END sstream_i[6]
  PIN sstream_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END sstream_i[7]
  PIN sstream_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END sstream_i[8]
  PIN sstream_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END sstream_i[9]
  PIN sstream_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.858500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END sstream_o
  PIN v0x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END v0x[0]
  PIN v0x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END v0x[10]
  PIN v0x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END v0x[11]
  PIN v0x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END v0x[12]
  PIN v0x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END v0x[13]
  PIN v0x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END v0x[14]
  PIN v0x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END v0x[15]
  PIN v0x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END v0x[16]
  PIN v0x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END v0x[17]
  PIN v0x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END v0x[18]
  PIN v0x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END v0x[19]
  PIN v0x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END v0x[1]
  PIN v0x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END v0x[20]
  PIN v0x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END v0x[21]
  PIN v0x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END v0x[22]
  PIN v0x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END v0x[23]
  PIN v0x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END v0x[24]
  PIN v0x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END v0x[25]
  PIN v0x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END v0x[26]
  PIN v0x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END v0x[27]
  PIN v0x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END v0x[28]
  PIN v0x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END v0x[29]
  PIN v0x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END v0x[2]
  PIN v0x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END v0x[30]
  PIN v0x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END v0x[31]
  PIN v0x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END v0x[3]
  PIN v0x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END v0x[4]
  PIN v0x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END v0x[5]
  PIN v0x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END v0x[6]
  PIN v0x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END v0x[7]
  PIN v0x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END v0x[8]
  PIN v0x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END v0x[9]
  PIN v0y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END v0y[0]
  PIN v0y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END v0y[10]
  PIN v0y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END v0y[11]
  PIN v0y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END v0y[12]
  PIN v0y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END v0y[13]
  PIN v0y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END v0y[14]
  PIN v0y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END v0y[15]
  PIN v0y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END v0y[16]
  PIN v0y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END v0y[17]
  PIN v0y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END v0y[18]
  PIN v0y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END v0y[19]
  PIN v0y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END v0y[1]
  PIN v0y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END v0y[20]
  PIN v0y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END v0y[21]
  PIN v0y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END v0y[22]
  PIN v0y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END v0y[23]
  PIN v0y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END v0y[24]
  PIN v0y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END v0y[25]
  PIN v0y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END v0y[26]
  PIN v0y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END v0y[27]
  PIN v0y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 4.000 ;
    END
  END v0y[28]
  PIN v0y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END v0y[29]
  PIN v0y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END v0y[2]
  PIN v0y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END v0y[30]
  PIN v0y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END v0y[31]
  PIN v0y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END v0y[3]
  PIN v0y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END v0y[4]
  PIN v0y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END v0y[5]
  PIN v0y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END v0y[6]
  PIN v0y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END v0y[7]
  PIN v0y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END v0y[8]
  PIN v0y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END v0y[9]
  PIN v0z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END v0z[0]
  PIN v0z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END v0z[10]
  PIN v0z[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END v0z[11]
  PIN v0z[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END v0z[12]
  PIN v0z[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END v0z[13]
  PIN v0z[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END v0z[14]
  PIN v0z[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END v0z[15]
  PIN v0z[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END v0z[16]
  PIN v0z[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END v0z[17]
  PIN v0z[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END v0z[18]
  PIN v0z[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END v0z[19]
  PIN v0z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END v0z[1]
  PIN v0z[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END v0z[20]
  PIN v0z[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END v0z[21]
  PIN v0z[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END v0z[22]
  PIN v0z[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END v0z[23]
  PIN v0z[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END v0z[24]
  PIN v0z[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END v0z[25]
  PIN v0z[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END v0z[26]
  PIN v0z[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END v0z[27]
  PIN v0z[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END v0z[28]
  PIN v0z[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END v0z[29]
  PIN v0z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END v0z[2]
  PIN v0z[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END v0z[30]
  PIN v0z[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END v0z[31]
  PIN v0z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END v0z[3]
  PIN v0z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END v0z[4]
  PIN v0z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END v0z[5]
  PIN v0z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END v0z[6]
  PIN v0z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END v0z[7]
  PIN v0z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END v0z[8]
  PIN v0z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END v0z[9]
  PIN v1x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END v1x[0]
  PIN v1x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END v1x[10]
  PIN v1x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END v1x[11]
  PIN v1x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END v1x[12]
  PIN v1x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END v1x[13]
  PIN v1x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END v1x[14]
  PIN v1x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END v1x[15]
  PIN v1x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END v1x[16]
  PIN v1x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END v1x[17]
  PIN v1x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END v1x[18]
  PIN v1x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END v1x[19]
  PIN v1x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END v1x[1]
  PIN v1x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END v1x[20]
  PIN v1x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END v1x[21]
  PIN v1x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END v1x[22]
  PIN v1x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END v1x[23]
  PIN v1x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END v1x[24]
  PIN v1x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END v1x[25]
  PIN v1x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END v1x[26]
  PIN v1x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END v1x[27]
  PIN v1x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END v1x[28]
  PIN v1x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END v1x[29]
  PIN v1x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END v1x[2]
  PIN v1x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END v1x[30]
  PIN v1x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END v1x[31]
  PIN v1x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END v1x[3]
  PIN v1x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END v1x[4]
  PIN v1x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END v1x[5]
  PIN v1x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END v1x[6]
  PIN v1x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END v1x[7]
  PIN v1x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END v1x[8]
  PIN v1x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END v1x[9]
  PIN v1y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END v1y[0]
  PIN v1y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END v1y[10]
  PIN v1y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END v1y[11]
  PIN v1y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END v1y[12]
  PIN v1y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END v1y[13]
  PIN v1y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END v1y[14]
  PIN v1y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END v1y[15]
  PIN v1y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END v1y[16]
  PIN v1y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END v1y[17]
  PIN v1y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END v1y[18]
  PIN v1y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END v1y[19]
  PIN v1y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END v1y[1]
  PIN v1y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END v1y[20]
  PIN v1y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END v1y[21]
  PIN v1y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END v1y[22]
  PIN v1y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END v1y[23]
  PIN v1y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END v1y[24]
  PIN v1y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END v1y[25]
  PIN v1y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END v1y[26]
  PIN v1y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END v1y[27]
  PIN v1y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END v1y[28]
  PIN v1y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END v1y[29]
  PIN v1y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END v1y[2]
  PIN v1y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END v1y[30]
  PIN v1y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END v1y[31]
  PIN v1y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END v1y[3]
  PIN v1y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END v1y[4]
  PIN v1y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END v1y[5]
  PIN v1y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END v1y[6]
  PIN v1y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END v1y[7]
  PIN v1y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END v1y[8]
  PIN v1y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END v1y[9]
  PIN v1z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END v1z[0]
  PIN v1z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END v1z[10]
  PIN v1z[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END v1z[11]
  PIN v1z[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END v1z[12]
  PIN v1z[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END v1z[13]
  PIN v1z[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END v1z[14]
  PIN v1z[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END v1z[15]
  PIN v1z[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END v1z[16]
  PIN v1z[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END v1z[17]
  PIN v1z[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END v1z[18]
  PIN v1z[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END v1z[19]
  PIN v1z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END v1z[1]
  PIN v1z[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END v1z[20]
  PIN v1z[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END v1z[21]
  PIN v1z[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END v1z[22]
  PIN v1z[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END v1z[23]
  PIN v1z[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END v1z[24]
  PIN v1z[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END v1z[25]
  PIN v1z[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END v1z[26]
  PIN v1z[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END v1z[27]
  PIN v1z[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END v1z[28]
  PIN v1z[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END v1z[29]
  PIN v1z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END v1z[2]
  PIN v1z[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END v1z[30]
  PIN v1z[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END v1z[31]
  PIN v1z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END v1z[3]
  PIN v1z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END v1z[4]
  PIN v1z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END v1z[5]
  PIN v1z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END v1z[6]
  PIN v1z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END v1z[7]
  PIN v1z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END v1z[8]
  PIN v1z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END v1z[9]
  PIN v2x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END v2x[0]
  PIN v2x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END v2x[10]
  PIN v2x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END v2x[11]
  PIN v2x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END v2x[12]
  PIN v2x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END v2x[13]
  PIN v2x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END v2x[14]
  PIN v2x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END v2x[15]
  PIN v2x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END v2x[16]
  PIN v2x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END v2x[17]
  PIN v2x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END v2x[18]
  PIN v2x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END v2x[19]
  PIN v2x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END v2x[1]
  PIN v2x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END v2x[20]
  PIN v2x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END v2x[21]
  PIN v2x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END v2x[22]
  PIN v2x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END v2x[23]
  PIN v2x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END v2x[24]
  PIN v2x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END v2x[25]
  PIN v2x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END v2x[26]
  PIN v2x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END v2x[27]
  PIN v2x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END v2x[28]
  PIN v2x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END v2x[29]
  PIN v2x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END v2x[2]
  PIN v2x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END v2x[30]
  PIN v2x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END v2x[31]
  PIN v2x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END v2x[3]
  PIN v2x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END v2x[4]
  PIN v2x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END v2x[5]
  PIN v2x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END v2x[6]
  PIN v2x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END v2x[7]
  PIN v2x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END v2x[8]
  PIN v2x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END v2x[9]
  PIN v2y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END v2y[0]
  PIN v2y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END v2y[10]
  PIN v2y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END v2y[11]
  PIN v2y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END v2y[12]
  PIN v2y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END v2y[13]
  PIN v2y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END v2y[14]
  PIN v2y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END v2y[15]
  PIN v2y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END v2y[16]
  PIN v2y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END v2y[17]
  PIN v2y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END v2y[18]
  PIN v2y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END v2y[19]
  PIN v2y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END v2y[1]
  PIN v2y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END v2y[20]
  PIN v2y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END v2y[21]
  PIN v2y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END v2y[22]
  PIN v2y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END v2y[23]
  PIN v2y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END v2y[24]
  PIN v2y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END v2y[25]
  PIN v2y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END v2y[26]
  PIN v2y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 651.450 0.000 651.730 4.000 ;
    END
  END v2y[27]
  PIN v2y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END v2y[28]
  PIN v2y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END v2y[29]
  PIN v2y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END v2y[2]
  PIN v2y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END v2y[30]
  PIN v2y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END v2y[31]
  PIN v2y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END v2y[3]
  PIN v2y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END v2y[4]
  PIN v2y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END v2y[5]
  PIN v2y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END v2y[6]
  PIN v2y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END v2y[7]
  PIN v2y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END v2y[8]
  PIN v2y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END v2y[9]
  PIN v2z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END v2z[0]
  PIN v2z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END v2z[10]
  PIN v2z[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END v2z[11]
  PIN v2z[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END v2z[12]
  PIN v2z[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END v2z[13]
  PIN v2z[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END v2z[14]
  PIN v2z[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END v2z[15]
  PIN v2z[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END v2z[16]
  PIN v2z[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END v2z[17]
  PIN v2z[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END v2z[18]
  PIN v2z[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END v2z[19]
  PIN v2z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END v2z[1]
  PIN v2z[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END v2z[20]
  PIN v2z[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END v2z[21]
  PIN v2z[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END v2z[22]
  PIN v2z[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END v2z[23]
  PIN v2z[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END v2z[24]
  PIN v2z[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END v2z[25]
  PIN v2z[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END v2z[26]
  PIN v2z[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END v2z[27]
  PIN v2z[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END v2z[28]
  PIN v2z[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 4.000 ;
    END
  END v2z[29]
  PIN v2z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END v2z[2]
  PIN v2z[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END v2z[30]
  PIN v2z[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END v2z[31]
  PIN v2z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END v2z[3]
  PIN v2z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END v2z[4]
  PIN v2z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END v2z[5]
  PIN v2z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END v2z[6]
  PIN v2z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END v2z[7]
  PIN v2z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END v2z[8]
  PIN v2z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END v2z[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 788.885 ;
      LAYER met1 ;
        RECT 5.520 0.380 796.650 789.040 ;
      LAYER met2 ;
        RECT 17.110 4.280 796.620 793.405 ;
        RECT 17.110 0.155 62.370 4.280 ;
        RECT 63.210 0.155 64.670 4.280 ;
        RECT 65.510 0.155 66.970 4.280 ;
        RECT 67.810 0.155 69.270 4.280 ;
        RECT 70.110 0.155 71.570 4.280 ;
        RECT 72.410 0.155 73.870 4.280 ;
        RECT 74.710 0.155 76.170 4.280 ;
        RECT 77.010 0.155 78.470 4.280 ;
        RECT 79.310 0.155 80.770 4.280 ;
        RECT 81.610 0.155 83.070 4.280 ;
        RECT 83.910 0.155 85.370 4.280 ;
        RECT 86.210 0.155 87.670 4.280 ;
        RECT 88.510 0.155 89.970 4.280 ;
        RECT 90.810 0.155 92.270 4.280 ;
        RECT 93.110 0.155 94.570 4.280 ;
        RECT 95.410 0.155 96.870 4.280 ;
        RECT 97.710 0.155 99.170 4.280 ;
        RECT 100.010 0.155 101.470 4.280 ;
        RECT 102.310 0.155 103.770 4.280 ;
        RECT 104.610 0.155 106.070 4.280 ;
        RECT 106.910 0.155 108.370 4.280 ;
        RECT 109.210 0.155 110.670 4.280 ;
        RECT 111.510 0.155 112.970 4.280 ;
        RECT 113.810 0.155 115.270 4.280 ;
        RECT 116.110 0.155 117.570 4.280 ;
        RECT 118.410 0.155 119.870 4.280 ;
        RECT 120.710 0.155 122.170 4.280 ;
        RECT 123.010 0.155 124.470 4.280 ;
        RECT 125.310 0.155 126.770 4.280 ;
        RECT 127.610 0.155 129.070 4.280 ;
        RECT 129.910 0.155 131.370 4.280 ;
        RECT 132.210 0.155 133.670 4.280 ;
        RECT 134.510 0.155 135.970 4.280 ;
        RECT 136.810 0.155 138.270 4.280 ;
        RECT 139.110 0.155 140.570 4.280 ;
        RECT 141.410 0.155 142.870 4.280 ;
        RECT 143.710 0.155 145.170 4.280 ;
        RECT 146.010 0.155 147.470 4.280 ;
        RECT 148.310 0.155 149.770 4.280 ;
        RECT 150.610 0.155 152.070 4.280 ;
        RECT 152.910 0.155 154.370 4.280 ;
        RECT 155.210 0.155 156.670 4.280 ;
        RECT 157.510 0.155 158.970 4.280 ;
        RECT 159.810 0.155 161.270 4.280 ;
        RECT 162.110 0.155 163.570 4.280 ;
        RECT 164.410 0.155 165.870 4.280 ;
        RECT 166.710 0.155 168.170 4.280 ;
        RECT 169.010 0.155 170.470 4.280 ;
        RECT 171.310 0.155 172.770 4.280 ;
        RECT 173.610 0.155 175.070 4.280 ;
        RECT 175.910 0.155 177.370 4.280 ;
        RECT 178.210 0.155 179.670 4.280 ;
        RECT 180.510 0.155 181.970 4.280 ;
        RECT 182.810 0.155 184.270 4.280 ;
        RECT 185.110 0.155 186.570 4.280 ;
        RECT 187.410 0.155 188.870 4.280 ;
        RECT 189.710 0.155 191.170 4.280 ;
        RECT 192.010 0.155 193.470 4.280 ;
        RECT 194.310 0.155 195.770 4.280 ;
        RECT 196.610 0.155 198.070 4.280 ;
        RECT 198.910 0.155 200.370 4.280 ;
        RECT 201.210 0.155 202.670 4.280 ;
        RECT 203.510 0.155 204.970 4.280 ;
        RECT 205.810 0.155 207.270 4.280 ;
        RECT 208.110 0.155 209.570 4.280 ;
        RECT 210.410 0.155 211.870 4.280 ;
        RECT 212.710 0.155 214.170 4.280 ;
        RECT 215.010 0.155 216.470 4.280 ;
        RECT 217.310 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.070 4.280 ;
        RECT 221.910 0.155 223.370 4.280 ;
        RECT 224.210 0.155 225.670 4.280 ;
        RECT 226.510 0.155 227.970 4.280 ;
        RECT 228.810 0.155 230.270 4.280 ;
        RECT 231.110 0.155 232.570 4.280 ;
        RECT 233.410 0.155 234.870 4.280 ;
        RECT 235.710 0.155 237.170 4.280 ;
        RECT 238.010 0.155 239.470 4.280 ;
        RECT 240.310 0.155 241.770 4.280 ;
        RECT 242.610 0.155 244.070 4.280 ;
        RECT 244.910 0.155 246.370 4.280 ;
        RECT 247.210 0.155 248.670 4.280 ;
        RECT 249.510 0.155 250.970 4.280 ;
        RECT 251.810 0.155 253.270 4.280 ;
        RECT 254.110 0.155 255.570 4.280 ;
        RECT 256.410 0.155 257.870 4.280 ;
        RECT 258.710 0.155 260.170 4.280 ;
        RECT 261.010 0.155 262.470 4.280 ;
        RECT 263.310 0.155 264.770 4.280 ;
        RECT 265.610 0.155 267.070 4.280 ;
        RECT 267.910 0.155 269.370 4.280 ;
        RECT 270.210 0.155 271.670 4.280 ;
        RECT 272.510 0.155 273.970 4.280 ;
        RECT 274.810 0.155 276.270 4.280 ;
        RECT 277.110 0.155 278.570 4.280 ;
        RECT 279.410 0.155 280.870 4.280 ;
        RECT 281.710 0.155 283.170 4.280 ;
        RECT 284.010 0.155 285.470 4.280 ;
        RECT 286.310 0.155 287.770 4.280 ;
        RECT 288.610 0.155 290.070 4.280 ;
        RECT 290.910 0.155 292.370 4.280 ;
        RECT 293.210 0.155 294.670 4.280 ;
        RECT 295.510 0.155 296.970 4.280 ;
        RECT 297.810 0.155 299.270 4.280 ;
        RECT 300.110 0.155 301.570 4.280 ;
        RECT 302.410 0.155 303.870 4.280 ;
        RECT 304.710 0.155 306.170 4.280 ;
        RECT 307.010 0.155 308.470 4.280 ;
        RECT 309.310 0.155 310.770 4.280 ;
        RECT 311.610 0.155 313.070 4.280 ;
        RECT 313.910 0.155 315.370 4.280 ;
        RECT 316.210 0.155 317.670 4.280 ;
        RECT 318.510 0.155 319.970 4.280 ;
        RECT 320.810 0.155 322.270 4.280 ;
        RECT 323.110 0.155 324.570 4.280 ;
        RECT 325.410 0.155 326.870 4.280 ;
        RECT 327.710 0.155 329.170 4.280 ;
        RECT 330.010 0.155 331.470 4.280 ;
        RECT 332.310 0.155 333.770 4.280 ;
        RECT 334.610 0.155 336.070 4.280 ;
        RECT 336.910 0.155 338.370 4.280 ;
        RECT 339.210 0.155 340.670 4.280 ;
        RECT 341.510 0.155 342.970 4.280 ;
        RECT 343.810 0.155 345.270 4.280 ;
        RECT 346.110 0.155 347.570 4.280 ;
        RECT 348.410 0.155 349.870 4.280 ;
        RECT 350.710 0.155 352.170 4.280 ;
        RECT 353.010 0.155 354.470 4.280 ;
        RECT 355.310 0.155 356.770 4.280 ;
        RECT 357.610 0.155 359.070 4.280 ;
        RECT 359.910 0.155 361.370 4.280 ;
        RECT 362.210 0.155 363.670 4.280 ;
        RECT 364.510 0.155 365.970 4.280 ;
        RECT 366.810 0.155 368.270 4.280 ;
        RECT 369.110 0.155 370.570 4.280 ;
        RECT 371.410 0.155 372.870 4.280 ;
        RECT 373.710 0.155 375.170 4.280 ;
        RECT 376.010 0.155 377.470 4.280 ;
        RECT 378.310 0.155 379.770 4.280 ;
        RECT 380.610 0.155 382.070 4.280 ;
        RECT 382.910 0.155 384.370 4.280 ;
        RECT 385.210 0.155 386.670 4.280 ;
        RECT 387.510 0.155 388.970 4.280 ;
        RECT 389.810 0.155 391.270 4.280 ;
        RECT 392.110 0.155 393.570 4.280 ;
        RECT 394.410 0.155 395.870 4.280 ;
        RECT 396.710 0.155 398.170 4.280 ;
        RECT 399.010 0.155 400.470 4.280 ;
        RECT 401.310 0.155 402.770 4.280 ;
        RECT 403.610 0.155 405.070 4.280 ;
        RECT 405.910 0.155 407.370 4.280 ;
        RECT 408.210 0.155 409.670 4.280 ;
        RECT 410.510 0.155 411.970 4.280 ;
        RECT 412.810 0.155 414.270 4.280 ;
        RECT 415.110 0.155 416.570 4.280 ;
        RECT 417.410 0.155 418.870 4.280 ;
        RECT 419.710 0.155 421.170 4.280 ;
        RECT 422.010 0.155 423.470 4.280 ;
        RECT 424.310 0.155 425.770 4.280 ;
        RECT 426.610 0.155 428.070 4.280 ;
        RECT 428.910 0.155 430.370 4.280 ;
        RECT 431.210 0.155 432.670 4.280 ;
        RECT 433.510 0.155 434.970 4.280 ;
        RECT 435.810 0.155 437.270 4.280 ;
        RECT 438.110 0.155 439.570 4.280 ;
        RECT 440.410 0.155 441.870 4.280 ;
        RECT 442.710 0.155 444.170 4.280 ;
        RECT 445.010 0.155 446.470 4.280 ;
        RECT 447.310 0.155 448.770 4.280 ;
        RECT 449.610 0.155 451.070 4.280 ;
        RECT 451.910 0.155 453.370 4.280 ;
        RECT 454.210 0.155 455.670 4.280 ;
        RECT 456.510 0.155 457.970 4.280 ;
        RECT 458.810 0.155 460.270 4.280 ;
        RECT 461.110 0.155 462.570 4.280 ;
        RECT 463.410 0.155 464.870 4.280 ;
        RECT 465.710 0.155 467.170 4.280 ;
        RECT 468.010 0.155 469.470 4.280 ;
        RECT 470.310 0.155 471.770 4.280 ;
        RECT 472.610 0.155 474.070 4.280 ;
        RECT 474.910 0.155 476.370 4.280 ;
        RECT 477.210 0.155 478.670 4.280 ;
        RECT 479.510 0.155 480.970 4.280 ;
        RECT 481.810 0.155 483.270 4.280 ;
        RECT 484.110 0.155 485.570 4.280 ;
        RECT 486.410 0.155 487.870 4.280 ;
        RECT 488.710 0.155 490.170 4.280 ;
        RECT 491.010 0.155 492.470 4.280 ;
        RECT 493.310 0.155 494.770 4.280 ;
        RECT 495.610 0.155 497.070 4.280 ;
        RECT 497.910 0.155 499.370 4.280 ;
        RECT 500.210 0.155 501.670 4.280 ;
        RECT 502.510 0.155 503.970 4.280 ;
        RECT 504.810 0.155 506.270 4.280 ;
        RECT 507.110 0.155 508.570 4.280 ;
        RECT 509.410 0.155 510.870 4.280 ;
        RECT 511.710 0.155 513.170 4.280 ;
        RECT 514.010 0.155 515.470 4.280 ;
        RECT 516.310 0.155 517.770 4.280 ;
        RECT 518.610 0.155 520.070 4.280 ;
        RECT 520.910 0.155 522.370 4.280 ;
        RECT 523.210 0.155 524.670 4.280 ;
        RECT 525.510 0.155 526.970 4.280 ;
        RECT 527.810 0.155 529.270 4.280 ;
        RECT 530.110 0.155 531.570 4.280 ;
        RECT 532.410 0.155 533.870 4.280 ;
        RECT 534.710 0.155 536.170 4.280 ;
        RECT 537.010 0.155 538.470 4.280 ;
        RECT 539.310 0.155 540.770 4.280 ;
        RECT 541.610 0.155 543.070 4.280 ;
        RECT 543.910 0.155 545.370 4.280 ;
        RECT 546.210 0.155 547.670 4.280 ;
        RECT 548.510 0.155 549.970 4.280 ;
        RECT 550.810 0.155 552.270 4.280 ;
        RECT 553.110 0.155 554.570 4.280 ;
        RECT 555.410 0.155 556.870 4.280 ;
        RECT 557.710 0.155 559.170 4.280 ;
        RECT 560.010 0.155 561.470 4.280 ;
        RECT 562.310 0.155 563.770 4.280 ;
        RECT 564.610 0.155 566.070 4.280 ;
        RECT 566.910 0.155 568.370 4.280 ;
        RECT 569.210 0.155 570.670 4.280 ;
        RECT 571.510 0.155 572.970 4.280 ;
        RECT 573.810 0.155 575.270 4.280 ;
        RECT 576.110 0.155 577.570 4.280 ;
        RECT 578.410 0.155 579.870 4.280 ;
        RECT 580.710 0.155 582.170 4.280 ;
        RECT 583.010 0.155 584.470 4.280 ;
        RECT 585.310 0.155 586.770 4.280 ;
        RECT 587.610 0.155 589.070 4.280 ;
        RECT 589.910 0.155 591.370 4.280 ;
        RECT 592.210 0.155 593.670 4.280 ;
        RECT 594.510 0.155 595.970 4.280 ;
        RECT 596.810 0.155 598.270 4.280 ;
        RECT 599.110 0.155 600.570 4.280 ;
        RECT 601.410 0.155 602.870 4.280 ;
        RECT 603.710 0.155 605.170 4.280 ;
        RECT 606.010 0.155 607.470 4.280 ;
        RECT 608.310 0.155 609.770 4.280 ;
        RECT 610.610 0.155 612.070 4.280 ;
        RECT 612.910 0.155 614.370 4.280 ;
        RECT 615.210 0.155 616.670 4.280 ;
        RECT 617.510 0.155 618.970 4.280 ;
        RECT 619.810 0.155 621.270 4.280 ;
        RECT 622.110 0.155 623.570 4.280 ;
        RECT 624.410 0.155 625.870 4.280 ;
        RECT 626.710 0.155 628.170 4.280 ;
        RECT 629.010 0.155 630.470 4.280 ;
        RECT 631.310 0.155 632.770 4.280 ;
        RECT 633.610 0.155 635.070 4.280 ;
        RECT 635.910 0.155 637.370 4.280 ;
        RECT 638.210 0.155 639.670 4.280 ;
        RECT 640.510 0.155 641.970 4.280 ;
        RECT 642.810 0.155 644.270 4.280 ;
        RECT 645.110 0.155 646.570 4.280 ;
        RECT 647.410 0.155 648.870 4.280 ;
        RECT 649.710 0.155 651.170 4.280 ;
        RECT 652.010 0.155 653.470 4.280 ;
        RECT 654.310 0.155 655.770 4.280 ;
        RECT 656.610 0.155 658.070 4.280 ;
        RECT 658.910 0.155 660.370 4.280 ;
        RECT 661.210 0.155 662.670 4.280 ;
        RECT 663.510 0.155 664.970 4.280 ;
        RECT 665.810 0.155 667.270 4.280 ;
        RECT 668.110 0.155 669.570 4.280 ;
        RECT 670.410 0.155 671.870 4.280 ;
        RECT 672.710 0.155 674.170 4.280 ;
        RECT 675.010 0.155 676.470 4.280 ;
        RECT 677.310 0.155 678.770 4.280 ;
        RECT 679.610 0.155 681.070 4.280 ;
        RECT 681.910 0.155 683.370 4.280 ;
        RECT 684.210 0.155 685.670 4.280 ;
        RECT 686.510 0.155 687.970 4.280 ;
        RECT 688.810 0.155 690.270 4.280 ;
        RECT 691.110 0.155 692.570 4.280 ;
        RECT 693.410 0.155 694.870 4.280 ;
        RECT 695.710 0.155 697.170 4.280 ;
        RECT 698.010 0.155 699.470 4.280 ;
        RECT 700.310 0.155 701.770 4.280 ;
        RECT 702.610 0.155 704.070 4.280 ;
        RECT 704.910 0.155 706.370 4.280 ;
        RECT 707.210 0.155 708.670 4.280 ;
        RECT 709.510 0.155 710.970 4.280 ;
        RECT 711.810 0.155 713.270 4.280 ;
        RECT 714.110 0.155 715.570 4.280 ;
        RECT 716.410 0.155 717.870 4.280 ;
        RECT 718.710 0.155 720.170 4.280 ;
        RECT 721.010 0.155 722.470 4.280 ;
        RECT 723.310 0.155 724.770 4.280 ;
        RECT 725.610 0.155 727.070 4.280 ;
        RECT 727.910 0.155 729.370 4.280 ;
        RECT 730.210 0.155 731.670 4.280 ;
        RECT 732.510 0.155 733.970 4.280 ;
        RECT 734.810 0.155 736.270 4.280 ;
        RECT 737.110 0.155 796.620 4.280 ;
      LAYER met3 ;
        RECT 4.000 792.520 795.600 793.385 ;
        RECT 4.000 787.120 796.000 792.520 ;
        RECT 4.000 785.720 795.600 787.120 ;
        RECT 4.000 780.320 796.000 785.720 ;
        RECT 4.400 778.920 795.600 780.320 ;
        RECT 4.000 773.520 796.000 778.920 ;
        RECT 4.000 772.120 795.600 773.520 ;
        RECT 4.000 766.720 796.000 772.120 ;
        RECT 4.000 765.320 795.600 766.720 ;
        RECT 4.000 759.920 796.000 765.320 ;
        RECT 4.000 758.520 795.600 759.920 ;
        RECT 4.000 753.120 796.000 758.520 ;
        RECT 4.000 751.720 795.600 753.120 ;
        RECT 4.000 746.320 796.000 751.720 ;
        RECT 4.000 744.920 795.600 746.320 ;
        RECT 4.000 742.240 796.000 744.920 ;
        RECT 4.400 740.840 796.000 742.240 ;
        RECT 4.000 739.520 796.000 740.840 ;
        RECT 4.000 738.120 795.600 739.520 ;
        RECT 4.000 732.720 796.000 738.120 ;
        RECT 4.000 731.320 795.600 732.720 ;
        RECT 4.000 725.920 796.000 731.320 ;
        RECT 4.000 724.520 795.600 725.920 ;
        RECT 4.000 719.120 796.000 724.520 ;
        RECT 4.000 717.720 795.600 719.120 ;
        RECT 4.000 712.320 796.000 717.720 ;
        RECT 4.000 710.920 795.600 712.320 ;
        RECT 4.000 705.520 796.000 710.920 ;
        RECT 4.000 704.160 795.600 705.520 ;
        RECT 4.400 704.120 795.600 704.160 ;
        RECT 4.400 702.760 796.000 704.120 ;
        RECT 4.000 698.720 796.000 702.760 ;
        RECT 4.000 697.320 795.600 698.720 ;
        RECT 4.000 691.920 796.000 697.320 ;
        RECT 4.000 690.520 795.600 691.920 ;
        RECT 4.000 685.120 796.000 690.520 ;
        RECT 4.000 683.720 795.600 685.120 ;
        RECT 4.000 678.320 796.000 683.720 ;
        RECT 4.000 676.920 795.600 678.320 ;
        RECT 4.000 671.520 796.000 676.920 ;
        RECT 4.000 670.120 795.600 671.520 ;
        RECT 4.000 666.080 796.000 670.120 ;
        RECT 4.400 664.720 796.000 666.080 ;
        RECT 4.400 664.680 795.600 664.720 ;
        RECT 4.000 663.320 795.600 664.680 ;
        RECT 4.000 657.920 796.000 663.320 ;
        RECT 4.000 656.520 795.600 657.920 ;
        RECT 4.000 651.120 796.000 656.520 ;
        RECT 4.000 649.720 795.600 651.120 ;
        RECT 4.000 644.320 796.000 649.720 ;
        RECT 4.000 642.920 795.600 644.320 ;
        RECT 4.000 637.520 796.000 642.920 ;
        RECT 4.000 636.120 795.600 637.520 ;
        RECT 4.000 630.720 796.000 636.120 ;
        RECT 4.000 629.320 795.600 630.720 ;
        RECT 4.000 628.000 796.000 629.320 ;
        RECT 4.400 626.600 796.000 628.000 ;
        RECT 4.000 623.920 796.000 626.600 ;
        RECT 4.000 622.520 795.600 623.920 ;
        RECT 4.000 617.120 796.000 622.520 ;
        RECT 4.000 615.720 795.600 617.120 ;
        RECT 4.000 610.320 796.000 615.720 ;
        RECT 4.000 608.920 795.600 610.320 ;
        RECT 4.000 603.520 796.000 608.920 ;
        RECT 4.000 602.120 795.600 603.520 ;
        RECT 4.000 596.720 796.000 602.120 ;
        RECT 4.000 595.320 795.600 596.720 ;
        RECT 4.000 589.920 796.000 595.320 ;
        RECT 4.400 588.520 795.600 589.920 ;
        RECT 4.000 583.120 796.000 588.520 ;
        RECT 4.000 581.720 795.600 583.120 ;
        RECT 4.000 576.320 796.000 581.720 ;
        RECT 4.000 574.920 795.600 576.320 ;
        RECT 4.000 569.520 796.000 574.920 ;
        RECT 4.000 568.120 795.600 569.520 ;
        RECT 4.000 562.720 796.000 568.120 ;
        RECT 4.000 561.320 795.600 562.720 ;
        RECT 4.000 555.920 796.000 561.320 ;
        RECT 4.000 554.520 795.600 555.920 ;
        RECT 4.000 551.840 796.000 554.520 ;
        RECT 4.400 550.440 796.000 551.840 ;
        RECT 4.000 549.120 796.000 550.440 ;
        RECT 4.000 547.720 795.600 549.120 ;
        RECT 4.000 542.320 796.000 547.720 ;
        RECT 4.000 540.920 795.600 542.320 ;
        RECT 4.000 535.520 796.000 540.920 ;
        RECT 4.000 534.120 795.600 535.520 ;
        RECT 4.000 528.720 796.000 534.120 ;
        RECT 4.000 527.320 795.600 528.720 ;
        RECT 4.000 521.920 796.000 527.320 ;
        RECT 4.000 520.520 795.600 521.920 ;
        RECT 4.000 515.120 796.000 520.520 ;
        RECT 4.000 513.760 795.600 515.120 ;
        RECT 4.400 513.720 795.600 513.760 ;
        RECT 4.400 512.360 796.000 513.720 ;
        RECT 4.000 508.320 796.000 512.360 ;
        RECT 4.000 506.920 795.600 508.320 ;
        RECT 4.000 501.520 796.000 506.920 ;
        RECT 4.000 500.120 795.600 501.520 ;
        RECT 4.000 494.720 796.000 500.120 ;
        RECT 4.000 493.320 795.600 494.720 ;
        RECT 4.000 487.920 796.000 493.320 ;
        RECT 4.000 486.520 795.600 487.920 ;
        RECT 4.000 481.120 796.000 486.520 ;
        RECT 4.000 479.720 795.600 481.120 ;
        RECT 4.000 475.680 796.000 479.720 ;
        RECT 4.400 474.320 796.000 475.680 ;
        RECT 4.400 474.280 795.600 474.320 ;
        RECT 4.000 472.920 795.600 474.280 ;
        RECT 4.000 467.520 796.000 472.920 ;
        RECT 4.000 466.120 795.600 467.520 ;
        RECT 4.000 460.720 796.000 466.120 ;
        RECT 4.000 459.320 795.600 460.720 ;
        RECT 4.000 453.920 796.000 459.320 ;
        RECT 4.000 452.520 795.600 453.920 ;
        RECT 4.000 447.120 796.000 452.520 ;
        RECT 4.000 445.720 795.600 447.120 ;
        RECT 4.000 440.320 796.000 445.720 ;
        RECT 4.000 438.920 795.600 440.320 ;
        RECT 4.000 437.600 796.000 438.920 ;
        RECT 4.400 436.200 796.000 437.600 ;
        RECT 4.000 433.520 796.000 436.200 ;
        RECT 4.000 432.120 795.600 433.520 ;
        RECT 4.000 426.720 796.000 432.120 ;
        RECT 4.000 425.320 795.600 426.720 ;
        RECT 4.000 419.920 796.000 425.320 ;
        RECT 4.000 418.520 795.600 419.920 ;
        RECT 4.000 413.120 796.000 418.520 ;
        RECT 4.000 411.720 795.600 413.120 ;
        RECT 4.000 406.320 796.000 411.720 ;
        RECT 4.000 404.920 795.600 406.320 ;
        RECT 4.000 399.520 796.000 404.920 ;
        RECT 4.400 398.120 795.600 399.520 ;
        RECT 4.000 392.720 796.000 398.120 ;
        RECT 4.000 391.320 795.600 392.720 ;
        RECT 4.000 385.920 796.000 391.320 ;
        RECT 4.000 384.520 795.600 385.920 ;
        RECT 4.000 379.120 796.000 384.520 ;
        RECT 4.000 377.720 795.600 379.120 ;
        RECT 4.000 372.320 796.000 377.720 ;
        RECT 4.000 370.920 795.600 372.320 ;
        RECT 4.000 365.520 796.000 370.920 ;
        RECT 4.000 364.120 795.600 365.520 ;
        RECT 4.000 361.440 796.000 364.120 ;
        RECT 4.400 360.040 796.000 361.440 ;
        RECT 4.000 358.720 796.000 360.040 ;
        RECT 4.000 357.320 795.600 358.720 ;
        RECT 4.000 351.920 796.000 357.320 ;
        RECT 4.000 350.520 795.600 351.920 ;
        RECT 4.000 345.120 796.000 350.520 ;
        RECT 4.000 343.720 795.600 345.120 ;
        RECT 4.000 338.320 796.000 343.720 ;
        RECT 4.000 336.920 795.600 338.320 ;
        RECT 4.000 331.520 796.000 336.920 ;
        RECT 4.000 330.120 795.600 331.520 ;
        RECT 4.000 324.720 796.000 330.120 ;
        RECT 4.000 323.360 795.600 324.720 ;
        RECT 4.400 323.320 795.600 323.360 ;
        RECT 4.400 321.960 796.000 323.320 ;
        RECT 4.000 317.920 796.000 321.960 ;
        RECT 4.000 316.520 795.600 317.920 ;
        RECT 4.000 311.120 796.000 316.520 ;
        RECT 4.000 309.720 795.600 311.120 ;
        RECT 4.000 304.320 796.000 309.720 ;
        RECT 4.000 302.920 795.600 304.320 ;
        RECT 4.000 297.520 796.000 302.920 ;
        RECT 4.000 296.120 795.600 297.520 ;
        RECT 4.000 290.720 796.000 296.120 ;
        RECT 4.000 289.320 795.600 290.720 ;
        RECT 4.000 285.280 796.000 289.320 ;
        RECT 4.400 283.920 796.000 285.280 ;
        RECT 4.400 283.880 795.600 283.920 ;
        RECT 4.000 282.520 795.600 283.880 ;
        RECT 4.000 277.120 796.000 282.520 ;
        RECT 4.000 275.720 795.600 277.120 ;
        RECT 4.000 270.320 796.000 275.720 ;
        RECT 4.000 268.920 795.600 270.320 ;
        RECT 4.000 263.520 796.000 268.920 ;
        RECT 4.000 262.120 795.600 263.520 ;
        RECT 4.000 256.720 796.000 262.120 ;
        RECT 4.000 255.320 795.600 256.720 ;
        RECT 4.000 249.920 796.000 255.320 ;
        RECT 4.000 248.520 795.600 249.920 ;
        RECT 4.000 247.200 796.000 248.520 ;
        RECT 4.400 245.800 796.000 247.200 ;
        RECT 4.000 243.120 796.000 245.800 ;
        RECT 4.000 241.720 795.600 243.120 ;
        RECT 4.000 236.320 796.000 241.720 ;
        RECT 4.000 234.920 795.600 236.320 ;
        RECT 4.000 229.520 796.000 234.920 ;
        RECT 4.000 228.120 795.600 229.520 ;
        RECT 4.000 222.720 796.000 228.120 ;
        RECT 4.000 221.320 795.600 222.720 ;
        RECT 4.000 215.920 796.000 221.320 ;
        RECT 4.000 214.520 795.600 215.920 ;
        RECT 4.000 209.120 796.000 214.520 ;
        RECT 4.400 207.720 795.600 209.120 ;
        RECT 4.000 202.320 796.000 207.720 ;
        RECT 4.000 200.920 795.600 202.320 ;
        RECT 4.000 195.520 796.000 200.920 ;
        RECT 4.000 194.120 795.600 195.520 ;
        RECT 4.000 188.720 796.000 194.120 ;
        RECT 4.000 187.320 795.600 188.720 ;
        RECT 4.000 181.920 796.000 187.320 ;
        RECT 4.000 180.520 795.600 181.920 ;
        RECT 4.000 175.120 796.000 180.520 ;
        RECT 4.000 173.720 795.600 175.120 ;
        RECT 4.000 171.040 796.000 173.720 ;
        RECT 4.400 169.640 796.000 171.040 ;
        RECT 4.000 168.320 796.000 169.640 ;
        RECT 4.000 166.920 795.600 168.320 ;
        RECT 4.000 161.520 796.000 166.920 ;
        RECT 4.000 160.120 795.600 161.520 ;
        RECT 4.000 154.720 796.000 160.120 ;
        RECT 4.000 153.320 795.600 154.720 ;
        RECT 4.000 147.920 796.000 153.320 ;
        RECT 4.000 146.520 795.600 147.920 ;
        RECT 4.000 141.120 796.000 146.520 ;
        RECT 4.000 139.720 795.600 141.120 ;
        RECT 4.000 134.320 796.000 139.720 ;
        RECT 4.000 132.960 795.600 134.320 ;
        RECT 4.400 132.920 795.600 132.960 ;
        RECT 4.400 131.560 796.000 132.920 ;
        RECT 4.000 127.520 796.000 131.560 ;
        RECT 4.000 126.120 795.600 127.520 ;
        RECT 4.000 120.720 796.000 126.120 ;
        RECT 4.000 119.320 795.600 120.720 ;
        RECT 4.000 113.920 796.000 119.320 ;
        RECT 4.000 112.520 795.600 113.920 ;
        RECT 4.000 107.120 796.000 112.520 ;
        RECT 4.000 105.720 795.600 107.120 ;
        RECT 4.000 100.320 796.000 105.720 ;
        RECT 4.000 98.920 795.600 100.320 ;
        RECT 4.000 94.880 796.000 98.920 ;
        RECT 4.400 93.520 796.000 94.880 ;
        RECT 4.400 93.480 795.600 93.520 ;
        RECT 4.000 92.120 795.600 93.480 ;
        RECT 4.000 86.720 796.000 92.120 ;
        RECT 4.000 85.320 795.600 86.720 ;
        RECT 4.000 79.920 796.000 85.320 ;
        RECT 4.000 78.520 795.600 79.920 ;
        RECT 4.000 73.120 796.000 78.520 ;
        RECT 4.000 71.720 795.600 73.120 ;
        RECT 4.000 66.320 796.000 71.720 ;
        RECT 4.000 64.920 795.600 66.320 ;
        RECT 4.000 59.520 796.000 64.920 ;
        RECT 4.000 58.120 795.600 59.520 ;
        RECT 4.000 56.800 796.000 58.120 ;
        RECT 4.400 55.400 796.000 56.800 ;
        RECT 4.000 52.720 796.000 55.400 ;
        RECT 4.000 51.320 795.600 52.720 ;
        RECT 4.000 45.920 796.000 51.320 ;
        RECT 4.000 44.520 795.600 45.920 ;
        RECT 4.000 39.120 796.000 44.520 ;
        RECT 4.000 37.720 795.600 39.120 ;
        RECT 4.000 32.320 796.000 37.720 ;
        RECT 4.000 30.920 795.600 32.320 ;
        RECT 4.000 25.520 796.000 30.920 ;
        RECT 4.000 24.120 795.600 25.520 ;
        RECT 4.000 18.720 796.000 24.120 ;
        RECT 4.400 17.320 795.600 18.720 ;
        RECT 4.000 11.920 796.000 17.320 ;
        RECT 4.000 10.520 795.600 11.920 ;
        RECT 4.000 5.120 796.000 10.520 ;
        RECT 4.000 3.720 795.600 5.120 ;
        RECT 4.000 0.175 796.000 3.720 ;
      LAYER met4 ;
        RECT 177.855 10.240 251.040 785.225 ;
        RECT 253.440 10.240 327.840 785.225 ;
        RECT 330.240 10.240 404.640 785.225 ;
        RECT 407.040 10.240 481.440 785.225 ;
        RECT 483.840 10.240 558.240 785.225 ;
        RECT 560.640 10.240 635.040 785.225 ;
        RECT 637.440 10.240 711.840 785.225 ;
        RECT 714.240 10.240 779.865 785.225 ;
        RECT 177.855 0.855 779.865 10.240 ;
  END
END bary_pipe_m
END LIBRARY

