VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO busarb_2_2
  CLASS BLOCK ;
  FOREIGN busarb_2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 450.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 13.890 446.000 14.170 450.000 ;
    END
  END clk_i
  PIN mports_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 17.570 446.000 17.850 450.000 ;
    END
  END mports_i[0]
  PIN mports_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 201.570 446.000 201.850 450.000 ;
    END
  END mports_i[100]
  PIN mports_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 446.000 203.690 450.000 ;
    END
  END mports_i[101]
  PIN mports_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 205.250 446.000 205.530 450.000 ;
    END
  END mports_i[102]
  PIN mports_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 207.090 446.000 207.370 450.000 ;
    END
  END mports_i[103]
  PIN mports_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 208.930 446.000 209.210 450.000 ;
    END
  END mports_i[104]
  PIN mports_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 210.770 446.000 211.050 450.000 ;
    END
  END mports_i[105]
  PIN mports_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 446.000 212.890 450.000 ;
    END
  END mports_i[106]
  PIN mports_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 214.450 446.000 214.730 450.000 ;
    END
  END mports_i[107]
  PIN mports_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 216.290 446.000 216.570 450.000 ;
    END
  END mports_i[108]
  PIN mports_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 218.130 446.000 218.410 450.000 ;
    END
  END mports_i[109]
  PIN mports_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 35.970 446.000 36.250 450.000 ;
    END
  END mports_i[10]
  PIN mports_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 219.970 446.000 220.250 450.000 ;
    END
  END mports_i[110]
  PIN mports_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 221.810 446.000 222.090 450.000 ;
    END
  END mports_i[111]
  PIN mports_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 223.650 446.000 223.930 450.000 ;
    END
  END mports_i[112]
  PIN mports_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 446.000 225.770 450.000 ;
    END
  END mports_i[113]
  PIN mports_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 227.330 446.000 227.610 450.000 ;
    END
  END mports_i[114]
  PIN mports_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 229.170 446.000 229.450 450.000 ;
    END
  END mports_i[115]
  PIN mports_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 446.000 231.290 450.000 ;
    END
  END mports_i[116]
  PIN mports_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 232.850 446.000 233.130 450.000 ;
    END
  END mports_i[117]
  PIN mports_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 234.690 446.000 234.970 450.000 ;
    END
  END mports_i[118]
  PIN mports_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 236.530 446.000 236.810 450.000 ;
    END
  END mports_i[119]
  PIN mports_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 37.810 446.000 38.090 450.000 ;
    END
  END mports_i[11]
  PIN mports_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 238.370 446.000 238.650 450.000 ;
    END
  END mports_i[120]
  PIN mports_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 240.210 446.000 240.490 450.000 ;
    END
  END mports_i[121]
  PIN mports_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 242.050 446.000 242.330 450.000 ;
    END
  END mports_i[122]
  PIN mports_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 446.000 244.170 450.000 ;
    END
  END mports_i[123]
  PIN mports_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 245.730 446.000 246.010 450.000 ;
    END
  END mports_i[124]
  PIN mports_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 247.570 446.000 247.850 450.000 ;
    END
  END mports_i[125]
  PIN mports_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 249.410 446.000 249.690 450.000 ;
    END
  END mports_i[126]
  PIN mports_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 251.250 446.000 251.530 450.000 ;
    END
  END mports_i[127]
  PIN mports_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 253.090 446.000 253.370 450.000 ;
    END
  END mports_i[128]
  PIN mports_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 254.930 446.000 255.210 450.000 ;
    END
  END mports_i[129]
  PIN mports_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 39.650 446.000 39.930 450.000 ;
    END
  END mports_i[12]
  PIN mports_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 256.770 446.000 257.050 450.000 ;
    END
  END mports_i[130]
  PIN mports_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 258.610 446.000 258.890 450.000 ;
    END
  END mports_i[131]
  PIN mports_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 446.000 260.730 450.000 ;
    END
  END mports_i[132]
  PIN mports_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 262.290 446.000 262.570 450.000 ;
    END
  END mports_i[133]
  PIN mports_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 264.130 446.000 264.410 450.000 ;
    END
  END mports_i[134]
  PIN mports_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 265.970 446.000 266.250 450.000 ;
    END
  END mports_i[135]
  PIN mports_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 267.810 446.000 268.090 450.000 ;
    END
  END mports_i[136]
  PIN mports_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 446.000 269.930 450.000 ;
    END
  END mports_i[137]
  PIN mports_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 271.490 446.000 271.770 450.000 ;
    END
  END mports_i[138]
  PIN mports_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 273.330 446.000 273.610 450.000 ;
    END
  END mports_i[139]
  PIN mports_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 41.490 446.000 41.770 450.000 ;
    END
  END mports_i[13]
  PIN mports_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 275.170 446.000 275.450 450.000 ;
    END
  END mports_i[140]
  PIN mports_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 277.010 446.000 277.290 450.000 ;
    END
  END mports_i[141]
  PIN mports_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 278.850 446.000 279.130 450.000 ;
    END
  END mports_i[142]
  PIN mports_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 280.690 446.000 280.970 450.000 ;
    END
  END mports_i[143]
  PIN mports_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 282.530 446.000 282.810 450.000 ;
    END
  END mports_i[144]
  PIN mports_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 284.370 446.000 284.650 450.000 ;
    END
  END mports_i[145]
  PIN mports_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 286.210 446.000 286.490 450.000 ;
    END
  END mports_i[146]
  PIN mports_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 288.050 446.000 288.330 450.000 ;
    END
  END mports_i[147]
  PIN mports_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 446.000 290.170 450.000 ;
    END
  END mports_i[148]
  PIN mports_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 291.730 446.000 292.010 450.000 ;
    END
  END mports_i[149]
  PIN mports_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 43.330 446.000 43.610 450.000 ;
    END
  END mports_i[14]
  PIN mports_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 293.570 446.000 293.850 450.000 ;
    END
  END mports_i[150]
  PIN mports_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 295.410 446.000 295.690 450.000 ;
    END
  END mports_i[151]
  PIN mports_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 297.250 446.000 297.530 450.000 ;
    END
  END mports_i[152]
  PIN mports_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 299.090 446.000 299.370 450.000 ;
    END
  END mports_i[153]
  PIN mports_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 300.930 446.000 301.210 450.000 ;
    END
  END mports_i[154]
  PIN mports_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 446.000 303.050 450.000 ;
    END
  END mports_i[155]
  PIN mports_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 304.610 446.000 304.890 450.000 ;
    END
  END mports_i[156]
  PIN mports_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 306.450 446.000 306.730 450.000 ;
    END
  END mports_i[157]
  PIN mports_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 308.290 446.000 308.570 450.000 ;
    END
  END mports_i[158]
  PIN mports_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 310.130 446.000 310.410 450.000 ;
    END
  END mports_i[159]
  PIN mports_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 446.000 45.450 450.000 ;
    END
  END mports_i[15]
  PIN mports_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 311.970 446.000 312.250 450.000 ;
    END
  END mports_i[160]
  PIN mports_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 313.810 446.000 314.090 450.000 ;
    END
  END mports_i[161]
  PIN mports_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 315.650 446.000 315.930 450.000 ;
    END
  END mports_i[162]
  PIN mports_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 317.490 446.000 317.770 450.000 ;
    END
  END mports_i[163]
  PIN mports_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 319.330 446.000 319.610 450.000 ;
    END
  END mports_i[164]
  PIN mports_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 321.170 446.000 321.450 450.000 ;
    END
  END mports_i[165]
  PIN mports_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 323.010 446.000 323.290 450.000 ;
    END
  END mports_i[166]
  PIN mports_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 324.850 446.000 325.130 450.000 ;
    END
  END mports_i[167]
  PIN mports_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 326.690 446.000 326.970 450.000 ;
    END
  END mports_i[168]
  PIN mports_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 328.530 446.000 328.810 450.000 ;
    END
  END mports_i[169]
  PIN mports_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 446.000 47.290 450.000 ;
    END
  END mports_i[16]
  PIN mports_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 330.370 446.000 330.650 450.000 ;
    END
  END mports_i[170]
  PIN mports_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 332.210 446.000 332.490 450.000 ;
    END
  END mports_i[171]
  PIN mports_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 334.050 446.000 334.330 450.000 ;
    END
  END mports_i[172]
  PIN mports_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 335.890 446.000 336.170 450.000 ;
    END
  END mports_i[173]
  PIN mports_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 337.730 446.000 338.010 450.000 ;
    END
  END mports_i[174]
  PIN mports_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 339.570 446.000 339.850 450.000 ;
    END
  END mports_i[175]
  PIN mports_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 446.000 341.690 450.000 ;
    END
  END mports_i[176]
  PIN mports_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 343.250 446.000 343.530 450.000 ;
    END
  END mports_i[177]
  PIN mports_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 345.090 446.000 345.370 450.000 ;
    END
  END mports_i[178]
  PIN mports_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 346.930 446.000 347.210 450.000 ;
    END
  END mports_i[179]
  PIN mports_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 446.000 49.130 450.000 ;
    END
  END mports_i[17]
  PIN mports_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 348.770 446.000 349.050 450.000 ;
    END
  END mports_i[180]
  PIN mports_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 350.610 446.000 350.890 450.000 ;
    END
  END mports_i[181]
  PIN mports_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 446.000 352.730 450.000 ;
    END
  END mports_i[182]
  PIN mports_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 354.290 446.000 354.570 450.000 ;
    END
  END mports_i[183]
  PIN mports_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 356.130 446.000 356.410 450.000 ;
    END
  END mports_i[184]
  PIN mports_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 357.970 446.000 358.250 450.000 ;
    END
  END mports_i[185]
  PIN mports_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 359.810 446.000 360.090 450.000 ;
    END
  END mports_i[186]
  PIN mports_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 446.000 361.930 450.000 ;
    END
  END mports_i[187]
  PIN mports_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 363.490 446.000 363.770 450.000 ;
    END
  END mports_i[188]
  PIN mports_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 446.000 365.610 450.000 ;
    END
  END mports_i[189]
  PIN mports_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 50.690 446.000 50.970 450.000 ;
    END
  END mports_i[18]
  PIN mports_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 367.170 446.000 367.450 450.000 ;
    END
  END mports_i[190]
  PIN mports_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 369.010 446.000 369.290 450.000 ;
    END
  END mports_i[191]
  PIN mports_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 370.850 446.000 371.130 450.000 ;
    END
  END mports_i[192]
  PIN mports_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 372.690 446.000 372.970 450.000 ;
    END
  END mports_i[193]
  PIN mports_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 374.530 446.000 374.810 450.000 ;
    END
  END mports_i[194]
  PIN mports_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 376.370 446.000 376.650 450.000 ;
    END
  END mports_i[195]
  PIN mports_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 378.210 446.000 378.490 450.000 ;
    END
  END mports_i[196]
  PIN mports_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 446.000 380.330 450.000 ;
    END
  END mports_i[197]
  PIN mports_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 381.890 446.000 382.170 450.000 ;
    END
  END mports_i[198]
  PIN mports_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 383.730 446.000 384.010 450.000 ;
    END
  END mports_i[199]
  PIN mports_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 52.530 446.000 52.810 450.000 ;
    END
  END mports_i[19]
  PIN mports_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 446.000 19.690 450.000 ;
    END
  END mports_i[1]
  PIN mports_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 385.570 446.000 385.850 450.000 ;
    END
  END mports_i[200]
  PIN mports_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 387.410 446.000 387.690 450.000 ;
    END
  END mports_i[201]
  PIN mports_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 389.250 446.000 389.530 450.000 ;
    END
  END mports_i[202]
  PIN mports_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 391.090 446.000 391.370 450.000 ;
    END
  END mports_i[203]
  PIN mports_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 446.000 393.210 450.000 ;
    END
  END mports_i[204]
  PIN mports_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 394.770 446.000 395.050 450.000 ;
    END
  END mports_i[205]
  PIN mports_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 396.610 446.000 396.890 450.000 ;
    END
  END mports_i[206]
  PIN mports_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 398.450 446.000 398.730 450.000 ;
    END
  END mports_i[207]
  PIN mports_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 400.290 446.000 400.570 450.000 ;
    END
  END mports_i[208]
  PIN mports_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 402.130 446.000 402.410 450.000 ;
    END
  END mports_i[209]
  PIN mports_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 54.370 446.000 54.650 450.000 ;
    END
  END mports_i[20]
  PIN mports_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 403.970 446.000 404.250 450.000 ;
    END
  END mports_i[210]
  PIN mports_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 405.810 446.000 406.090 450.000 ;
    END
  END mports_i[211]
  PIN mports_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 407.650 446.000 407.930 450.000 ;
    END
  END mports_i[212]
  PIN mports_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 446.000 409.770 450.000 ;
    END
  END mports_i[213]
  PIN mports_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 411.330 446.000 411.610 450.000 ;
    END
  END mports_i[214]
  PIN mports_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 413.170 446.000 413.450 450.000 ;
    END
  END mports_i[215]
  PIN mports_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 415.010 446.000 415.290 450.000 ;
    END
  END mports_i[216]
  PIN mports_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 416.850 446.000 417.130 450.000 ;
    END
  END mports_i[217]
  PIN mports_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 418.690 446.000 418.970 450.000 ;
    END
  END mports_i[218]
  PIN mports_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 420.530 446.000 420.810 450.000 ;
    END
  END mports_i[219]
  PIN mports_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 56.210 446.000 56.490 450.000 ;
    END
  END mports_i[21]
  PIN mports_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 422.370 446.000 422.650 450.000 ;
    END
  END mports_i[220]
  PIN mports_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 424.210 446.000 424.490 450.000 ;
    END
  END mports_i[221]
  PIN mports_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 426.050 446.000 426.330 450.000 ;
    END
  END mports_i[222]
  PIN mports_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 427.890 446.000 428.170 450.000 ;
    END
  END mports_i[223]
  PIN mports_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 429.730 446.000 430.010 450.000 ;
    END
  END mports_i[224]
  PIN mports_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 431.570 446.000 431.850 450.000 ;
    END
  END mports_i[225]
  PIN mports_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 433.410 446.000 433.690 450.000 ;
    END
  END mports_i[226]
  PIN mports_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 435.250 446.000 435.530 450.000 ;
    END
  END mports_i[227]
  PIN mports_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 446.000 58.330 450.000 ;
    END
  END mports_i[22]
  PIN mports_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 59.890 446.000 60.170 450.000 ;
    END
  END mports_i[23]
  PIN mports_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 61.730 446.000 62.010 450.000 ;
    END
  END mports_i[24]
  PIN mports_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 63.570 446.000 63.850 450.000 ;
    END
  END mports_i[25]
  PIN mports_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 65.410 446.000 65.690 450.000 ;
    END
  END mports_i[26]
  PIN mports_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 446.000 67.530 450.000 ;
    END
  END mports_i[27]
  PIN mports_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 69.090 446.000 69.370 450.000 ;
    END
  END mports_i[28]
  PIN mports_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 446.000 71.210 450.000 ;
    END
  END mports_i[29]
  PIN mports_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 21.250 446.000 21.530 450.000 ;
    END
  END mports_i[2]
  PIN mports_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 72.770 446.000 73.050 450.000 ;
    END
  END mports_i[30]
  PIN mports_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 446.000 74.890 450.000 ;
    END
  END mports_i[31]
  PIN mports_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 76.450 446.000 76.730 450.000 ;
    END
  END mports_i[32]
  PIN mports_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 446.000 78.570 450.000 ;
    END
  END mports_i[33]
  PIN mports_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 80.130 446.000 80.410 450.000 ;
    END
  END mports_i[34]
  PIN mports_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 81.970 446.000 82.250 450.000 ;
    END
  END mports_i[35]
  PIN mports_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 446.000 84.090 450.000 ;
    END
  END mports_i[36]
  PIN mports_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 85.650 446.000 85.930 450.000 ;
    END
  END mports_i[37]
  PIN mports_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 446.000 87.770 450.000 ;
    END
  END mports_i[38]
  PIN mports_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 89.330 446.000 89.610 450.000 ;
    END
  END mports_i[39]
  PIN mports_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 446.000 23.370 450.000 ;
    END
  END mports_i[3]
  PIN mports_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 91.170 446.000 91.450 450.000 ;
    END
  END mports_i[40]
  PIN mports_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 93.010 446.000 93.290 450.000 ;
    END
  END mports_i[41]
  PIN mports_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 446.000 95.130 450.000 ;
    END
  END mports_i[42]
  PIN mports_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 446.000 96.970 450.000 ;
    END
  END mports_i[43]
  PIN mports_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 446.000 98.810 450.000 ;
    END
  END mports_i[44]
  PIN mports_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 100.370 446.000 100.650 450.000 ;
    END
  END mports_i[45]
  PIN mports_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 102.210 446.000 102.490 450.000 ;
    END
  END mports_i[46]
  PIN mports_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 104.050 446.000 104.330 450.000 ;
    END
  END mports_i[47]
  PIN mports_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 105.890 446.000 106.170 450.000 ;
    END
  END mports_i[48]
  PIN mports_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 446.000 108.010 450.000 ;
    END
  END mports_i[49]
  PIN mports_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 24.930 446.000 25.210 450.000 ;
    END
  END mports_i[4]
  PIN mports_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 446.000 109.850 450.000 ;
    END
  END mports_i[50]
  PIN mports_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 111.410 446.000 111.690 450.000 ;
    END
  END mports_i[51]
  PIN mports_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 113.250 446.000 113.530 450.000 ;
    END
  END mports_i[52]
  PIN mports_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 446.000 115.370 450.000 ;
    END
  END mports_i[53]
  PIN mports_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 116.930 446.000 117.210 450.000 ;
    END
  END mports_i[54]
  PIN mports_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 118.770 446.000 119.050 450.000 ;
    END
  END mports_i[55]
  PIN mports_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 120.610 446.000 120.890 450.000 ;
    END
  END mports_i[56]
  PIN mports_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 446.000 122.730 450.000 ;
    END
  END mports_i[57]
  PIN mports_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 124.290 446.000 124.570 450.000 ;
    END
  END mports_i[58]
  PIN mports_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 446.000 126.410 450.000 ;
    END
  END mports_i[59]
  PIN mports_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 26.770 446.000 27.050 450.000 ;
    END
  END mports_i[5]
  PIN mports_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 127.970 446.000 128.250 450.000 ;
    END
  END mports_i[60]
  PIN mports_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 446.000 130.090 450.000 ;
    END
  END mports_i[61]
  PIN mports_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 131.650 446.000 131.930 450.000 ;
    END
  END mports_i[62]
  PIN mports_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 133.490 446.000 133.770 450.000 ;
    END
  END mports_i[63]
  PIN mports_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 446.000 135.610 450.000 ;
    END
  END mports_i[64]
  PIN mports_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 446.000 137.450 450.000 ;
    END
  END mports_i[65]
  PIN mports_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 139.010 446.000 139.290 450.000 ;
    END
  END mports_i[66]
  PIN mports_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 140.850 446.000 141.130 450.000 ;
    END
  END mports_i[67]
  PIN mports_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 142.690 446.000 142.970 450.000 ;
    END
  END mports_i[68]
  PIN mports_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 446.000 144.810 450.000 ;
    END
  END mports_i[69]
  PIN mports_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 28.610 446.000 28.890 450.000 ;
    END
  END mports_i[6]
  PIN mports_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 146.370 446.000 146.650 450.000 ;
    END
  END mports_i[70]
  PIN mports_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 446.000 148.490 450.000 ;
    END
  END mports_i[71]
  PIN mports_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 150.050 446.000 150.330 450.000 ;
    END
  END mports_i[72]
  PIN mports_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 151.890 446.000 152.170 450.000 ;
    END
  END mports_i[73]
  PIN mports_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 153.730 446.000 154.010 450.000 ;
    END
  END mports_i[74]
  PIN mports_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 446.000 155.850 450.000 ;
    END
  END mports_i[75]
  PIN mports_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 157.410 446.000 157.690 450.000 ;
    END
  END mports_i[76]
  PIN mports_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 446.000 159.530 450.000 ;
    END
  END mports_i[77]
  PIN mports_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 446.000 161.370 450.000 ;
    END
  END mports_i[78]
  PIN mports_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 162.930 446.000 163.210 450.000 ;
    END
  END mports_i[79]
  PIN mports_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 446.000 30.730 450.000 ;
    END
  END mports_i[7]
  PIN mports_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 164.770 446.000 165.050 450.000 ;
    END
  END mports_i[80]
  PIN mports_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 166.610 446.000 166.890 450.000 ;
    END
  END mports_i[81]
  PIN mports_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 446.000 168.730 450.000 ;
    END
  END mports_i[82]
  PIN mports_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 446.000 170.570 450.000 ;
    END
  END mports_i[83]
  PIN mports_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 172.130 446.000 172.410 450.000 ;
    END
  END mports_i[84]
  PIN mports_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 446.000 174.250 450.000 ;
    END
  END mports_i[85]
  PIN mports_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 175.810 446.000 176.090 450.000 ;
    END
  END mports_i[86]
  PIN mports_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 177.650 446.000 177.930 450.000 ;
    END
  END mports_i[87]
  PIN mports_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 179.490 446.000 179.770 450.000 ;
    END
  END mports_i[88]
  PIN mports_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 181.330 446.000 181.610 450.000 ;
    END
  END mports_i[89]
  PIN mports_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 446.000 32.570 450.000 ;
    END
  END mports_i[8]
  PIN mports_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 183.170 446.000 183.450 450.000 ;
    END
  END mports_i[90]
  PIN mports_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 185.010 446.000 185.290 450.000 ;
    END
  END mports_i[91]
  PIN mports_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 446.000 187.130 450.000 ;
    END
  END mports_i[92]
  PIN mports_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 188.690 446.000 188.970 450.000 ;
    END
  END mports_i[93]
  PIN mports_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 446.000 190.810 450.000 ;
    END
  END mports_i[94]
  PIN mports_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 192.370 446.000 192.650 450.000 ;
    END
  END mports_i[95]
  PIN mports_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 446.000 194.490 450.000 ;
    END
  END mports_i[96]
  PIN mports_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 446.000 196.330 450.000 ;
    END
  END mports_i[97]
  PIN mports_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 197.890 446.000 198.170 450.000 ;
    END
  END mports_i[98]
  PIN mports_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 446.000 200.010 450.000 ;
    END
  END mports_i[99]
  PIN mports_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 34.130 446.000 34.410 450.000 ;
    END
  END mports_i[9]
  PIN mports_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END mports_o[0]
  PIN mports_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END mports_o[100]
  PIN mports_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END mports_o[101]
  PIN mports_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END mports_o[102]
  PIN mports_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END mports_o[103]
  PIN mports_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END mports_o[104]
  PIN mports_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END mports_o[105]
  PIN mports_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END mports_o[106]
  PIN mports_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END mports_o[107]
  PIN mports_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END mports_o[108]
  PIN mports_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END mports_o[109]
  PIN mports_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END mports_o[10]
  PIN mports_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END mports_o[110]
  PIN mports_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END mports_o[111]
  PIN mports_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END mports_o[112]
  PIN mports_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END mports_o[113]
  PIN mports_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END mports_o[114]
  PIN mports_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END mports_o[115]
  PIN mports_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END mports_o[116]
  PIN mports_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END mports_o[117]
  PIN mports_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END mports_o[118]
  PIN mports_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END mports_o[119]
  PIN mports_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END mports_o[11]
  PIN mports_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END mports_o[120]
  PIN mports_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END mports_o[121]
  PIN mports_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END mports_o[122]
  PIN mports_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END mports_o[123]
  PIN mports_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END mports_o[124]
  PIN mports_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END mports_o[125]
  PIN mports_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END mports_o[126]
  PIN mports_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END mports_o[127]
  PIN mports_o[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END mports_o[128]
  PIN mports_o[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END mports_o[129]
  PIN mports_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END mports_o[12]
  PIN mports_o[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END mports_o[130]
  PIN mports_o[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END mports_o[131]
  PIN mports_o[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END mports_o[132]
  PIN mports_o[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END mports_o[133]
  PIN mports_o[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END mports_o[134]
  PIN mports_o[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END mports_o[135]
  PIN mports_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END mports_o[13]
  PIN mports_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END mports_o[14]
  PIN mports_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END mports_o[15]
  PIN mports_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END mports_o[16]
  PIN mports_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END mports_o[17]
  PIN mports_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END mports_o[18]
  PIN mports_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END mports_o[19]
  PIN mports_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END mports_o[1]
  PIN mports_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END mports_o[20]
  PIN mports_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END mports_o[21]
  PIN mports_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END mports_o[22]
  PIN mports_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END mports_o[23]
  PIN mports_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END mports_o[24]
  PIN mports_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END mports_o[25]
  PIN mports_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END mports_o[26]
  PIN mports_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END mports_o[27]
  PIN mports_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END mports_o[28]
  PIN mports_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END mports_o[29]
  PIN mports_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END mports_o[2]
  PIN mports_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END mports_o[30]
  PIN mports_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END mports_o[31]
  PIN mports_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END mports_o[32]
  PIN mports_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END mports_o[33]
  PIN mports_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END mports_o[34]
  PIN mports_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END mports_o[35]
  PIN mports_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END mports_o[36]
  PIN mports_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END mports_o[37]
  PIN mports_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END mports_o[38]
  PIN mports_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END mports_o[39]
  PIN mports_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END mports_o[3]
  PIN mports_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END mports_o[40]
  PIN mports_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END mports_o[41]
  PIN mports_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END mports_o[42]
  PIN mports_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END mports_o[43]
  PIN mports_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END mports_o[44]
  PIN mports_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END mports_o[45]
  PIN mports_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END mports_o[46]
  PIN mports_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END mports_o[47]
  PIN mports_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END mports_o[48]
  PIN mports_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END mports_o[49]
  PIN mports_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END mports_o[4]
  PIN mports_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END mports_o[50]
  PIN mports_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END mports_o[51]
  PIN mports_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END mports_o[52]
  PIN mports_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END mports_o[53]
  PIN mports_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END mports_o[54]
  PIN mports_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END mports_o[55]
  PIN mports_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END mports_o[56]
  PIN mports_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END mports_o[57]
  PIN mports_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END mports_o[58]
  PIN mports_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END mports_o[59]
  PIN mports_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END mports_o[5]
  PIN mports_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END mports_o[60]
  PIN mports_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END mports_o[61]
  PIN mports_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END mports_o[62]
  PIN mports_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END mports_o[63]
  PIN mports_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END mports_o[64]
  PIN mports_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END mports_o[65]
  PIN mports_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END mports_o[66]
  PIN mports_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END mports_o[67]
  PIN mports_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END mports_o[68]
  PIN mports_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END mports_o[69]
  PIN mports_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END mports_o[6]
  PIN mports_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END mports_o[70]
  PIN mports_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END mports_o[71]
  PIN mports_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END mports_o[72]
  PIN mports_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END mports_o[73]
  PIN mports_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END mports_o[74]
  PIN mports_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END mports_o[75]
  PIN mports_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END mports_o[76]
  PIN mports_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END mports_o[77]
  PIN mports_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END mports_o[78]
  PIN mports_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END mports_o[79]
  PIN mports_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END mports_o[7]
  PIN mports_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END mports_o[80]
  PIN mports_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END mports_o[81]
  PIN mports_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END mports_o[82]
  PIN mports_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END mports_o[83]
  PIN mports_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END mports_o[84]
  PIN mports_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END mports_o[85]
  PIN mports_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END mports_o[86]
  PIN mports_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END mports_o[87]
  PIN mports_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END mports_o[88]
  PIN mports_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END mports_o[89]
  PIN mports_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END mports_o[8]
  PIN mports_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END mports_o[90]
  PIN mports_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END mports_o[91]
  PIN mports_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END mports_o[92]
  PIN mports_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END mports_o[93]
  PIN mports_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END mports_o[94]
  PIN mports_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END mports_o[95]
  PIN mports_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END mports_o[96]
  PIN mports_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END mports_o[97]
  PIN mports_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END mports_o[98]
  PIN mports_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END mports_o[99]
  PIN mports_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END mports_o[9]
  PIN nrst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 15.730 446.000 16.010 450.000 ;
    END
  END nrst_i
  PIN sports_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 40.840 450.000 41.440 ;
    END
  END sports_i[0]
  PIN sports_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 312.840 450.000 313.440 ;
    END
  END sports_i[100]
  PIN sports_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 315.560 450.000 316.160 ;
    END
  END sports_i[101]
  PIN sports_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 318.280 450.000 318.880 ;
    END
  END sports_i[102]
  PIN sports_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 321.000 450.000 321.600 ;
    END
  END sports_i[103]
  PIN sports_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 323.720 450.000 324.320 ;
    END
  END sports_i[104]
  PIN sports_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 326.440 450.000 327.040 ;
    END
  END sports_i[105]
  PIN sports_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 329.160 450.000 329.760 ;
    END
  END sports_i[106]
  PIN sports_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 331.880 450.000 332.480 ;
    END
  END sports_i[107]
  PIN sports_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 334.600 450.000 335.200 ;
    END
  END sports_i[108]
  PIN sports_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 337.320 450.000 337.920 ;
    END
  END sports_i[109]
  PIN sports_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 68.040 450.000 68.640 ;
    END
  END sports_i[10]
  PIN sports_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 340.040 450.000 340.640 ;
    END
  END sports_i[110]
  PIN sports_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 342.760 450.000 343.360 ;
    END
  END sports_i[111]
  PIN sports_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 345.480 450.000 346.080 ;
    END
  END sports_i[112]
  PIN sports_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 348.200 450.000 348.800 ;
    END
  END sports_i[113]
  PIN sports_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 350.920 450.000 351.520 ;
    END
  END sports_i[114]
  PIN sports_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 353.640 450.000 354.240 ;
    END
  END sports_i[115]
  PIN sports_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 356.360 450.000 356.960 ;
    END
  END sports_i[116]
  PIN sports_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 359.080 450.000 359.680 ;
    END
  END sports_i[117]
  PIN sports_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 361.800 450.000 362.400 ;
    END
  END sports_i[118]
  PIN sports_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 364.520 450.000 365.120 ;
    END
  END sports_i[119]
  PIN sports_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 70.760 450.000 71.360 ;
    END
  END sports_i[11]
  PIN sports_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 367.240 450.000 367.840 ;
    END
  END sports_i[120]
  PIN sports_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 369.960 450.000 370.560 ;
    END
  END sports_i[121]
  PIN sports_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 372.680 450.000 373.280 ;
    END
  END sports_i[122]
  PIN sports_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 375.400 450.000 376.000 ;
    END
  END sports_i[123]
  PIN sports_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 378.120 450.000 378.720 ;
    END
  END sports_i[124]
  PIN sports_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 380.840 450.000 381.440 ;
    END
  END sports_i[125]
  PIN sports_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 383.560 450.000 384.160 ;
    END
  END sports_i[126]
  PIN sports_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 386.280 450.000 386.880 ;
    END
  END sports_i[127]
  PIN sports_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 389.000 450.000 389.600 ;
    END
  END sports_i[128]
  PIN sports_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 391.720 450.000 392.320 ;
    END
  END sports_i[129]
  PIN sports_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 73.480 450.000 74.080 ;
    END
  END sports_i[12]
  PIN sports_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 394.440 450.000 395.040 ;
    END
  END sports_i[130]
  PIN sports_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 397.160 450.000 397.760 ;
    END
  END sports_i[131]
  PIN sports_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 399.880 450.000 400.480 ;
    END
  END sports_i[132]
  PIN sports_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 402.600 450.000 403.200 ;
    END
  END sports_i[133]
  PIN sports_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 405.320 450.000 405.920 ;
    END
  END sports_i[134]
  PIN sports_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 408.040 450.000 408.640 ;
    END
  END sports_i[135]
  PIN sports_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 76.200 450.000 76.800 ;
    END
  END sports_i[13]
  PIN sports_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 78.920 450.000 79.520 ;
    END
  END sports_i[14]
  PIN sports_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 81.640 450.000 82.240 ;
    END
  END sports_i[15]
  PIN sports_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 84.360 450.000 84.960 ;
    END
  END sports_i[16]
  PIN sports_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 87.080 450.000 87.680 ;
    END
  END sports_i[17]
  PIN sports_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 89.800 450.000 90.400 ;
    END
  END sports_i[18]
  PIN sports_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 92.520 450.000 93.120 ;
    END
  END sports_i[19]
  PIN sports_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 43.560 450.000 44.160 ;
    END
  END sports_i[1]
  PIN sports_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 95.240 450.000 95.840 ;
    END
  END sports_i[20]
  PIN sports_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 97.960 450.000 98.560 ;
    END
  END sports_i[21]
  PIN sports_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 100.680 450.000 101.280 ;
    END
  END sports_i[22]
  PIN sports_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 103.400 450.000 104.000 ;
    END
  END sports_i[23]
  PIN sports_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 106.120 450.000 106.720 ;
    END
  END sports_i[24]
  PIN sports_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 108.840 450.000 109.440 ;
    END
  END sports_i[25]
  PIN sports_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 111.560 450.000 112.160 ;
    END
  END sports_i[26]
  PIN sports_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 114.280 450.000 114.880 ;
    END
  END sports_i[27]
  PIN sports_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 117.000 450.000 117.600 ;
    END
  END sports_i[28]
  PIN sports_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 119.720 450.000 120.320 ;
    END
  END sports_i[29]
  PIN sports_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 46.280 450.000 46.880 ;
    END
  END sports_i[2]
  PIN sports_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 122.440 450.000 123.040 ;
    END
  END sports_i[30]
  PIN sports_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 125.160 450.000 125.760 ;
    END
  END sports_i[31]
  PIN sports_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 127.880 450.000 128.480 ;
    END
  END sports_i[32]
  PIN sports_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 130.600 450.000 131.200 ;
    END
  END sports_i[33]
  PIN sports_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 133.320 450.000 133.920 ;
    END
  END sports_i[34]
  PIN sports_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 136.040 450.000 136.640 ;
    END
  END sports_i[35]
  PIN sports_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 138.760 450.000 139.360 ;
    END
  END sports_i[36]
  PIN sports_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 141.480 450.000 142.080 ;
    END
  END sports_i[37]
  PIN sports_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 144.200 450.000 144.800 ;
    END
  END sports_i[38]
  PIN sports_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 146.920 450.000 147.520 ;
    END
  END sports_i[39]
  PIN sports_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 49.000 450.000 49.600 ;
    END
  END sports_i[3]
  PIN sports_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 149.640 450.000 150.240 ;
    END
  END sports_i[40]
  PIN sports_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 152.360 450.000 152.960 ;
    END
  END sports_i[41]
  PIN sports_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 155.080 450.000 155.680 ;
    END
  END sports_i[42]
  PIN sports_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 157.800 450.000 158.400 ;
    END
  END sports_i[43]
  PIN sports_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 160.520 450.000 161.120 ;
    END
  END sports_i[44]
  PIN sports_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 163.240 450.000 163.840 ;
    END
  END sports_i[45]
  PIN sports_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 165.960 450.000 166.560 ;
    END
  END sports_i[46]
  PIN sports_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 168.680 450.000 169.280 ;
    END
  END sports_i[47]
  PIN sports_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 171.400 450.000 172.000 ;
    END
  END sports_i[48]
  PIN sports_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 174.120 450.000 174.720 ;
    END
  END sports_i[49]
  PIN sports_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 51.720 450.000 52.320 ;
    END
  END sports_i[4]
  PIN sports_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 176.840 450.000 177.440 ;
    END
  END sports_i[50]
  PIN sports_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 179.560 450.000 180.160 ;
    END
  END sports_i[51]
  PIN sports_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 182.280 450.000 182.880 ;
    END
  END sports_i[52]
  PIN sports_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 185.000 450.000 185.600 ;
    END
  END sports_i[53]
  PIN sports_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 187.720 450.000 188.320 ;
    END
  END sports_i[54]
  PIN sports_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 190.440 450.000 191.040 ;
    END
  END sports_i[55]
  PIN sports_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 193.160 450.000 193.760 ;
    END
  END sports_i[56]
  PIN sports_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 195.880 450.000 196.480 ;
    END
  END sports_i[57]
  PIN sports_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 198.600 450.000 199.200 ;
    END
  END sports_i[58]
  PIN sports_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 201.320 450.000 201.920 ;
    END
  END sports_i[59]
  PIN sports_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 54.440 450.000 55.040 ;
    END
  END sports_i[5]
  PIN sports_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 204.040 450.000 204.640 ;
    END
  END sports_i[60]
  PIN sports_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 206.760 450.000 207.360 ;
    END
  END sports_i[61]
  PIN sports_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 209.480 450.000 210.080 ;
    END
  END sports_i[62]
  PIN sports_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 212.200 450.000 212.800 ;
    END
  END sports_i[63]
  PIN sports_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 214.920 450.000 215.520 ;
    END
  END sports_i[64]
  PIN sports_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 217.640 450.000 218.240 ;
    END
  END sports_i[65]
  PIN sports_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 220.360 450.000 220.960 ;
    END
  END sports_i[66]
  PIN sports_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 223.080 450.000 223.680 ;
    END
  END sports_i[67]
  PIN sports_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 225.800 450.000 226.400 ;
    END
  END sports_i[68]
  PIN sports_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 228.520 450.000 229.120 ;
    END
  END sports_i[69]
  PIN sports_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 57.160 450.000 57.760 ;
    END
  END sports_i[6]
  PIN sports_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 231.240 450.000 231.840 ;
    END
  END sports_i[70]
  PIN sports_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 233.960 450.000 234.560 ;
    END
  END sports_i[71]
  PIN sports_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 236.680 450.000 237.280 ;
    END
  END sports_i[72]
  PIN sports_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 239.400 450.000 240.000 ;
    END
  END sports_i[73]
  PIN sports_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 242.120 450.000 242.720 ;
    END
  END sports_i[74]
  PIN sports_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 244.840 450.000 245.440 ;
    END
  END sports_i[75]
  PIN sports_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 247.560 450.000 248.160 ;
    END
  END sports_i[76]
  PIN sports_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 250.280 450.000 250.880 ;
    END
  END sports_i[77]
  PIN sports_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 253.000 450.000 253.600 ;
    END
  END sports_i[78]
  PIN sports_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 255.720 450.000 256.320 ;
    END
  END sports_i[79]
  PIN sports_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 59.880 450.000 60.480 ;
    END
  END sports_i[7]
  PIN sports_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 258.440 450.000 259.040 ;
    END
  END sports_i[80]
  PIN sports_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 261.160 450.000 261.760 ;
    END
  END sports_i[81]
  PIN sports_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 263.880 450.000 264.480 ;
    END
  END sports_i[82]
  PIN sports_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 266.600 450.000 267.200 ;
    END
  END sports_i[83]
  PIN sports_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 269.320 450.000 269.920 ;
    END
  END sports_i[84]
  PIN sports_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 272.040 450.000 272.640 ;
    END
  END sports_i[85]
  PIN sports_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 274.760 450.000 275.360 ;
    END
  END sports_i[86]
  PIN sports_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 277.480 450.000 278.080 ;
    END
  END sports_i[87]
  PIN sports_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 280.200 450.000 280.800 ;
    END
  END sports_i[88]
  PIN sports_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 282.920 450.000 283.520 ;
    END
  END sports_i[89]
  PIN sports_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 62.600 450.000 63.200 ;
    END
  END sports_i[8]
  PIN sports_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 285.640 450.000 286.240 ;
    END
  END sports_i[90]
  PIN sports_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 288.360 450.000 288.960 ;
    END
  END sports_i[91]
  PIN sports_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 291.080 450.000 291.680 ;
    END
  END sports_i[92]
  PIN sports_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 293.800 450.000 294.400 ;
    END
  END sports_i[93]
  PIN sports_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 296.520 450.000 297.120 ;
    END
  END sports_i[94]
  PIN sports_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 299.240 450.000 299.840 ;
    END
  END sports_i[95]
  PIN sports_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 301.960 450.000 302.560 ;
    END
  END sports_i[96]
  PIN sports_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 304.680 450.000 305.280 ;
    END
  END sports_i[97]
  PIN sports_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 307.400 450.000 308.000 ;
    END
  END sports_i[98]
  PIN sports_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 446.000 310.120 450.000 310.720 ;
    END
  END sports_i[99]
  PIN sports_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 65.320 450.000 65.920 ;
    END
  END sports_i[9]
  PIN sports_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END sports_o[0]
  PIN sports_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END sports_o[100]
  PIN sports_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END sports_o[101]
  PIN sports_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END sports_o[102]
  PIN sports_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END sports_o[103]
  PIN sports_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END sports_o[104]
  PIN sports_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END sports_o[105]
  PIN sports_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END sports_o[106]
  PIN sports_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END sports_o[107]
  PIN sports_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END sports_o[108]
  PIN sports_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END sports_o[109]
  PIN sports_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END sports_o[10]
  PIN sports_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END sports_o[110]
  PIN sports_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END sports_o[111]
  PIN sports_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END sports_o[112]
  PIN sports_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END sports_o[113]
  PIN sports_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END sports_o[114]
  PIN sports_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END sports_o[115]
  PIN sports_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END sports_o[116]
  PIN sports_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END sports_o[117]
  PIN sports_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END sports_o[118]
  PIN sports_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END sports_o[119]
  PIN sports_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END sports_o[11]
  PIN sports_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END sports_o[120]
  PIN sports_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END sports_o[121]
  PIN sports_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END sports_o[122]
  PIN sports_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END sports_o[123]
  PIN sports_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END sports_o[124]
  PIN sports_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END sports_o[125]
  PIN sports_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END sports_o[126]
  PIN sports_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END sports_o[127]
  PIN sports_o[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END sports_o[128]
  PIN sports_o[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END sports_o[129]
  PIN sports_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END sports_o[12]
  PIN sports_o[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END sports_o[130]
  PIN sports_o[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END sports_o[131]
  PIN sports_o[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END sports_o[132]
  PIN sports_o[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END sports_o[133]
  PIN sports_o[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END sports_o[134]
  PIN sports_o[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END sports_o[135]
  PIN sports_o[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END sports_o[136]
  PIN sports_o[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END sports_o[137]
  PIN sports_o[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END sports_o[138]
  PIN sports_o[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END sports_o[139]
  PIN sports_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END sports_o[13]
  PIN sports_o[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END sports_o[140]
  PIN sports_o[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END sports_o[141]
  PIN sports_o[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END sports_o[142]
  PIN sports_o[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END sports_o[143]
  PIN sports_o[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END sports_o[144]
  PIN sports_o[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END sports_o[145]
  PIN sports_o[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END sports_o[146]
  PIN sports_o[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END sports_o[147]
  PIN sports_o[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END sports_o[148]
  PIN sports_o[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END sports_o[149]
  PIN sports_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END sports_o[14]
  PIN sports_o[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END sports_o[150]
  PIN sports_o[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END sports_o[151]
  PIN sports_o[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END sports_o[152]
  PIN sports_o[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END sports_o[153]
  PIN sports_o[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END sports_o[154]
  PIN sports_o[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END sports_o[155]
  PIN sports_o[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END sports_o[156]
  PIN sports_o[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END sports_o[157]
  PIN sports_o[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END sports_o[158]
  PIN sports_o[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END sports_o[159]
  PIN sports_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END sports_o[15]
  PIN sports_o[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END sports_o[160]
  PIN sports_o[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END sports_o[161]
  PIN sports_o[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END sports_o[162]
  PIN sports_o[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END sports_o[163]
  PIN sports_o[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END sports_o[164]
  PIN sports_o[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END sports_o[165]
  PIN sports_o[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END sports_o[166]
  PIN sports_o[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END sports_o[167]
  PIN sports_o[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END sports_o[168]
  PIN sports_o[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END sports_o[169]
  PIN sports_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END sports_o[16]
  PIN sports_o[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END sports_o[170]
  PIN sports_o[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END sports_o[171]
  PIN sports_o[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END sports_o[172]
  PIN sports_o[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END sports_o[173]
  PIN sports_o[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END sports_o[174]
  PIN sports_o[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END sports_o[175]
  PIN sports_o[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END sports_o[176]
  PIN sports_o[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END sports_o[177]
  PIN sports_o[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END sports_o[178]
  PIN sports_o[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END sports_o[179]
  PIN sports_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END sports_o[17]
  PIN sports_o[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END sports_o[180]
  PIN sports_o[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END sports_o[181]
  PIN sports_o[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END sports_o[182]
  PIN sports_o[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END sports_o[183]
  PIN sports_o[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END sports_o[184]
  PIN sports_o[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END sports_o[185]
  PIN sports_o[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END sports_o[186]
  PIN sports_o[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END sports_o[187]
  PIN sports_o[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END sports_o[188]
  PIN sports_o[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END sports_o[189]
  PIN sports_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END sports_o[18]
  PIN sports_o[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END sports_o[190]
  PIN sports_o[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END sports_o[191]
  PIN sports_o[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END sports_o[192]
  PIN sports_o[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END sports_o[193]
  PIN sports_o[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END sports_o[194]
  PIN sports_o[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END sports_o[195]
  PIN sports_o[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END sports_o[196]
  PIN sports_o[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END sports_o[197]
  PIN sports_o[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END sports_o[198]
  PIN sports_o[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END sports_o[199]
  PIN sports_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END sports_o[19]
  PIN sports_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END sports_o[1]
  PIN sports_o[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END sports_o[200]
  PIN sports_o[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END sports_o[201]
  PIN sports_o[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END sports_o[202]
  PIN sports_o[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END sports_o[203]
  PIN sports_o[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END sports_o[204]
  PIN sports_o[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END sports_o[205]
  PIN sports_o[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END sports_o[206]
  PIN sports_o[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END sports_o[207]
  PIN sports_o[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END sports_o[208]
  PIN sports_o[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END sports_o[209]
  PIN sports_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END sports_o[20]
  PIN sports_o[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END sports_o[210]
  PIN sports_o[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END sports_o[211]
  PIN sports_o[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END sports_o[212]
  PIN sports_o[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END sports_o[213]
  PIN sports_o[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END sports_o[214]
  PIN sports_o[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END sports_o[215]
  PIN sports_o[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END sports_o[216]
  PIN sports_o[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END sports_o[217]
  PIN sports_o[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END sports_o[218]
  PIN sports_o[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END sports_o[219]
  PIN sports_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END sports_o[21]
  PIN sports_o[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END sports_o[220]
  PIN sports_o[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END sports_o[221]
  PIN sports_o[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END sports_o[222]
  PIN sports_o[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END sports_o[223]
  PIN sports_o[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END sports_o[224]
  PIN sports_o[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END sports_o[225]
  PIN sports_o[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END sports_o[226]
  PIN sports_o[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END sports_o[227]
  PIN sports_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END sports_o[22]
  PIN sports_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END sports_o[23]
  PIN sports_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END sports_o[24]
  PIN sports_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END sports_o[25]
  PIN sports_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END sports_o[26]
  PIN sports_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END sports_o[27]
  PIN sports_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END sports_o[28]
  PIN sports_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END sports_o[29]
  PIN sports_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END sports_o[2]
  PIN sports_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END sports_o[30]
  PIN sports_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END sports_o[31]
  PIN sports_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END sports_o[32]
  PIN sports_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END sports_o[33]
  PIN sports_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END sports_o[34]
  PIN sports_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END sports_o[35]
  PIN sports_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END sports_o[36]
  PIN sports_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END sports_o[37]
  PIN sports_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END sports_o[38]
  PIN sports_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END sports_o[39]
  PIN sports_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END sports_o[3]
  PIN sports_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END sports_o[40]
  PIN sports_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END sports_o[41]
  PIN sports_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END sports_o[42]
  PIN sports_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END sports_o[43]
  PIN sports_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END sports_o[44]
  PIN sports_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END sports_o[45]
  PIN sports_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END sports_o[46]
  PIN sports_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END sports_o[47]
  PIN sports_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END sports_o[48]
  PIN sports_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END sports_o[49]
  PIN sports_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END sports_o[4]
  PIN sports_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END sports_o[50]
  PIN sports_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END sports_o[51]
  PIN sports_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END sports_o[52]
  PIN sports_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END sports_o[53]
  PIN sports_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END sports_o[54]
  PIN sports_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END sports_o[55]
  PIN sports_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END sports_o[56]
  PIN sports_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END sports_o[57]
  PIN sports_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END sports_o[58]
  PIN sports_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END sports_o[59]
  PIN sports_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END sports_o[5]
  PIN sports_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END sports_o[60]
  PIN sports_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END sports_o[61]
  PIN sports_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END sports_o[62]
  PIN sports_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END sports_o[63]
  PIN sports_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END sports_o[64]
  PIN sports_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END sports_o[65]
  PIN sports_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END sports_o[66]
  PIN sports_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END sports_o[67]
  PIN sports_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END sports_o[68]
  PIN sports_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END sports_o[69]
  PIN sports_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END sports_o[6]
  PIN sports_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END sports_o[70]
  PIN sports_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END sports_o[71]
  PIN sports_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END sports_o[72]
  PIN sports_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END sports_o[73]
  PIN sports_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END sports_o[74]
  PIN sports_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END sports_o[75]
  PIN sports_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END sports_o[76]
  PIN sports_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END sports_o[77]
  PIN sports_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END sports_o[78]
  PIN sports_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END sports_o[79]
  PIN sports_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END sports_o[7]
  PIN sports_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END sports_o[80]
  PIN sports_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END sports_o[81]
  PIN sports_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END sports_o[82]
  PIN sports_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END sports_o[83]
  PIN sports_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END sports_o[84]
  PIN sports_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END sports_o[85]
  PIN sports_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END sports_o[86]
  PIN sports_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END sports_o[87]
  PIN sports_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END sports_o[88]
  PIN sports_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END sports_o[89]
  PIN sports_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END sports_o[8]
  PIN sports_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END sports_o[90]
  PIN sports_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END sports_o[91]
  PIN sports_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END sports_o[92]
  PIN sports_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END sports_o[93]
  PIN sports_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END sports_o[94]
  PIN sports_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END sports_o[95]
  PIN sports_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END sports_o[96]
  PIN sports_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END sports_o[97]
  PIN sports_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END sports_o[98]
  PIN sports_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END sports_o[99]
  PIN sports_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END sports_o[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 438.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 438.160 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 444.360 438.005 ;
      LAYER met1 ;
        RECT 0.070 4.800 449.810 449.780 ;
      LAYER met2 ;
        RECT 0.100 445.720 13.610 449.810 ;
        RECT 14.450 445.720 15.450 449.810 ;
        RECT 16.290 445.720 17.290 449.810 ;
        RECT 18.130 445.720 19.130 449.810 ;
        RECT 19.970 445.720 20.970 449.810 ;
        RECT 21.810 445.720 22.810 449.810 ;
        RECT 23.650 445.720 24.650 449.810 ;
        RECT 25.490 445.720 26.490 449.810 ;
        RECT 27.330 445.720 28.330 449.810 ;
        RECT 29.170 445.720 30.170 449.810 ;
        RECT 31.010 445.720 32.010 449.810 ;
        RECT 32.850 445.720 33.850 449.810 ;
        RECT 34.690 445.720 35.690 449.810 ;
        RECT 36.530 445.720 37.530 449.810 ;
        RECT 38.370 445.720 39.370 449.810 ;
        RECT 40.210 445.720 41.210 449.810 ;
        RECT 42.050 445.720 43.050 449.810 ;
        RECT 43.890 445.720 44.890 449.810 ;
        RECT 45.730 445.720 46.730 449.810 ;
        RECT 47.570 445.720 48.570 449.810 ;
        RECT 49.410 445.720 50.410 449.810 ;
        RECT 51.250 445.720 52.250 449.810 ;
        RECT 53.090 445.720 54.090 449.810 ;
        RECT 54.930 445.720 55.930 449.810 ;
        RECT 56.770 445.720 57.770 449.810 ;
        RECT 58.610 445.720 59.610 449.810 ;
        RECT 60.450 445.720 61.450 449.810 ;
        RECT 62.290 445.720 63.290 449.810 ;
        RECT 64.130 445.720 65.130 449.810 ;
        RECT 65.970 445.720 66.970 449.810 ;
        RECT 67.810 445.720 68.810 449.810 ;
        RECT 69.650 445.720 70.650 449.810 ;
        RECT 71.490 445.720 72.490 449.810 ;
        RECT 73.330 445.720 74.330 449.810 ;
        RECT 75.170 445.720 76.170 449.810 ;
        RECT 77.010 445.720 78.010 449.810 ;
        RECT 78.850 445.720 79.850 449.810 ;
        RECT 80.690 445.720 81.690 449.810 ;
        RECT 82.530 445.720 83.530 449.810 ;
        RECT 84.370 445.720 85.370 449.810 ;
        RECT 86.210 445.720 87.210 449.810 ;
        RECT 88.050 445.720 89.050 449.810 ;
        RECT 89.890 445.720 90.890 449.810 ;
        RECT 91.730 445.720 92.730 449.810 ;
        RECT 93.570 445.720 94.570 449.810 ;
        RECT 95.410 445.720 96.410 449.810 ;
        RECT 97.250 445.720 98.250 449.810 ;
        RECT 99.090 445.720 100.090 449.810 ;
        RECT 100.930 445.720 101.930 449.810 ;
        RECT 102.770 445.720 103.770 449.810 ;
        RECT 104.610 445.720 105.610 449.810 ;
        RECT 106.450 445.720 107.450 449.810 ;
        RECT 108.290 445.720 109.290 449.810 ;
        RECT 110.130 445.720 111.130 449.810 ;
        RECT 111.970 445.720 112.970 449.810 ;
        RECT 113.810 445.720 114.810 449.810 ;
        RECT 115.650 445.720 116.650 449.810 ;
        RECT 117.490 445.720 118.490 449.810 ;
        RECT 119.330 445.720 120.330 449.810 ;
        RECT 121.170 445.720 122.170 449.810 ;
        RECT 123.010 445.720 124.010 449.810 ;
        RECT 124.850 445.720 125.850 449.810 ;
        RECT 126.690 445.720 127.690 449.810 ;
        RECT 128.530 445.720 129.530 449.810 ;
        RECT 130.370 445.720 131.370 449.810 ;
        RECT 132.210 445.720 133.210 449.810 ;
        RECT 134.050 445.720 135.050 449.810 ;
        RECT 135.890 445.720 136.890 449.810 ;
        RECT 137.730 445.720 138.730 449.810 ;
        RECT 139.570 445.720 140.570 449.810 ;
        RECT 141.410 445.720 142.410 449.810 ;
        RECT 143.250 445.720 144.250 449.810 ;
        RECT 145.090 445.720 146.090 449.810 ;
        RECT 146.930 445.720 147.930 449.810 ;
        RECT 148.770 445.720 149.770 449.810 ;
        RECT 150.610 445.720 151.610 449.810 ;
        RECT 152.450 445.720 153.450 449.810 ;
        RECT 154.290 445.720 155.290 449.810 ;
        RECT 156.130 445.720 157.130 449.810 ;
        RECT 157.970 445.720 158.970 449.810 ;
        RECT 159.810 445.720 160.810 449.810 ;
        RECT 161.650 445.720 162.650 449.810 ;
        RECT 163.490 445.720 164.490 449.810 ;
        RECT 165.330 445.720 166.330 449.810 ;
        RECT 167.170 445.720 168.170 449.810 ;
        RECT 169.010 445.720 170.010 449.810 ;
        RECT 170.850 445.720 171.850 449.810 ;
        RECT 172.690 445.720 173.690 449.810 ;
        RECT 174.530 445.720 175.530 449.810 ;
        RECT 176.370 445.720 177.370 449.810 ;
        RECT 178.210 445.720 179.210 449.810 ;
        RECT 180.050 445.720 181.050 449.810 ;
        RECT 181.890 445.720 182.890 449.810 ;
        RECT 183.730 445.720 184.730 449.810 ;
        RECT 185.570 445.720 186.570 449.810 ;
        RECT 187.410 445.720 188.410 449.810 ;
        RECT 189.250 445.720 190.250 449.810 ;
        RECT 191.090 445.720 192.090 449.810 ;
        RECT 192.930 445.720 193.930 449.810 ;
        RECT 194.770 445.720 195.770 449.810 ;
        RECT 196.610 445.720 197.610 449.810 ;
        RECT 198.450 445.720 199.450 449.810 ;
        RECT 200.290 445.720 201.290 449.810 ;
        RECT 202.130 445.720 203.130 449.810 ;
        RECT 203.970 445.720 204.970 449.810 ;
        RECT 205.810 445.720 206.810 449.810 ;
        RECT 207.650 445.720 208.650 449.810 ;
        RECT 209.490 445.720 210.490 449.810 ;
        RECT 211.330 445.720 212.330 449.810 ;
        RECT 213.170 445.720 214.170 449.810 ;
        RECT 215.010 445.720 216.010 449.810 ;
        RECT 216.850 445.720 217.850 449.810 ;
        RECT 218.690 445.720 219.690 449.810 ;
        RECT 220.530 445.720 221.530 449.810 ;
        RECT 222.370 445.720 223.370 449.810 ;
        RECT 224.210 445.720 225.210 449.810 ;
        RECT 226.050 445.720 227.050 449.810 ;
        RECT 227.890 445.720 228.890 449.810 ;
        RECT 229.730 445.720 230.730 449.810 ;
        RECT 231.570 445.720 232.570 449.810 ;
        RECT 233.410 445.720 234.410 449.810 ;
        RECT 235.250 445.720 236.250 449.810 ;
        RECT 237.090 445.720 238.090 449.810 ;
        RECT 238.930 445.720 239.930 449.810 ;
        RECT 240.770 445.720 241.770 449.810 ;
        RECT 242.610 445.720 243.610 449.810 ;
        RECT 244.450 445.720 245.450 449.810 ;
        RECT 246.290 445.720 247.290 449.810 ;
        RECT 248.130 445.720 249.130 449.810 ;
        RECT 249.970 445.720 250.970 449.810 ;
        RECT 251.810 445.720 252.810 449.810 ;
        RECT 253.650 445.720 254.650 449.810 ;
        RECT 255.490 445.720 256.490 449.810 ;
        RECT 257.330 445.720 258.330 449.810 ;
        RECT 259.170 445.720 260.170 449.810 ;
        RECT 261.010 445.720 262.010 449.810 ;
        RECT 262.850 445.720 263.850 449.810 ;
        RECT 264.690 445.720 265.690 449.810 ;
        RECT 266.530 445.720 267.530 449.810 ;
        RECT 268.370 445.720 269.370 449.810 ;
        RECT 270.210 445.720 271.210 449.810 ;
        RECT 272.050 445.720 273.050 449.810 ;
        RECT 273.890 445.720 274.890 449.810 ;
        RECT 275.730 445.720 276.730 449.810 ;
        RECT 277.570 445.720 278.570 449.810 ;
        RECT 279.410 445.720 280.410 449.810 ;
        RECT 281.250 445.720 282.250 449.810 ;
        RECT 283.090 445.720 284.090 449.810 ;
        RECT 284.930 445.720 285.930 449.810 ;
        RECT 286.770 445.720 287.770 449.810 ;
        RECT 288.610 445.720 289.610 449.810 ;
        RECT 290.450 445.720 291.450 449.810 ;
        RECT 292.290 445.720 293.290 449.810 ;
        RECT 294.130 445.720 295.130 449.810 ;
        RECT 295.970 445.720 296.970 449.810 ;
        RECT 297.810 445.720 298.810 449.810 ;
        RECT 299.650 445.720 300.650 449.810 ;
        RECT 301.490 445.720 302.490 449.810 ;
        RECT 303.330 445.720 304.330 449.810 ;
        RECT 305.170 445.720 306.170 449.810 ;
        RECT 307.010 445.720 308.010 449.810 ;
        RECT 308.850 445.720 309.850 449.810 ;
        RECT 310.690 445.720 311.690 449.810 ;
        RECT 312.530 445.720 313.530 449.810 ;
        RECT 314.370 445.720 315.370 449.810 ;
        RECT 316.210 445.720 317.210 449.810 ;
        RECT 318.050 445.720 319.050 449.810 ;
        RECT 319.890 445.720 320.890 449.810 ;
        RECT 321.730 445.720 322.730 449.810 ;
        RECT 323.570 445.720 324.570 449.810 ;
        RECT 325.410 445.720 326.410 449.810 ;
        RECT 327.250 445.720 328.250 449.810 ;
        RECT 329.090 445.720 330.090 449.810 ;
        RECT 330.930 445.720 331.930 449.810 ;
        RECT 332.770 445.720 333.770 449.810 ;
        RECT 334.610 445.720 335.610 449.810 ;
        RECT 336.450 445.720 337.450 449.810 ;
        RECT 338.290 445.720 339.290 449.810 ;
        RECT 340.130 445.720 341.130 449.810 ;
        RECT 341.970 445.720 342.970 449.810 ;
        RECT 343.810 445.720 344.810 449.810 ;
        RECT 345.650 445.720 346.650 449.810 ;
        RECT 347.490 445.720 348.490 449.810 ;
        RECT 349.330 445.720 350.330 449.810 ;
        RECT 351.170 445.720 352.170 449.810 ;
        RECT 353.010 445.720 354.010 449.810 ;
        RECT 354.850 445.720 355.850 449.810 ;
        RECT 356.690 445.720 357.690 449.810 ;
        RECT 358.530 445.720 359.530 449.810 ;
        RECT 360.370 445.720 361.370 449.810 ;
        RECT 362.210 445.720 363.210 449.810 ;
        RECT 364.050 445.720 365.050 449.810 ;
        RECT 365.890 445.720 366.890 449.810 ;
        RECT 367.730 445.720 368.730 449.810 ;
        RECT 369.570 445.720 370.570 449.810 ;
        RECT 371.410 445.720 372.410 449.810 ;
        RECT 373.250 445.720 374.250 449.810 ;
        RECT 375.090 445.720 376.090 449.810 ;
        RECT 376.930 445.720 377.930 449.810 ;
        RECT 378.770 445.720 379.770 449.810 ;
        RECT 380.610 445.720 381.610 449.810 ;
        RECT 382.450 445.720 383.450 449.810 ;
        RECT 384.290 445.720 385.290 449.810 ;
        RECT 386.130 445.720 387.130 449.810 ;
        RECT 387.970 445.720 388.970 449.810 ;
        RECT 389.810 445.720 390.810 449.810 ;
        RECT 391.650 445.720 392.650 449.810 ;
        RECT 393.490 445.720 394.490 449.810 ;
        RECT 395.330 445.720 396.330 449.810 ;
        RECT 397.170 445.720 398.170 449.810 ;
        RECT 399.010 445.720 400.010 449.810 ;
        RECT 400.850 445.720 401.850 449.810 ;
        RECT 402.690 445.720 403.690 449.810 ;
        RECT 404.530 445.720 405.530 449.810 ;
        RECT 406.370 445.720 407.370 449.810 ;
        RECT 408.210 445.720 409.210 449.810 ;
        RECT 410.050 445.720 411.050 449.810 ;
        RECT 411.890 445.720 412.890 449.810 ;
        RECT 413.730 445.720 414.730 449.810 ;
        RECT 415.570 445.720 416.570 449.810 ;
        RECT 417.410 445.720 418.410 449.810 ;
        RECT 419.250 445.720 420.250 449.810 ;
        RECT 421.090 445.720 422.090 449.810 ;
        RECT 422.930 445.720 423.930 449.810 ;
        RECT 424.770 445.720 425.770 449.810 ;
        RECT 426.610 445.720 427.610 449.810 ;
        RECT 428.450 445.720 429.450 449.810 ;
        RECT 430.290 445.720 431.290 449.810 ;
        RECT 432.130 445.720 433.130 449.810 ;
        RECT 433.970 445.720 434.970 449.810 ;
        RECT 435.810 445.720 449.780 449.810 ;
        RECT 0.100 4.280 449.780 445.720 ;
        RECT 0.100 3.670 7.170 4.280 ;
        RECT 8.010 3.670 10.390 4.280 ;
        RECT 11.230 3.670 13.610 4.280 ;
        RECT 14.450 3.670 16.830 4.280 ;
        RECT 17.670 3.670 20.050 4.280 ;
        RECT 20.890 3.670 23.270 4.280 ;
        RECT 24.110 3.670 26.490 4.280 ;
        RECT 27.330 3.670 29.710 4.280 ;
        RECT 30.550 3.670 32.930 4.280 ;
        RECT 33.770 3.670 36.150 4.280 ;
        RECT 36.990 3.670 39.370 4.280 ;
        RECT 40.210 3.670 42.590 4.280 ;
        RECT 43.430 3.670 45.810 4.280 ;
        RECT 46.650 3.670 49.030 4.280 ;
        RECT 49.870 3.670 52.250 4.280 ;
        RECT 53.090 3.670 55.470 4.280 ;
        RECT 56.310 3.670 58.690 4.280 ;
        RECT 59.530 3.670 61.910 4.280 ;
        RECT 62.750 3.670 65.130 4.280 ;
        RECT 65.970 3.670 68.350 4.280 ;
        RECT 69.190 3.670 71.570 4.280 ;
        RECT 72.410 3.670 74.790 4.280 ;
        RECT 75.630 3.670 78.010 4.280 ;
        RECT 78.850 3.670 81.230 4.280 ;
        RECT 82.070 3.670 84.450 4.280 ;
        RECT 85.290 3.670 87.670 4.280 ;
        RECT 88.510 3.670 90.890 4.280 ;
        RECT 91.730 3.670 94.110 4.280 ;
        RECT 94.950 3.670 97.330 4.280 ;
        RECT 98.170 3.670 100.550 4.280 ;
        RECT 101.390 3.670 103.770 4.280 ;
        RECT 104.610 3.670 106.990 4.280 ;
        RECT 107.830 3.670 110.210 4.280 ;
        RECT 111.050 3.670 113.430 4.280 ;
        RECT 114.270 3.670 116.650 4.280 ;
        RECT 117.490 3.670 119.870 4.280 ;
        RECT 120.710 3.670 123.090 4.280 ;
        RECT 123.930 3.670 126.310 4.280 ;
        RECT 127.150 3.670 129.530 4.280 ;
        RECT 130.370 3.670 132.750 4.280 ;
        RECT 133.590 3.670 135.970 4.280 ;
        RECT 136.810 3.670 139.190 4.280 ;
        RECT 140.030 3.670 142.410 4.280 ;
        RECT 143.250 3.670 145.630 4.280 ;
        RECT 146.470 3.670 148.850 4.280 ;
        RECT 149.690 3.670 152.070 4.280 ;
        RECT 152.910 3.670 155.290 4.280 ;
        RECT 156.130 3.670 158.510 4.280 ;
        RECT 159.350 3.670 161.730 4.280 ;
        RECT 162.570 3.670 164.950 4.280 ;
        RECT 165.790 3.670 168.170 4.280 ;
        RECT 169.010 3.670 171.390 4.280 ;
        RECT 172.230 3.670 174.610 4.280 ;
        RECT 175.450 3.670 177.830 4.280 ;
        RECT 178.670 3.670 181.050 4.280 ;
        RECT 181.890 3.670 184.270 4.280 ;
        RECT 185.110 3.670 187.490 4.280 ;
        RECT 188.330 3.670 190.710 4.280 ;
        RECT 191.550 3.670 193.930 4.280 ;
        RECT 194.770 3.670 197.150 4.280 ;
        RECT 197.990 3.670 200.370 4.280 ;
        RECT 201.210 3.670 203.590 4.280 ;
        RECT 204.430 3.670 206.810 4.280 ;
        RECT 207.650 3.670 210.030 4.280 ;
        RECT 210.870 3.670 213.250 4.280 ;
        RECT 214.090 3.670 216.470 4.280 ;
        RECT 217.310 3.670 219.690 4.280 ;
        RECT 220.530 3.670 222.910 4.280 ;
        RECT 223.750 3.670 226.130 4.280 ;
        RECT 226.970 3.670 229.350 4.280 ;
        RECT 230.190 3.670 232.570 4.280 ;
        RECT 233.410 3.670 235.790 4.280 ;
        RECT 236.630 3.670 239.010 4.280 ;
        RECT 239.850 3.670 242.230 4.280 ;
        RECT 243.070 3.670 245.450 4.280 ;
        RECT 246.290 3.670 248.670 4.280 ;
        RECT 249.510 3.670 251.890 4.280 ;
        RECT 252.730 3.670 255.110 4.280 ;
        RECT 255.950 3.670 258.330 4.280 ;
        RECT 259.170 3.670 261.550 4.280 ;
        RECT 262.390 3.670 264.770 4.280 ;
        RECT 265.610 3.670 267.990 4.280 ;
        RECT 268.830 3.670 271.210 4.280 ;
        RECT 272.050 3.670 274.430 4.280 ;
        RECT 275.270 3.670 277.650 4.280 ;
        RECT 278.490 3.670 280.870 4.280 ;
        RECT 281.710 3.670 284.090 4.280 ;
        RECT 284.930 3.670 287.310 4.280 ;
        RECT 288.150 3.670 290.530 4.280 ;
        RECT 291.370 3.670 293.750 4.280 ;
        RECT 294.590 3.670 296.970 4.280 ;
        RECT 297.810 3.670 300.190 4.280 ;
        RECT 301.030 3.670 303.410 4.280 ;
        RECT 304.250 3.670 306.630 4.280 ;
        RECT 307.470 3.670 309.850 4.280 ;
        RECT 310.690 3.670 313.070 4.280 ;
        RECT 313.910 3.670 316.290 4.280 ;
        RECT 317.130 3.670 319.510 4.280 ;
        RECT 320.350 3.670 322.730 4.280 ;
        RECT 323.570 3.670 325.950 4.280 ;
        RECT 326.790 3.670 329.170 4.280 ;
        RECT 330.010 3.670 332.390 4.280 ;
        RECT 333.230 3.670 335.610 4.280 ;
        RECT 336.450 3.670 338.830 4.280 ;
        RECT 339.670 3.670 342.050 4.280 ;
        RECT 342.890 3.670 345.270 4.280 ;
        RECT 346.110 3.670 348.490 4.280 ;
        RECT 349.330 3.670 351.710 4.280 ;
        RECT 352.550 3.670 354.930 4.280 ;
        RECT 355.770 3.670 358.150 4.280 ;
        RECT 358.990 3.670 361.370 4.280 ;
        RECT 362.210 3.670 364.590 4.280 ;
        RECT 365.430 3.670 367.810 4.280 ;
        RECT 368.650 3.670 371.030 4.280 ;
        RECT 371.870 3.670 374.250 4.280 ;
        RECT 375.090 3.670 377.470 4.280 ;
        RECT 378.310 3.670 380.690 4.280 ;
        RECT 381.530 3.670 383.910 4.280 ;
        RECT 384.750 3.670 387.130 4.280 ;
        RECT 387.970 3.670 390.350 4.280 ;
        RECT 391.190 3.670 393.570 4.280 ;
        RECT 394.410 3.670 396.790 4.280 ;
        RECT 397.630 3.670 400.010 4.280 ;
        RECT 400.850 3.670 403.230 4.280 ;
        RECT 404.070 3.670 406.450 4.280 ;
        RECT 407.290 3.670 409.670 4.280 ;
        RECT 410.510 3.670 412.890 4.280 ;
        RECT 413.730 3.670 416.110 4.280 ;
        RECT 416.950 3.670 419.330 4.280 ;
        RECT 420.170 3.670 422.550 4.280 ;
        RECT 423.390 3.670 425.770 4.280 ;
        RECT 426.610 3.670 428.990 4.280 ;
        RECT 429.830 3.670 432.210 4.280 ;
        RECT 433.050 3.670 435.430 4.280 ;
        RECT 436.270 3.670 438.650 4.280 ;
        RECT 439.490 3.670 441.870 4.280 ;
        RECT 442.710 3.670 449.780 4.280 ;
      LAYER met3 ;
        RECT 4.000 409.040 446.135 449.305 ;
        RECT 4.000 407.640 445.600 409.040 ;
        RECT 4.000 406.320 446.135 407.640 ;
        RECT 4.000 404.920 445.600 406.320 ;
        RECT 4.000 403.600 446.135 404.920 ;
        RECT 4.000 402.200 445.600 403.600 ;
        RECT 4.000 400.880 446.135 402.200 ;
        RECT 4.000 399.480 445.600 400.880 ;
        RECT 4.000 398.160 446.135 399.480 ;
        RECT 4.000 396.760 445.600 398.160 ;
        RECT 4.000 395.440 446.135 396.760 ;
        RECT 4.000 394.040 445.600 395.440 ;
        RECT 4.000 392.720 446.135 394.040 ;
        RECT 4.000 391.320 445.600 392.720 ;
        RECT 4.000 390.000 446.135 391.320 ;
        RECT 4.000 388.600 445.600 390.000 ;
        RECT 4.000 387.280 446.135 388.600 ;
        RECT 4.000 385.880 445.600 387.280 ;
        RECT 4.000 384.560 446.135 385.880 ;
        RECT 4.000 383.160 445.600 384.560 ;
        RECT 4.000 381.840 446.135 383.160 ;
        RECT 4.000 380.440 445.600 381.840 ;
        RECT 4.000 379.120 446.135 380.440 ;
        RECT 4.400 377.720 445.600 379.120 ;
        RECT 4.400 376.400 446.135 377.720 ;
        RECT 4.400 375.000 445.600 376.400 ;
        RECT 4.400 373.680 446.135 375.000 ;
        RECT 4.400 372.280 445.600 373.680 ;
        RECT 4.400 370.960 446.135 372.280 ;
        RECT 4.400 369.560 445.600 370.960 ;
        RECT 4.400 368.240 446.135 369.560 ;
        RECT 4.400 366.840 445.600 368.240 ;
        RECT 4.400 365.520 446.135 366.840 ;
        RECT 4.400 364.120 445.600 365.520 ;
        RECT 4.400 362.800 446.135 364.120 ;
        RECT 4.400 361.400 445.600 362.800 ;
        RECT 4.400 360.080 446.135 361.400 ;
        RECT 4.400 358.680 445.600 360.080 ;
        RECT 4.400 357.360 446.135 358.680 ;
        RECT 4.400 355.960 445.600 357.360 ;
        RECT 4.400 354.640 446.135 355.960 ;
        RECT 4.400 353.240 445.600 354.640 ;
        RECT 4.400 351.920 446.135 353.240 ;
        RECT 4.400 350.520 445.600 351.920 ;
        RECT 4.400 349.200 446.135 350.520 ;
        RECT 4.400 347.800 445.600 349.200 ;
        RECT 4.400 346.480 446.135 347.800 ;
        RECT 4.400 345.080 445.600 346.480 ;
        RECT 4.400 343.760 446.135 345.080 ;
        RECT 4.400 342.360 445.600 343.760 ;
        RECT 4.400 341.040 446.135 342.360 ;
        RECT 4.400 339.640 445.600 341.040 ;
        RECT 4.400 338.320 446.135 339.640 ;
        RECT 4.400 336.920 445.600 338.320 ;
        RECT 4.400 335.600 446.135 336.920 ;
        RECT 4.400 334.200 445.600 335.600 ;
        RECT 4.400 332.880 446.135 334.200 ;
        RECT 4.400 331.480 445.600 332.880 ;
        RECT 4.400 330.160 446.135 331.480 ;
        RECT 4.400 328.760 445.600 330.160 ;
        RECT 4.400 327.440 446.135 328.760 ;
        RECT 4.400 326.040 445.600 327.440 ;
        RECT 4.400 324.720 446.135 326.040 ;
        RECT 4.400 323.320 445.600 324.720 ;
        RECT 4.400 322.000 446.135 323.320 ;
        RECT 4.400 320.600 445.600 322.000 ;
        RECT 4.400 319.280 446.135 320.600 ;
        RECT 4.400 317.880 445.600 319.280 ;
        RECT 4.400 316.560 446.135 317.880 ;
        RECT 4.400 315.160 445.600 316.560 ;
        RECT 4.400 313.840 446.135 315.160 ;
        RECT 4.400 312.440 445.600 313.840 ;
        RECT 4.400 311.120 446.135 312.440 ;
        RECT 4.400 309.720 445.600 311.120 ;
        RECT 4.400 308.400 446.135 309.720 ;
        RECT 4.400 307.000 445.600 308.400 ;
        RECT 4.400 305.680 446.135 307.000 ;
        RECT 4.400 304.280 445.600 305.680 ;
        RECT 4.400 302.960 446.135 304.280 ;
        RECT 4.400 301.560 445.600 302.960 ;
        RECT 4.400 300.240 446.135 301.560 ;
        RECT 4.400 298.840 445.600 300.240 ;
        RECT 4.400 297.520 446.135 298.840 ;
        RECT 4.400 296.120 445.600 297.520 ;
        RECT 4.400 294.800 446.135 296.120 ;
        RECT 4.400 293.400 445.600 294.800 ;
        RECT 4.400 292.080 446.135 293.400 ;
        RECT 4.400 290.680 445.600 292.080 ;
        RECT 4.400 289.360 446.135 290.680 ;
        RECT 4.400 287.960 445.600 289.360 ;
        RECT 4.400 286.640 446.135 287.960 ;
        RECT 4.400 285.240 445.600 286.640 ;
        RECT 4.400 283.920 446.135 285.240 ;
        RECT 4.400 282.520 445.600 283.920 ;
        RECT 4.400 281.200 446.135 282.520 ;
        RECT 4.400 279.800 445.600 281.200 ;
        RECT 4.400 278.480 446.135 279.800 ;
        RECT 4.400 277.080 445.600 278.480 ;
        RECT 4.400 275.760 446.135 277.080 ;
        RECT 4.400 274.360 445.600 275.760 ;
        RECT 4.400 273.040 446.135 274.360 ;
        RECT 4.400 271.640 445.600 273.040 ;
        RECT 4.400 270.320 446.135 271.640 ;
        RECT 4.400 268.920 445.600 270.320 ;
        RECT 4.400 267.600 446.135 268.920 ;
        RECT 4.400 266.200 445.600 267.600 ;
        RECT 4.400 264.880 446.135 266.200 ;
        RECT 4.400 263.480 445.600 264.880 ;
        RECT 4.400 262.160 446.135 263.480 ;
        RECT 4.400 260.760 445.600 262.160 ;
        RECT 4.400 259.440 446.135 260.760 ;
        RECT 4.400 258.040 445.600 259.440 ;
        RECT 4.400 256.720 446.135 258.040 ;
        RECT 4.400 255.320 445.600 256.720 ;
        RECT 4.400 254.000 446.135 255.320 ;
        RECT 4.400 252.600 445.600 254.000 ;
        RECT 4.400 251.280 446.135 252.600 ;
        RECT 4.400 249.880 445.600 251.280 ;
        RECT 4.400 248.560 446.135 249.880 ;
        RECT 4.400 247.160 445.600 248.560 ;
        RECT 4.400 245.840 446.135 247.160 ;
        RECT 4.400 244.440 445.600 245.840 ;
        RECT 4.400 243.120 446.135 244.440 ;
        RECT 4.400 241.720 445.600 243.120 ;
        RECT 4.400 240.400 446.135 241.720 ;
        RECT 4.400 239.000 445.600 240.400 ;
        RECT 4.400 237.680 446.135 239.000 ;
        RECT 4.400 236.280 445.600 237.680 ;
        RECT 4.400 234.960 446.135 236.280 ;
        RECT 4.400 233.560 445.600 234.960 ;
        RECT 4.400 232.240 446.135 233.560 ;
        RECT 4.400 230.840 445.600 232.240 ;
        RECT 4.400 229.520 446.135 230.840 ;
        RECT 4.400 228.120 445.600 229.520 ;
        RECT 4.400 226.800 446.135 228.120 ;
        RECT 4.400 225.400 445.600 226.800 ;
        RECT 4.400 224.080 446.135 225.400 ;
        RECT 4.400 222.680 445.600 224.080 ;
        RECT 4.400 221.360 446.135 222.680 ;
        RECT 4.400 219.960 445.600 221.360 ;
        RECT 4.400 218.640 446.135 219.960 ;
        RECT 4.400 217.240 445.600 218.640 ;
        RECT 4.400 215.920 446.135 217.240 ;
        RECT 4.400 214.520 445.600 215.920 ;
        RECT 4.400 213.200 446.135 214.520 ;
        RECT 4.400 211.800 445.600 213.200 ;
        RECT 4.400 210.480 446.135 211.800 ;
        RECT 4.400 209.080 445.600 210.480 ;
        RECT 4.400 207.760 446.135 209.080 ;
        RECT 4.400 206.360 445.600 207.760 ;
        RECT 4.400 205.040 446.135 206.360 ;
        RECT 4.400 203.640 445.600 205.040 ;
        RECT 4.400 202.320 446.135 203.640 ;
        RECT 4.400 200.920 445.600 202.320 ;
        RECT 4.400 199.600 446.135 200.920 ;
        RECT 4.400 198.200 445.600 199.600 ;
        RECT 4.400 196.880 446.135 198.200 ;
        RECT 4.400 195.480 445.600 196.880 ;
        RECT 4.400 194.160 446.135 195.480 ;
        RECT 4.400 192.760 445.600 194.160 ;
        RECT 4.400 191.440 446.135 192.760 ;
        RECT 4.400 190.040 445.600 191.440 ;
        RECT 4.400 188.720 446.135 190.040 ;
        RECT 4.400 187.320 445.600 188.720 ;
        RECT 4.400 186.000 446.135 187.320 ;
        RECT 4.400 184.600 445.600 186.000 ;
        RECT 4.400 183.280 446.135 184.600 ;
        RECT 4.400 181.880 445.600 183.280 ;
        RECT 4.400 180.560 446.135 181.880 ;
        RECT 4.400 179.160 445.600 180.560 ;
        RECT 4.400 177.840 446.135 179.160 ;
        RECT 4.400 176.440 445.600 177.840 ;
        RECT 4.400 175.120 446.135 176.440 ;
        RECT 4.400 173.720 445.600 175.120 ;
        RECT 4.400 172.400 446.135 173.720 ;
        RECT 4.400 171.000 445.600 172.400 ;
        RECT 4.400 169.680 446.135 171.000 ;
        RECT 4.400 168.280 445.600 169.680 ;
        RECT 4.400 166.960 446.135 168.280 ;
        RECT 4.400 165.560 445.600 166.960 ;
        RECT 4.400 164.240 446.135 165.560 ;
        RECT 4.400 162.840 445.600 164.240 ;
        RECT 4.400 161.520 446.135 162.840 ;
        RECT 4.400 160.120 445.600 161.520 ;
        RECT 4.400 158.800 446.135 160.120 ;
        RECT 4.400 157.400 445.600 158.800 ;
        RECT 4.400 156.080 446.135 157.400 ;
        RECT 4.400 154.680 445.600 156.080 ;
        RECT 4.400 153.360 446.135 154.680 ;
        RECT 4.400 151.960 445.600 153.360 ;
        RECT 4.400 150.640 446.135 151.960 ;
        RECT 4.400 149.240 445.600 150.640 ;
        RECT 4.400 147.920 446.135 149.240 ;
        RECT 4.400 146.520 445.600 147.920 ;
        RECT 4.400 145.200 446.135 146.520 ;
        RECT 4.400 143.800 445.600 145.200 ;
        RECT 4.400 142.480 446.135 143.800 ;
        RECT 4.400 141.080 445.600 142.480 ;
        RECT 4.400 139.760 446.135 141.080 ;
        RECT 4.400 138.360 445.600 139.760 ;
        RECT 4.400 137.040 446.135 138.360 ;
        RECT 4.400 135.640 445.600 137.040 ;
        RECT 4.400 134.320 446.135 135.640 ;
        RECT 4.400 132.920 445.600 134.320 ;
        RECT 4.400 131.600 446.135 132.920 ;
        RECT 4.400 130.200 445.600 131.600 ;
        RECT 4.400 128.880 446.135 130.200 ;
        RECT 4.400 127.480 445.600 128.880 ;
        RECT 4.400 126.160 446.135 127.480 ;
        RECT 4.400 124.760 445.600 126.160 ;
        RECT 4.400 123.440 446.135 124.760 ;
        RECT 4.400 122.040 445.600 123.440 ;
        RECT 4.400 120.720 446.135 122.040 ;
        RECT 4.400 119.320 445.600 120.720 ;
        RECT 4.400 118.000 446.135 119.320 ;
        RECT 4.400 116.600 445.600 118.000 ;
        RECT 4.400 115.280 446.135 116.600 ;
        RECT 4.400 113.880 445.600 115.280 ;
        RECT 4.400 112.560 446.135 113.880 ;
        RECT 4.400 111.160 445.600 112.560 ;
        RECT 4.400 109.840 446.135 111.160 ;
        RECT 4.400 108.440 445.600 109.840 ;
        RECT 4.400 107.120 446.135 108.440 ;
        RECT 4.400 105.720 445.600 107.120 ;
        RECT 4.400 104.400 446.135 105.720 ;
        RECT 4.400 103.000 445.600 104.400 ;
        RECT 4.400 101.680 446.135 103.000 ;
        RECT 4.400 100.280 445.600 101.680 ;
        RECT 4.400 98.960 446.135 100.280 ;
        RECT 4.400 97.560 445.600 98.960 ;
        RECT 4.400 96.240 446.135 97.560 ;
        RECT 4.400 94.840 445.600 96.240 ;
        RECT 4.400 93.520 446.135 94.840 ;
        RECT 4.400 92.120 445.600 93.520 ;
        RECT 4.400 90.800 446.135 92.120 ;
        RECT 4.400 89.400 445.600 90.800 ;
        RECT 4.400 88.080 446.135 89.400 ;
        RECT 4.400 86.680 445.600 88.080 ;
        RECT 4.400 85.360 446.135 86.680 ;
        RECT 4.400 83.960 445.600 85.360 ;
        RECT 4.400 82.640 446.135 83.960 ;
        RECT 4.400 81.240 445.600 82.640 ;
        RECT 4.400 79.920 446.135 81.240 ;
        RECT 4.400 78.520 445.600 79.920 ;
        RECT 4.400 77.200 446.135 78.520 ;
        RECT 4.400 75.800 445.600 77.200 ;
        RECT 4.400 74.480 446.135 75.800 ;
        RECT 4.400 73.080 445.600 74.480 ;
        RECT 4.400 71.760 446.135 73.080 ;
        RECT 4.400 70.360 445.600 71.760 ;
        RECT 4.400 69.040 446.135 70.360 ;
        RECT 4.400 69.000 445.600 69.040 ;
        RECT 4.000 67.640 445.600 69.000 ;
        RECT 4.000 66.320 446.135 67.640 ;
        RECT 4.000 64.920 445.600 66.320 ;
        RECT 4.000 63.600 446.135 64.920 ;
        RECT 4.000 62.200 445.600 63.600 ;
        RECT 4.000 60.880 446.135 62.200 ;
        RECT 4.000 59.480 445.600 60.880 ;
        RECT 4.000 58.160 446.135 59.480 ;
        RECT 4.000 56.760 445.600 58.160 ;
        RECT 4.000 55.440 446.135 56.760 ;
        RECT 4.000 54.040 445.600 55.440 ;
        RECT 4.000 52.720 446.135 54.040 ;
        RECT 4.000 51.320 445.600 52.720 ;
        RECT 4.000 50.000 446.135 51.320 ;
        RECT 4.000 48.600 445.600 50.000 ;
        RECT 4.000 47.280 446.135 48.600 ;
        RECT 4.000 45.880 445.600 47.280 ;
        RECT 4.000 44.560 446.135 45.880 ;
        RECT 4.000 43.160 445.600 44.560 ;
        RECT 4.000 41.840 446.135 43.160 ;
        RECT 4.000 40.440 445.600 41.840 ;
        RECT 4.000 5.615 446.135 40.440 ;
      LAYER met4 ;
        RECT 2.150 438.560 444.065 449.305 ;
        RECT 2.150 10.240 20.640 438.560 ;
        RECT 23.040 10.240 97.440 438.560 ;
        RECT 99.840 10.240 174.240 438.560 ;
        RECT 176.640 10.240 251.040 438.560 ;
        RECT 253.440 10.240 327.840 438.560 ;
        RECT 330.240 10.240 404.640 438.560 ;
        RECT 407.040 10.240 444.065 438.560 ;
        RECT 2.150 5.615 444.065 10.240 ;
  END
END busarb_2_2
END LIBRARY

