* NGSPICE file created from mac_piped.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

.subckt mac_piped a_i[0] a_i[10] a_i[11] a_i[12] a_i[13] a_i[14] a_i[15] a_i[16] a_i[17]
+ a_i[18] a_i[19] a_i[1] a_i[20] a_i[21] a_i[22] a_i[23] a_i[24] a_i[25] a_i[26] a_i[27]
+ a_i[28] a_i[29] a_i[2] a_i[30] a_i[31] a_i[3] a_i[4] a_i[5] a_i[6] a_i[7] a_i[8]
+ a_i[9] b_i[0] b_i[10] b_i[11] b_i[12] b_i[13] b_i[14] b_i[15] b_i[16] b_i[17] b_i[18]
+ b_i[19] b_i[1] b_i[20] b_i[21] b_i[22] b_i[23] b_i[24] b_i[25] b_i[26] b_i[27] b_i[28]
+ b_i[29] b_i[2] b_i[30] b_i[31] b_i[3] b_i[4] b_i[5] b_i[6] b_i[7] b_i[8] b_i[9]
+ clk nrst vccd1 vssd1 y_o[0] y_o[10] y_o[11] y_o[12] y_o[13] y_o[14] y_o[15] y_o[16]
+ y_o[17] y_o[18] y_o[19] y_o[1] y_o[20] y_o[21] y_o[22] y_o[23] y_o[24] y_o[25] y_o[26]
+ y_o[27] y_o[28] y_o[29] y_o[2] y_o[30] y_o[31] y_o[3] y_o[4] y_o[5] y_o[6] y_o[7]
+ y_o[8] y_o[9]
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05903_ _05903_/A _05903_/B _05903_/C vssd1 vssd1 vccd1 vccd1 _05906_/B sky130_fd_sc_hd__nand3_1
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__nand2_1
X_06883_ _06883_/A _06884_/A vssd1 vssd1 vccd1 vccd1 _06886_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08622_ _08624_/B _08886_/C vssd1 vssd1 vccd1 vccd1 _08623_/A sky130_fd_sc_hd__nand2_1
X_05834_ input5/X _08688_/A vssd1 vssd1 vccd1 vccd1 _05948_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08553_ _08557_/C vssd1 vssd1 vccd1 vccd1 _08553_/Y sky130_fd_sc_hd__inv_2
X_05765_ _05766_/B _05765_/B vssd1 vssd1 vccd1 vccd1 _05787_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08484_ _08737_/B _08485_/C _08485_/B vssd1 vssd1 vccd1 vccd1 _08490_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_9_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07504_ _07540_/C _07571_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07539_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_64_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05696_ _06175_/B _05696_/B vssd1 vssd1 vccd1 vccd1 _05729_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07435_ _09854_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _07440_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07366_ _07366_/A _07366_/B vssd1 vssd1 vccd1 vccd1 _07366_/Y sky130_fd_sc_hd__nor2_1
X_09105_ _09108_/B _09406_/B vssd1 vssd1 vccd1 vccd1 _09107_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06317_ _06330_/B _05954_/Y _05955_/Y vssd1 vssd1 vccd1 vccd1 _06318_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07297_ _09951_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _07298_/A sky130_fd_sc_hd__nand2_1
X_09036_ _09083_/A _10084_/D _09035_/C vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06248_ _09720_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _06696_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09211__B2 _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06179_ _06179_/A _06179_/B _06179_/C vssd1 vssd1 vccd1 vccd1 _06180_/B sky130_fd_sc_hd__nand3_1
X_09938_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06411__B _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09869_ _09869_/A _09869_/B _10100_/B vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09722__B _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06139__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10009_ _10010_/A _10010_/C _10010_/B vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07433__A _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08248__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05550_ _05550_/A _05551_/A vssd1 vssd1 vccd1 vccd1 _05562_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05481_ input38/X vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ _07220_/A _07221_/A vssd1 vssd1 vccd1 vccd1 _07223_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07151_ _07151_/A _07151_/B vssd1 vssd1 vccd1 vccd1 _07706_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06102_ _06402_/A _06404_/A _06103_/B vssd1 vssd1 vccd1 vccd1 _06183_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_14_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07082_ _07082_/A _07082_/B _07082_/C vssd1 vssd1 vccd1 vccd1 _07083_/B sky130_fd_sc_hd__nand3_1
X_06033_ _10026_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _06034_/B sky130_fd_sc_hd__nand2_1
X_07984_ _07984_/A _08091_/B vssd1 vssd1 vccd1 vccd1 _08087_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09723_ input46/X _10051_/B _10051_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _09723_/X
+ sky130_fd_sc_hd__a22o_1
X_06935_ _07090_/A _07090_/C vssd1 vssd1 vccd1 vccd1 _06940_/A sky130_fd_sc_hd__nand2_1
X_09654_ _09654_/A _09655_/A vssd1 vssd1 vccd1 vccd1 _09661_/B sky130_fd_sc_hd__nand2_1
X_06866_ _07024_/B _07024_/C vssd1 vssd1 vccd1 vccd1 _07023_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08605_ _08603_/Y _08381_/B _08604_/Y vssd1 vssd1 vccd1 vccd1 _08628_/A sky130_fd_sc_hd__a21oi_2
X_05817_ _05817_/A vssd1 vssd1 vccd1 vccd1 _05824_/B sky130_fd_sc_hd__inv_2
X_09585_ _09585_/A _09586_/A vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__nand2_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06797_ _06797_/A _06797_/B vssd1 vssd1 vccd1 vccd1 _06843_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08536_ _08540_/A _08540_/B vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__nand2_1
X_05748_ _05748_/A _05748_/B vssd1 vssd1 vccd1 vccd1 _05886_/C sky130_fd_sc_hd__nand2_1
X_08467_ _08467_/A _08467_/B _08467_/C vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07997__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05679_ _05448_/C _05448_/B _05678_/Y vssd1 vssd1 vccd1 vccd1 _06107_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08398_ _08620_/B _08398_/B vssd1 vssd1 vccd1 vccd1 _08401_/B sky130_fd_sc_hd__nand2_1
X_07418_ _07418_/A _07418_/B _07418_/C vssd1 vssd1 vccd1 vccd1 _07419_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07349_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07352_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ _10360_/A hold60/X vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__nand2_1
X_09019_ _09046_/B _09046_/C vssd1 vssd1 vccd1 vccd1 _09045_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10291_ _10495_/Q hold113/X vssd1 vssd1 vccd1 vccd1 hold114/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09499__B2 _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__A1 _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10489_ _10495_/CLK hold42/X fanout99/X vssd1 vssd1 vccd1 vccd1 _10489_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07428__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06720_ _06720_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _06982_/B sky130_fd_sc_hd__or2b_1
X_06651_ _06651_/A _06651_/B vssd1 vssd1 vccd1 vccd1 _06654_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07163__A _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05602_ input38/X _08810_/B vssd1 vssd1 vccd1 vccd1 _05604_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _09608_/A _09370_/B vssd1 vssd1 vccd1 vccd1 _09372_/A sky130_fd_sc_hd__nand2_1
X_06582_ _06582_/A _06582_/B vssd1 vssd1 vccd1 vccd1 _06590_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08321_ _08386_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__nand2_1
X_05533_ _05533_/A vssd1 vssd1 vccd1 vccd1 _05534_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08706__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ _08253_/B _08253_/A vssd1 vssd1 vccd1 vccd1 _08464_/A sky130_fd_sc_hd__or2_1
X_05464_ _05464_/A _05464_/B _05464_/C vssd1 vssd1 vccd1 vccd1 _05826_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ _07203_/A _07203_/B vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05411__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _08140_/Y _08144_/Y _08182_/X vssd1 vssd1 vccd1 vccd1 _08184_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06226__B _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05395_ _05395_/A _05395_/B _05398_/A vssd1 vssd1 vccd1 vccd1 _05400_/A sky130_fd_sc_hd__nand3_1
XANTENNA__10024__A2 _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07134_ _07659_/A _07658_/A vssd1 vssd1 vccd1 vccd1 _07134_/Y sky130_fd_sc_hd__nor2_1
X_07065_ _07079_/B _07080_/B _07080_/A vssd1 vssd1 vccd1 vccd1 _07092_/B sky130_fd_sc_hd__nand3_1
X_06016_ _06016_/A _06463_/A _06016_/C vssd1 vssd1 vccd1 vccd1 _06408_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07967_ _07989_/A _07989_/C _07989_/B vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__a21boi_2
X_09706_ _09701_/Y _09706_/B vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__nand2b_1
X_06918_ _10083_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _07110_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07073__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _07898_/A _07898_/B _07898_/C vssd1 vssd1 vccd1 vccd1 _07907_/B sky130_fd_sc_hd__nand3_1
X_09637_ _09637_/A _09637_/B vssd1 vssd1 vccd1 vccd1 _09917_/A sky130_fd_sc_hd__nand2_1
X_06849_ _06849_/A _06849_/B vssd1 vssd1 vccd1 vccd1 _07008_/B sky130_fd_sc_hd__nand2_1
X_09568_ _09568_/A _09568_/B _09568_/C vssd1 vssd1 vccd1 vccd1 _09569_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08519_ _08854_/A _08672_/A _08520_/A vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _09963_/A _09960_/B _09962_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _09692_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05321__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10412_ _10413_/B _10413_/A vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__or2_1
X_10343_ hold66/X _10344_/A vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10274_ hold106/X vssd1 vssd1 vccd1 vccd1 _10492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09463__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05231__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08870_ _08870_/A vssd1 vssd1 vccd1 vccd1 _08870_/Y sky130_fd_sc_hd__inv_2
X_07821_ _07821_/A _07821_/B vssd1 vssd1 vccd1 vccd1 _07822_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07752_ _07752_/A _07753_/A vssd1 vssd1 vccd1 vccd1 _07755_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07683_ _07683_/A _07683_/B vssd1 vssd1 vccd1 vccd1 _07692_/B sky130_fd_sc_hd__nand2_1
X_06703_ _06703_/A _06703_/B _06703_/C vssd1 vssd1 vccd1 vccd1 _06946_/B sky130_fd_sc_hd__nand3_1
X_09422_ _09427_/A _09669_/A vssd1 vssd1 vccd1 vccd1 _09426_/A sky130_fd_sc_hd__nand2_1
X_06634_ _06634_/A _06634_/B vssd1 vssd1 vccd1 vccd1 _08656_/A sky130_fd_sc_hd__nand2_1
X_09353_ _09353_/A _09353_/B vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06565_ _06565_/A _06565_/B vssd1 vssd1 vccd1 vccd1 _06566_/B sky130_fd_sc_hd__nand2_1
X_08304_ _08511_/A _08304_/B _08582_/A vssd1 vssd1 vccd1 vccd1 _08308_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09284_ _09448_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _09286_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06496_ _06502_/B vssd1 vssd1 vccd1 vccd1 _06499_/B sky130_fd_sc_hd__inv_2
X_05516_ _05516_/A _05998_/A vssd1 vssd1 vccd1 vccd1 _05518_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08236_/B sky130_fd_sc_hd__nand2_1
X_05447_ _05447_/A vssd1 vssd1 vccd1 vccd1 _05448_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09548__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ _10385_/B _08196_/C vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__nor2_1
X_05378_ _05397_/A _05397_/C vssd1 vssd1 vccd1 vccd1 _05405_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08452__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07117_ _07357_/B _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07363_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09267__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08097_ _10111_/B _09986_/A vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__nand2_1
X_07048_ _07051_/B _07060_/A vssd1 vssd1 vccd1 vccd1 _07050_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07068__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08999_ _10027_/A _10044_/D _08999_/C vssd1 vssd1 vccd1 vccd1 _09234_/A sky130_fd_sc_hd__nor3_1
XANTENNA__05316__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10326_ _10326_/A hold15/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__xor2_1
XFILLER_0_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _10491_/Q hold102/X vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__nor2_1
X_10188_ _10482_/Q hold17/X vssd1 vssd1 vccd1 vccd1 _10190_/A sky130_fd_sc_hd__or2_1
XANTENNA__07425__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06350_ _06756_/B _06755_/A vssd1 vssd1 vccd1 vccd1 _06350_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05301_ _05303_/B vssd1 vssd1 vccd1 vccd1 _05302_/B sky130_fd_sc_hd__inv_2
X_06281_ _06296_/C _06299_/A vssd1 vssd1 vccd1 vccd1 _06291_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08020_ _08020_/A _08020_/B vssd1 vssd1 vccd1 vccd1 _08020_/Y sky130_fd_sc_hd__nor2_1
X_05232_ _05311_/A vssd1 vssd1 vccd1 vccd1 _05243_/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08272__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09971_ _09971_/A _09971_/B vssd1 vssd1 vccd1 vccd1 _09971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10026__B _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _09291_/A sky130_fd_sc_hd__nand2_1
X_08853_ _08854_/B _08854_/A vssd1 vssd1 vccd1 vccd1 _08853_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08784_ _10026_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _08785_/B sky130_fd_sc_hd__nand2_1
X_05996_ _05996_/A _05996_/B _05996_/C vssd1 vssd1 vccd1 vccd1 _06018_/C sky130_fd_sc_hd__nand3_2
X_07804_ _07803_/B _07804_/B _07804_/C vssd1 vssd1 vccd1 vccd1 _07893_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07735_ _07744_/B _07744_/C vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _09408_/B _09408_/C vssd1 vssd1 vccd1 vccd1 _09407_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__nand2_1
X_06617_ _06617_/A _08388_/A _06617_/C vssd1 vssd1 vccd1 vccd1 _06618_/B sky130_fd_sc_hd__nand3_1
X_07597_ _07719_/B _07717_/A vssd1 vssd1 vccd1 vccd1 _07597_/Y sky130_fd_sc_hd__nand2_1
X_09336_ _09339_/B _09339_/C vssd1 vssd1 vccd1 vccd1 _09338_/A sky130_fd_sc_hd__nand2_1
X_06548_ _06549_/A _06549_/B vssd1 vssd1 vccd1 vccd1 _08322_/B sky130_fd_sc_hd__or2_1
XANTENNA__07070__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _09980_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08218_ _08219_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08221_/A sky130_fd_sc_hd__nor2_1
X_06479_ _09951_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _06481_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ _10043_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _09204_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _08151_/B _08151_/A vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ input56/X _10111_/B vssd1 vssd1 vccd1 vccd1 _10120_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10042_ _10060_/A _10060_/C vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__nand2_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09188__A _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10309_ _10497_/Q hold117/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__nand2_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05850_ _05851_/B _05850_/B _05850_/C vssd1 vssd1 vccd1 vccd1 _06366_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07520_ _07520_/A _07520_/B vssd1 vssd1 vccd1 vccd1 _07523_/B sky130_fd_sc_hd__nand2_1
X_05781_ _05781_/A _05781_/B _05781_/C vssd1 vssd1 vccd1 vccd1 _05782_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07451_ _07451_/A _07451_/B _07451_/C vssd1 vssd1 vccd1 vccd1 _07453_/B sky130_fd_sc_hd__nand3_1
X_06402_ _06402_/A _06402_/B vssd1 vssd1 vccd1 vccd1 _06402_/Y sky130_fd_sc_hd__nor2_1
X_07382_ _07382_/A _07382_/B vssd1 vssd1 vccd1 vccd1 _07525_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09121_ _09127_/B vssd1 vssd1 vccd1 vccd1 _09125_/B sky130_fd_sc_hd__inv_2
X_06333_ _06333_/A _06333_/B vssd1 vssd1 vccd1 vccd1 _06335_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09052_ _09399_/B _09052_/B vssd1 vssd1 vccd1 vccd1 _09060_/A sky130_fd_sc_hd__nand2_1
X_06264_ _06264_/A _06264_/B _06264_/C vssd1 vssd1 vccd1 vccd1 _06658_/B sky130_fd_sc_hd__nand3_1
X_08003_ _08003_/A _08003_/B vssd1 vssd1 vccd1 vccd1 _08010_/B sky130_fd_sc_hd__xnor2_1
X_05215_ _05215_/A _05215_/B _05217_/A vssd1 vssd1 vccd1 vccd1 _05338_/B sky130_fd_sc_hd__nand3_1
X_06195_ _06399_/B _06399_/A vssd1 vssd1 vccd1 vccd1 _06196_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06234__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _09485_/C _09775_/B _09804_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09955_/B
+ sky130_fd_sc_hd__a22o_1
X_09885_ _09885_/A _09885_/B _10140_/A vssd1 vssd1 vccd1 vccd1 _09908_/C sky130_fd_sc_hd__nand3_1
X_08905_ _08905_/A vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__inv_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06250__A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08836_ _08836_/A _08836_/B _08836_/C vssd1 vssd1 vccd1 vccd1 _08843_/C sky130_fd_sc_hd__nand3_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _08773_/B vssd1 vssd1 vccd1 vccd1 _08771_/B sky130_fd_sc_hd__inv_2
X_05979_ _05979_/A _05979_/B vssd1 vssd1 vccd1 vccd1 _05979_/Y sky130_fd_sc_hd__nor2_1
X_08698_ _08697_/B _08927_/B _08698_/C vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__nand3b_1
X_07718_ _07574_/Y _07730_/B _07595_/Y vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07649_ _07649_/A _07913_/B vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06409__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ _09319_/A _09484_/A vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput75 _10498_/Q vssd1 vssd1 vccd1 vccd1 y_o[18] sky130_fd_sc_hd__buf_12
Xoutput86 hold69/A vssd1 vssd1 vccd1 vccd1 y_o[28] sky130_fd_sc_hd__buf_12
Xoutput97 _10489_/Q vssd1 vssd1 vccd1 vccd1 y_o[9] sky130_fd_sc_hd__buf_12
XANTENNA__07256__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10025_ _10025_/A vssd1 vssd1 vccd1 vccd1 _10032_/B sky130_fd_sc_hd__inv_2
XFILLER_0_98_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06054__B _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08550__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06070__A _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07166__A _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _06951_/A _06951_/B vssd1 vssd1 vccd1 vccd1 _06952_/A sky130_fd_sc_hd__nand2_1
X_09670_ _09672_/A vssd1 vssd1 vccd1 vccd1 _09671_/B sky130_fd_sc_hd__inv_2
X_05902_ _05902_/A _05902_/B vssd1 vssd1 vccd1 vccd1 _05906_/A sky130_fd_sc_hd__nand2_1
X_08621_ _08886_/B _08621_/B _08621_/C vssd1 vssd1 vccd1 vccd1 _08886_/C sky130_fd_sc_hd__nand3_2
X_06882_ _09022_/C _07960_/B vssd1 vssd1 vccd1 vccd1 _06884_/A sky130_fd_sc_hd__nand2_1
X_05833_ _05949_/C vssd1 vssd1 vccd1 vccd1 _05918_/B sky130_fd_sc_hd__inv_2
X_08552_ _10044_/A _10084_/B _08551_/C vssd1 vssd1 vccd1 vccd1 _08557_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05764_ _09528_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _05765_/B sky130_fd_sc_hd__nand2_1
X_08483_ _08483_/A vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07503_ _07503_/A _07503_/B _07503_/C vssd1 vssd1 vccd1 vccd1 _07571_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05695_ _05748_/B _05693_/Y _05749_/B vssd1 vssd1 vccd1 vccd1 _05696_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07434_ _07440_/A vssd1 vssd1 vccd1 vccd1 _07437_/A sky130_fd_sc_hd__inv_2
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07365_ _07366_/B _07366_/A vssd1 vssd1 vccd1 vccd1 _07365_/Y sky130_fd_sc_hd__nand2_1
X_09104_ _09104_/A _09104_/B _09385_/A vssd1 vssd1 vccd1 vccd1 _09406_/B sky130_fd_sc_hd__nand3_1
X_06316_ _06316_/A _06316_/B _06316_/C vssd1 vssd1 vccd1 vccd1 _06321_/A sky130_fd_sc_hd__nand3_1
X_07296_ _07299_/A _07299_/B vssd1 vssd1 vccd1 vccd1 _07323_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ _09083_/A _10084_/D _09035_/C vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__nor3_1
X_06247_ _09560_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _06695_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09211__A2 _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06178_ _06178_/A vssd1 vssd1 vccd1 vccd1 _06179_/C sky130_fd_sc_hd__inv_2
XFILLER_0_40_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09937_ _09939_/B _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _10171_/B sky130_fd_sc_hd__nand3b_4
XANTENNA__06411__C _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ _10091_/A _09868_/B _09868_/C vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__nand3_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09799_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09722__C _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ _08819_/A vssd1 vssd1 vccd1 vccd1 _08832_/A sky130_fd_sc_hd__inv_2
XFILLER_0_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10045__B1 _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__A1 _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06155__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10511__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _10008_/A _10008_/B vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07433__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05480_ _05486_/C vssd1 vssd1 vccd1 vccd1 _05480_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07150_ _07154_/B _07150_/B vssd1 vssd1 vccd1 vccd1 _07151_/A sky130_fd_sc_hd__nand2_1
X_06101_ _06101_/A _06101_/B _06101_/C vssd1 vssd1 vccd1 vccd1 _06103_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_14_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07081_ _07081_/A vssd1 vssd1 vccd1 vccd1 _07082_/C sky130_fd_sc_hd__inv_2
X_06032_ _07216_/B vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ input46/X _10051_/A _10051_/B _10050_/B vssd1 vssd1 vccd1 vccd1 _09724_/A
+ sky130_fd_sc_hd__and4_1
X_07983_ _07983_/A _08040_/B _08040_/A vssd1 vssd1 vccd1 vccd1 _08091_/B sky130_fd_sc_hd__nand3_2
X_06934_ _06934_/A _06934_/B _06934_/C vssd1 vssd1 vccd1 vccd1 _07090_/C sky130_fd_sc_hd__nand3_1
X_09653_ _09932_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__nand2_1
X_06865_ _06865_/A _06865_/B _06865_/C vssd1 vssd1 vccd1 vccd1 _07024_/C sky130_fd_sc_hd__nand3_1
X_09584_ _09911_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10050__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _08604_/A _08604_/B vssd1 vssd1 vccd1 vccd1 _08604_/Y sky130_fd_sc_hd__nor2_1
X_05816_ _06213_/B _06216_/B vssd1 vssd1 vccd1 vccd1 _05817_/A sky130_fd_sc_hd__nor2_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _08800_/A _08802_/A _08800_/B vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__nand3_1
X_06796_ _06796_/A _06796_/B vssd1 vssd1 vccd1 vccd1 _06797_/B sky130_fd_sc_hd__nand2_1
X_05747_ _05749_/A _05749_/B vssd1 vssd1 vccd1 vccd1 _05748_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08455__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ _08467_/A _08467_/C _08467_/B vssd1 vssd1 vccd1 vccd1 _08468_/A sky130_fd_sc_hd__a21o_1
X_05678_ _05678_/A _05678_/B vssd1 vssd1 vccd1 vccd1 _05678_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08397_ _08397_/A _08397_/B vssd1 vssd1 vccd1 vccd1 _08398_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07417_ _07417_/A _07417_/B _07417_/C vssd1 vssd1 vccd1 vccd1 _07418_/B sky130_fd_sc_hd__nand3_1
X_07348_ _07350_/A _07350_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07279_ _07315_/B _07283_/B vssd1 vssd1 vccd1 vccd1 _07281_/B sky130_fd_sc_hd__nand2_1
X_09018_ _09018_/A _09217_/A _09018_/C vssd1 vssd1 vccd1 vccd1 _09046_/C sky130_fd_sc_hd__nand3_1
X_10290_ _10495_/Q hold113/X vssd1 vssd1 vccd1 vccd1 _10290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09499__A2 _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08349__B _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10488_ _10494_/CLK _10488_/D fanout99/X vssd1 vssd1 vccd1 vccd1 _10488_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07709__A _07709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06650_ _06831_/B _06650_/B vssd1 vssd1 vccd1 vccd1 _06651_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07163__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05601_ _05605_/A _05605_/C vssd1 vssd1 vccd1 vccd1 _05603_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06581_ _06583_/B vssd1 vssd1 vccd1 vccd1 _06582_/B sky130_fd_sc_hd__inv_2
X_08320_ _08521_/A _08320_/B _08597_/A vssd1 vssd1 vccd1 vccd1 _08386_/B sky130_fd_sc_hd__nand3_1
X_05532_ _05532_/A _05533_/A vssd1 vssd1 vccd1 vccd1 _05535_/A sky130_fd_sc_hd__nand2_1
X_08251_ _08464_/B _08251_/B vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__nand2_1
X_05463_ _05462_/B _05463_/B vssd1 vssd1 vccd1 vccd1 _05464_/B sky130_fd_sc_hd__nand2b_1
X_07202_ _07202_/A vssd1 vssd1 vccd1 vccd1 _07203_/B sky130_fd_sc_hd__inv_2
XANTENNA__05411__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _09890_/D _09986_/A _09392_/D _09751_/A _08142_/C vssd1 vssd1 vccd1 vccd1
+ _08182_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05394_ _05920_/B _05829_/A vssd1 vssd1 vccd1 vccd1 _05398_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10024__A3 _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07133_ _07133_/A _07133_/B vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__nor2_2
X_07064_ _07064_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _07080_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06015_ _06019_/C vssd1 vssd1 vccd1 vccd1 _06016_/C sky130_fd_sc_hd__inv_2
XFILLER_0_100_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _07966_/A _07966_/B _07966_/C vssd1 vssd1 vccd1 vccd1 _07989_/B sky130_fd_sc_hd__nand3_1
X_09705_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09706_/B sky130_fd_sc_hd__nor2_1
X_06917_ _09854_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _07111_/B sky130_fd_sc_hd__nand2_2
X_09636_ _09638_/C vssd1 vssd1 vccd1 vccd1 _09637_/B sky130_fd_sc_hd__inv_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07073__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ _07606_/Y _07803_/B _07607_/Y vssd1 vssd1 vccd1 vccd1 _07898_/A sky130_fd_sc_hd__a21o_1
X_06848_ _06850_/A _06850_/B vssd1 vssd1 vccd1 vccd1 _06849_/A sky130_fd_sc_hd__nand2_1
X_09567_ _09567_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09569_/A sky130_fd_sc_hd__nand2_1
X_06779_ _06847_/B _06845_/A vssd1 vssd1 vccd1 vccd1 _06779_/Y sky130_fd_sc_hd__nand2_1
X_09498_ _09498_/A vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__inv_2
X_08518_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08520_/A sky130_fd_sc_hd__nand2_1
X_08449_ _08449_/A _08449_/B _08449_/C vssd1 vssd1 vccd1 vccd1 _08471_/C sky130_fd_sc_hd__nand3_2
XANTENNA__05602__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10411_ _10407_/B _10409_/A _10407_/A _07678_/Y vssd1 vssd1 vccd1 vccd1 _10413_/A
+ sky130_fd_sc_hd__a31o_1
X_10342_ hold110/A _10333_/B _10340_/A _10341_/Y vssd1 vssd1 vccd1 vccd1 _10344_/A
+ sky130_fd_sc_hd__a31o_1
X_10273_ hold105/X _10278_/A vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__and2_1
XANTENNA__09463__B input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05512__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05231__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _07921_/B _07921_/C vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07751_ _09361_/D _07960_/B vssd1 vssd1 vccd1 vccd1 _07753_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06702_ _06702_/A _06702_/B vssd1 vssd1 vccd1 vccd1 _06946_/A sky130_fd_sc_hd__nand2_1
X_07682_ _07132_/Y _07666_/B _07134_/Y vssd1 vssd1 vccd1 vccd1 _07683_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09421_ _09421_/A _09669_/B _09421_/C vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__nand3_1
X_06633_ _06633_/A _09188_/A _06633_/C vssd1 vssd1 vccd1 vccd1 _06640_/A sky130_fd_sc_hd__nand3_2
X_09352_ _09352_/A _09352_/B vssd1 vssd1 vccd1 vccd1 _09353_/B sky130_fd_sc_hd__and2_1
X_06564_ _06564_/A _06564_/B vssd1 vssd1 vccd1 vccd1 _06565_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08303_ _08582_/B _08303_/B vssd1 vssd1 vccd1 vccd1 _08308_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05515_ _05515_/A _05515_/B _05515_/C vssd1 vssd1 vccd1 vccd1 _05539_/C sky130_fd_sc_hd__nand3_1
XANTENNA__10493__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05422__A _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ _10000_/A _09775_/B _09999_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09284_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06495_ _06495_/A _08356_/A vssd1 vssd1 vccd1 vccd1 _06502_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_51_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08234_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08236_/A sky130_fd_sc_hd__or2_1
X_05446_ _05446_/A _05447_/A vssd1 vssd1 vccd1 vccd1 _05449_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08165_ _08195_/B _08194_/A _08194_/B vssd1 vssd1 vccd1 vccd1 _08196_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05377_ _05377_/A _05377_/B vssd1 vssd1 vccd1 vccd1 _05397_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08452__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07116_ _07116_/A _07116_/B vssd1 vssd1 vccd1 vccd1 _07356_/B sky130_fd_sc_hd__nand2_1
X_08096_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08112_/B sky130_fd_sc_hd__xor2_1
X_07047_ _07060_/B vssd1 vssd1 vccd1 vccd1 _07051_/B sky130_fd_sc_hd__inv_2
XANTENNA__07068__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08998_ _09685_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _08999_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07949_ _07950_/A _07950_/B vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05316__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ _09616_/B _09619_/B _09619_/C vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_85_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06428__A _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ _10325_/A hold14/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__nand2_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ hold101/X vssd1 vssd1 vccd1 vccd1 _10490_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__05820__B1 _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05507__A _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ hold56/X vssd1 vssd1 vccd1 vccd1 _10481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05300_ input6/X _08248_/B vssd1 vssd1 vccd1 vccd1 _05303_/B sky130_fd_sc_hd__nand2_1
X_06280_ _06280_/A _06280_/B vssd1 vssd1 vccd1 vccd1 _06296_/C sky130_fd_sc_hd__nand2_1
X_05231_ _09496_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _05311_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08272__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06073__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09970_ _09949_/Y _09950_/Y _09969_/Y vssd1 vssd1 vccd1 vccd1 _09977_/B sky130_fd_sc_hd__o21ai_1
X_08921_ _08922_/B _08922_/A vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__or2_1
X_08852_ _09141_/B _09141_/C vssd1 vssd1 vccd1 vccd1 _09140_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05417__A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _07803_/A _07803_/B vssd1 vssd1 vccd1 vccd1 _07893_/A sky130_fd_sc_hd__nand2_1
X_08783_ _08995_/B _08786_/C vssd1 vssd1 vccd1 vccd1 _08785_/A sky130_fd_sc_hd__nand2_1
X_05995_ _05995_/A vssd1 vssd1 vccd1 vccd1 _05996_/B sky130_fd_sc_hd__inv_2
X_07734_ _07734_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08728__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07695_/B sky130_fd_sc_hd__nand2_1
X_09404_ _09648_/A _09404_/B _09663_/A vssd1 vssd1 vccd1 vccd1 _09408_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06616_ _06616_/A _06616_/B vssd1 vssd1 vccd1 vccd1 _06618_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06248__A _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07596_ _07574_/Y _07730_/B _07595_/Y vssd1 vssd1 vccd1 vccd1 _07717_/A sky130_fd_sc_hd__a21oi_1
X_09335_ _09335_/A _09335_/B _09575_/A vssd1 vssd1 vccd1 vccd1 _09339_/C sky130_fd_sc_hd__nand3_1
X_06547_ _09199_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _06549_/B sky130_fd_sc_hd__nand2_1
X_09266_ _09275_/B _09473_/B vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__nand2_1
X_06478_ _08281_/B _06482_/B vssd1 vssd1 vccd1 vccd1 _06480_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08217_ _08422_/A input17/X vssd1 vssd1 vccd1 vccd1 _08219_/B sky130_fd_sc_hd__nand2_1
X_05429_ _09951_/A _09022_/D vssd1 vssd1 vccd1 vccd1 _05464_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09197_ _09023_/X _09026_/B _09024_/A vssd1 vssd1 vccd1 vccd1 _09594_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08148_ _08148_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__nand2_1
X_08079_ _08079_/A _08079_/B _08079_/C vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__nand3_1
X_10110_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10110_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout98_A fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _10041_/A _10041_/B _10041_/C vssd1 vssd1 vccd1 vccd1 _10060_/C sky130_fd_sc_hd__nand3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10308_ _10497_/Q hold117/X vssd1 vssd1 vccd1 vccd1 _10308_/Y sky130_fd_sc_hd__nor2_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ hold92/X _10244_/A vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__and2_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05780_ _05780_/A _05780_/B vssd1 vssd1 vccd1 vccd1 _06187_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06068__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07450_ _07450_/A _07450_/B vssd1 vssd1 vccd1 vccd1 _07453_/A sky130_fd_sc_hd__nand2_1
X_06401_ _06402_/B _06402_/A vssd1 vssd1 vccd1 vccd1 _06401_/Y sky130_fd_sc_hd__nand2_1
X_07381_ _07410_/A _07528_/B vssd1 vssd1 vccd1 vccd1 _07526_/B sky130_fd_sc_hd__nor2b_1
X_09120_ _09120_/A _09418_/A vssd1 vssd1 vccd1 vccd1 _09127_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06332_ _06736_/B _06736_/C vssd1 vssd1 vccd1 vccd1 _06735_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09051_ _09399_/A vssd1 vssd1 vccd1 vccd1 _09052_/B sky130_fd_sc_hd__inv_2
X_08002_ _08002_/A vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__inv_2
X_06263_ _06263_/A _06263_/B vssd1 vssd1 vccd1 vccd1 _06658_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05214_ _09960_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _05217_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06194_ _05976_/Y _05784_/B _05977_/Y vssd1 vssd1 vccd1 vccd1 _06399_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout100_A fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ _09953_/A _09953_/B _09953_/C _09775_/B vssd1 vssd1 vccd1 vccd1 _09955_/A
+ sky130_fd_sc_hd__or4b_1
X_09884_ _10140_/B _09884_/B vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__nand2_1
X_08904_ _09751_/A _09762_/B _08904_/C vssd1 vssd1 vccd1 vccd1 _08905_/A sky130_fd_sc_hd__nor3_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06250__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08835_ _08835_/A _08835_/B vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__nand2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08766_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08773_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05978_ _05976_/Y _05784_/B _05977_/Y vssd1 vssd1 vccd1 vccd1 _06197_/B sky130_fd_sc_hd__a21o_1
X_07717_ _07717_/A _07717_/B _07717_/C vssd1 vssd1 vccd1 vccd1 _07722_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08697_ _08697_/A _08697_/B vssd1 vssd1 vccd1 vccd1 _08703_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07648_ _07697_/A _07651_/C vssd1 vssd1 vccd1 vccd1 _07649_/A sky130_fd_sc_hd__nand2_1
X_07579_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07592_/B sky130_fd_sc_hd__nand2_1
X_09318_ _09318_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09289__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _09252_/B _09252_/C vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput76 _10499_/Q vssd1 vssd1 vccd1 vccd1 y_o[19] sky130_fd_sc_hd__buf_12
XANTENNA__06441__A _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 hold1/A vssd1 vssd1 vccd1 vccd1 y_o[29] sky130_fd_sc_hd__buf_12
XANTENNA__07256__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10024_ _09819_/B _09960_/A _09816_/B _09817_/X vssd1 vssd1 vccd1 vccd1 _10025_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_98_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09199__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08550__B _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06070__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07166__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ _06952_/B _06951_/A _06951_/B vssd1 vssd1 vccd1 vccd1 _06953_/A sky130_fd_sc_hd__nand3b_1
X_06881_ _06885_/A _06885_/C vssd1 vssd1 vccd1 vccd1 _06883_/A sky130_fd_sc_hd__nand2_1
X_05901_ _05903_/A vssd1 vssd1 vccd1 vccd1 _05902_/B sky130_fd_sc_hd__inv_2
XANTENNA__08731__A2 _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _08620_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__nand2_1
X_05832_ _09533_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _05949_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _10044_/A _10084_/B _08551_/C vssd1 vssd1 vccd1 vccd1 _08551_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05763_ _09685_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _05766_/B sky130_fd_sc_hd__nand2_1
X_08482_ _09951_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__nand2_1
X_05694_ _05694_/A _05694_/B _05694_/C vssd1 vssd1 vccd1 vccd1 _05749_/B sky130_fd_sc_hd__nand3_1
X_07502_ _07556_/C _07496_/Y _07556_/A vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07433_ _09601_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _07440_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09103_ _08882_/C _08882_/B _08878_/Y vssd1 vssd1 vccd1 vccd1 _09104_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06526__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07364_ _07370_/A _07370_/B vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06315_ _06654_/A vssd1 vssd1 vccd1 vccd1 _06653_/B sky130_fd_sc_hd__inv_2
X_07295_ _09601_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _07299_/B sky130_fd_sc_hd__nand2_1
X_09034_ _10051_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _09035_/C sky130_fd_sc_hd__nand2_1
X_06246_ _06376_/A _06377_/A vssd1 vssd1 vccd1 vccd1 _06246_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06177_ _06177_/A _06178_/A vssd1 vssd1 vccd1 vccd1 _06180_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ _09936_/A _09936_/B _09936_/C vssd1 vssd1 vccd1 vccd1 _09938_/B sky130_fd_sc_hd__nand3_2
X_09867_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__nand2_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _09798_/A _09799_/B _09799_/A vssd1 vssd1 vccd1 vccd1 _09835_/B sky130_fd_sc_hd__nand3_2
XANTENNA__09722__D _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ _08820_/B _08820_/A vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10463__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _08750_/B _08750_/A vssd1 vssd1 vccd1 vccd1 _08751_/A sky130_fd_sc_hd__or2_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08916__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10045__A1 _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__B2 _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06155__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06171__A _06173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10007_ _10007_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _10008_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08098__A _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06346__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06100_ _06594_/A _06100_/B _06100_/C vssd1 vssd1 vccd1 vccd1 _06101_/B sky130_fd_sc_hd__nand3_1
X_07080_ _07080_/A _07080_/B _07088_/A vssd1 vssd1 vccd1 vccd1 _07082_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06031_ _06457_/B _06035_/C vssd1 vssd1 vccd1 vccd1 _06034_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07982_ _07929_/B _07928_/B _07928_/C vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10486__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _09721_/A vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__inv_2
X_06933_ _06933_/A _06933_/B vssd1 vssd1 vccd1 vccd1 _07090_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09652_ _09652_/A _09652_/B _09652_/C vssd1 vssd1 vccd1 vccd1 _09653_/B sky130_fd_sc_hd__nand3_1
X_06864_ _06864_/A _06864_/B vssd1 vssd1 vccd1 vccd1 _06865_/A sky130_fd_sc_hd__nand2_1
X_09583_ _09582_/B _09583_/B _09583_/C vssd1 vssd1 vccd1 vccd1 _09584_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__10050__B _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ _08604_/B _08604_/A vssd1 vssd1 vccd1 vccd1 _08603_/Y sky130_fd_sc_hd__nand2_1
X_06795_ _06795_/A _06795_/B vssd1 vssd1 vccd1 vccd1 _06796_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05425__A _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05815_ _05815_/A _05815_/B vssd1 vssd1 vccd1 vccd1 _06216_/B sky130_fd_sc_hd__nand2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08534_ _08800_/A _08800_/B _08802_/A vssd1 vssd1 vccd1 vccd1 _08540_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05746_ _05891_/C vssd1 vssd1 vccd1 vccd1 _05890_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08455__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ _08465_/A vssd1 vssd1 vccd1 vccd1 _08467_/B sky130_fd_sc_hd__inv_2
X_05677_ _05686_/A _06126_/A vssd1 vssd1 vccd1 vccd1 _06107_/B sky130_fd_sc_hd__nand2_1
X_08396_ _08621_/B vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07416_ _07416_/A _07416_/B vssd1 vssd1 vccd1 vccd1 _07418_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07347_ _07347_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07350_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09017_ _09017_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _09046_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07278_ _07315_/A vssd1 vssd1 vccd1 vccd1 _07283_/B sky130_fd_sc_hd__inv_2
X_06229_ _06357_/B vssd1 vssd1 vccd1 vccd1 _06358_/B sky130_fd_sc_hd__inv_2
XFILLER_0_20_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09919_ _09921_/C vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__inv_2
XFILLER_0_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10487_ _10495_/CLK hold38/X fanout99/X vssd1 vssd1 vccd1 vccd1 _10487_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07709__B _07709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09940__A _10171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05600_ _06121_/A _06121_/B vssd1 vssd1 vccd1 vccd1 _05605_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06580_ _06578_/Y _06094_/B _06579_/Y vssd1 vssd1 vccd1 vccd1 _06583_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05531_ _09816_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _05533_/A sky130_fd_sc_hd__nand2_1
X_08250_ _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__nand2_1
X_05462_ _05463_/B _05462_/B vssd1 vssd1 vccd1 vccd1 _05464_/A sky130_fd_sc_hd__nand2b_1
X_08181_ _08181_/A vssd1 vssd1 vccd1 vccd1 _08186_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07201_ _07228_/B _07227_/A vssd1 vssd1 vccd1 vccd1 _07202_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07132_ _07658_/A _07659_/A vssd1 vssd1 vccd1 vccd1 _07132_/Y sky130_fd_sc_hd__nand2_1
X_05393_ _05830_/B _05829_/A _05829_/B vssd1 vssd1 vccd1 vccd1 _05920_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07063_ _07063_/A _07063_/B vssd1 vssd1 vccd1 vccd1 _07064_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06014_ _06014_/A _06014_/B vssd1 vssd1 vccd1 vccd1 _06019_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07965_ _07988_/B vssd1 vssd1 vccd1 vccd1 _07989_/C sky130_fd_sc_hd__inv_2
X_09704_ _09540_/A _09540_/B _09541_/A vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__a21oi_1
X_06916_ _07007_/A _07008_/A vssd1 vssd1 vccd1 vccd1 _06916_/Y sky130_fd_sc_hd__nand2_1
X_09635_ _09903_/B _09635_/B vssd1 vssd1 vccd1 vccd1 _09638_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07896_ _08055_/A _07896_/B _08055_/B vssd1 vssd1 vccd1 vccd1 _08065_/B sky130_fd_sc_hd__nand3_2
X_06847_ _06847_/A _06847_/B vssd1 vssd1 vccd1 vccd1 _06850_/B sky130_fd_sc_hd__nand2_1
X_09566_ _09568_/B vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06778_ _06768_/Y _06856_/B _06777_/Y vssd1 vssd1 vccd1 vccd1 _06845_/A sky130_fd_sc_hd__a21oi_1
X_09497_ _09963_/A _09962_/A _09960_/B _09816_/B vssd1 vssd1 vccd1 vccd1 _09498_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10501__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ _08517_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__nand2_1
X_05729_ _05729_/A _05729_/B _05729_/C vssd1 vssd1 vccd1 vccd1 _05736_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_81_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08448_ _08449_/A _08448_/B vssd1 vssd1 vccd1 vccd1 _08673_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__05602__B _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08379_ _08382_/B _08382_/C vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__nand2_1
X_10410_ _10410_/A vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10341_ hold6/X _10336_/Y _10338_/B vssd1 vssd1 vccd1 vccd1 _10341_/Y sky130_fd_sc_hd__o21ai_1
X_10272_ _10272_/A _10299_/B vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09760__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05512__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07750_ _07767_/B _07754_/C vssd1 vssd1 vccd1 vccd1 _07752_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06701_ _06703_/A vssd1 vssd1 vccd1 vccd1 _06702_/B sky130_fd_sc_hd__inv_2
X_07681_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _07683_/A sky130_fd_sc_hd__nand2_1
X_09420_ _09420_/A _09420_/B vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08286__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06632_ _06638_/A _06632_/B _06632_/C vssd1 vssd1 vccd1 vccd1 _06633_/C sky130_fd_sc_hd__nand3_1
X_09351_ _09433_/A _09354_/C vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__nand2_1
X_06563_ _06564_/A _06564_/B vssd1 vssd1 vccd1 vccd1 _06565_/A sky130_fd_sc_hd__or2_1
XFILLER_0_59_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09282_ _10000_/A _09999_/A _09437_/B _09775_/B vssd1 vssd1 vccd1 vccd1 _09448_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08302_ _08582_/A vssd1 vssd1 vccd1 vccd1 _08303_/B sky130_fd_sc_hd__inv_2
X_05514_ _05998_/A _05998_/B vssd1 vssd1 vccd1 vccd1 _05515_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08233_ _09981_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__nand2_1
X_06494_ _06493_/B _08356_/B _06494_/C vssd1 vssd1 vccd1 vccd1 _08356_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05445_ input38/X _08814_/B vssd1 vssd1 vccd1 vccd1 _05447_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08164_ _08164_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08194_/B sky130_fd_sc_hd__nand2_1
X_05376_ _05376_/A _05376_/B vssd1 vssd1 vccd1 vccd1 _05377_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08095_ _08010_/Y _08095_/B vssd1 vssd1 vccd1 vccd1 _08096_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07115_ _07292_/C _07292_/B _07104_/Y vssd1 vssd1 vccd1 vccd1 _07116_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07046_ _07051_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08997_ _08997_/A vssd1 vssd1 vccd1 vccd1 _09003_/B sky130_fd_sc_hd__inv_2
X_07948_ _10083_/B _09988_/A vssd1 vssd1 vccd1 vccd1 _07950_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07879_ _07932_/B _07878_/Y vssd1 vssd1 vccd1 vccd1 _07928_/C sky130_fd_sc_hd__nor2b_1
X_09618_ _09612_/A _09612_/B _09615_/B vssd1 vssd1 vccd1 vccd1 _09619_/C sky130_fd_sc_hd__a21o_1
X_09549_ _10044_/A _10044_/C _09710_/D _10052_/A vssd1 vssd1 vccd1 vccd1 _09716_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06428__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10324_ _10322_/Y hold108/A vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__and2b_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10255_/A hold100/X vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__and2_1
XANTENNA__05820__B2 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05820__A1 _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ _10191_/A hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__and2_1
XANTENNA__05507__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05523__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05230_ input59/X vssd1 vssd1 vccd1 vccd1 _08688_/A sky130_fd_sc_hd__buf_8
XFILLER_0_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06073__B _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08920_ _09289_/C _08920_/B vssd1 vssd1 vccd1 vccd1 _08922_/A sky130_fd_sc_hd__xor2_1
X_08851_ _08899_/B _08851_/B _08851_/C vssd1 vssd1 vccd1 vccd1 _09141_/C sky130_fd_sc_hd__nand3_2
X_07802_ _07804_/B _07804_/C vssd1 vssd1 vccd1 vccd1 _07803_/A sky130_fd_sc_hd__nand2_1
X_08782_ _10027_/A _09710_/D _08781_/C vssd1 vssd1 vccd1 vccd1 _08786_/C sky130_fd_sc_hd__o21ai_1
X_05994_ _05994_/A _05995_/A vssd1 vssd1 vccd1 vccd1 _06018_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05417__B _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ _07733_/A _07733_/B vssd1 vssd1 vccd1 vccd1 _07734_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08728__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _07664_/A _07664_/B vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__nand2_1
X_09403_ _09663_/B _09403_/B vssd1 vssd1 vccd1 vccd1 _09408_/B sky130_fd_sc_hd__nand2_1
X_06615_ _08413_/B _06615_/B _06615_/C vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06248__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ _07728_/B _07725_/B vssd1 vssd1 vccd1 vccd1 _07595_/Y sky130_fd_sc_hd__nor2_1
X_09334_ _09334_/A vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__inv_2
XANTENNA__08744__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06546_ _09548_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _06549_/A sky130_fd_sc_hd__nand2_1
X_09265_ _09265_/A _09265_/B _09265_/C vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_62_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06477_ _06477_/A _06477_/B vssd1 vssd1 vccd1 vccd1 _06482_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09196_ _09196_/A _09196_/B vssd1 vssd1 vccd1 vccd1 _10452_/A sky130_fd_sc_hd__nand2_1
X_08216_ _08420_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _08219_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05428_ input31/X vssd1 vssd1 vccd1 vccd1 _09022_/D sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08147_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _08148_/B sky130_fd_sc_hd__nand2_1
X_05359_ _10026_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _05380_/A sky130_fd_sc_hd__nand2_1
X_08078_ _08176_/C vssd1 vssd1 vccd1 vccd1 _08079_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07029_ _07029_/A vssd1 vssd1 vccd1 vccd1 _07032_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10040_ _10039_/Y _10023_/B _10022_/Y vssd1 vssd1 vccd1 vccd1 _10041_/C sky130_fd_sc_hd__a21oi_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09485__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06902__A _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ hold116/X vssd1 vssd1 vccd1 vccd1 _10496_/D sky130_fd_sc_hd__clkbuf_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ hold91/X _10250_/B vssd1 vssd1 vccd1 vccd1 _10244_/A sky130_fd_sc_hd__nand2_1
X_10169_ _10168_/B _10169_/B _10169_/C vssd1 vssd1 vccd1 vccd1 _10172_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05253__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06068__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06400_ _06196_/C _06196_/B _06399_/Y vssd1 vssd1 vccd1 vccd1 _08655_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07380_ _07380_/A _07380_/B vssd1 vssd1 vccd1 vccd1 _07528_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06331_ _06331_/A _06331_/B _06331_/C vssd1 vssd1 vccd1 vccd1 _06736_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09050_ _09048_/Y _08764_/B _09049_/Y vssd1 vssd1 vccd1 vccd1 _09399_/A sky130_fd_sc_hd__a21oi_2
X_06262_ _06264_/A vssd1 vssd1 vccd1 vccd1 _06263_/B sky130_fd_sc_hd__inv_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08001_ _08001_/A _08014_/A vssd1 vssd1 vccd1 vccd1 _08002_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05213_ input55/X vssd1 vssd1 vccd1 vccd1 _08214_/A sky130_fd_sc_hd__buf_8
XFILLER_0_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06193_ _06198_/B _06198_/C vssd1 vssd1 vccd1 vccd1 _06399_/B sky130_fd_sc_hd__nand2_1
X_09952_ _09952_/A vssd1 vssd1 vccd1 vccd1 _09956_/A sky130_fd_sc_hd__inv_2
X_08903_ _09987_/A input19/X vssd1 vssd1 vccd1 vccd1 _08904_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09883_ _10140_/A vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__inv_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08836_/B vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__inv_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _08764_/B _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07716_ _07716_/A vssd1 vssd1 vccd1 vccd1 _08210_/A sky130_fd_sc_hd__inv_2
X_05977_ _05977_/A _05977_/B vssd1 vssd1 vccd1 vccd1 _05977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08696_ _08696_/A _08933_/A vssd1 vssd1 vccd1 vccd1 _08697_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07647_ _07647_/A _07647_/B _07647_/C vssd1 vssd1 vccd1 vccd1 _07651_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ _07564_/B _07761_/A _07562_/Y vssd1 vssd1 vccd1 vccd1 _07579_/B sky130_fd_sc_hd__a21oi_1
X_09317_ _09318_/B _09318_/A vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__or2_1
X_06529_ _06537_/A _08361_/A vssd1 vssd1 vccd1 vccd1 _06536_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09248_ _09581_/A _09248_/B _09641_/A vssd1 vssd1 vccd1 vccd1 _09252_/C sky130_fd_sc_hd__nand3_1
X_09179_ _09182_/B _09182_/C vssd1 vssd1 vccd1 vccd1 _09180_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06722__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 _10480_/Q vssd1 vssd1 vccd1 vccd1 y_o[0] sky130_fd_sc_hd__buf_12
Xoutput88 _10482_/Q vssd1 vssd1 vccd1 vccd1 y_o[2] sky130_fd_sc_hd__buf_12
Xoutput77 hold85/A vssd1 vssd1 vccd1 vccd1 y_o[1] sky130_fd_sc_hd__buf_12
X_10023_ _10023_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _10023_/X sky130_fd_sc_hd__and2_1
XFILLER_0_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09199__B _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06880_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _06885_/C sky130_fd_sc_hd__nand2_1
X_05900_ _05900_/A vssd1 vssd1 vccd1 vccd1 _06211_/B sky130_fd_sc_hd__inv_2
X_05831_ _05920_/C _05920_/B vssd1 vssd1 vccd1 vccd1 _05852_/B sky130_fd_sc_hd__nand2_1
X_08550_ input43/X _08814_/B vssd1 vssd1 vccd1 vccd1 _08551_/C sky130_fd_sc_hd__nand2_1
X_05762_ _05762_/A _05772_/A vssd1 vssd1 vccd1 vccd1 _05814_/B sky130_fd_sc_hd__nand2_1
X_08481_ _10027_/B _09953_/A _08479_/C vssd1 vssd1 vccd1 vccd1 _08485_/C sky130_fd_sc_hd__o21ai_1
X_05693_ _05694_/C _05694_/B _05694_/A vssd1 vssd1 vccd1 vccd1 _05693_/Y sky130_fd_sc_hd__a21oi_1
X_07501_ _07501_/A _07501_/B vssd1 vssd1 vccd1 vccd1 _07571_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07432_ _07507_/A _07508_/C vssd1 vssd1 vccd1 vccd1 _07432_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09102_ _09102_/A _09102_/B vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06526__B _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ _07363_/A _07363_/B _07363_/C vssd1 vssd1 vccd1 vccd1 _07370_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07294_ _08337_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _07299_/A sky130_fd_sc_hd__nand2_1
X_06314_ _06314_/A _06314_/B vssd1 vssd1 vccd1 vccd1 _06654_/A sky130_fd_sc_hd__nand2_1
X_09033_ _10050_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09039_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06245_ _06232_/Y _06368_/B _06244_/Y vssd1 vssd1 vccd1 vccd1 _06377_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06176_ _06176_/A _06176_/B vssd1 vssd1 vccd1 vccd1 _06178_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _09935_/A vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__inv_2
XFILLER_0_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09866_ _09869_/B _09866_/B _09866_/C vssd1 vssd1 vccd1 vccd1 _09877_/C sky130_fd_sc_hd__nand3b_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _08817_/A _09028_/A vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__nand2_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09797_ _09800_/B _09800_/C vssd1 vssd1 vccd1 vccd1 _09798_/A sky130_fd_sc_hd__nand2_1
X_08748_ _08748_/A _08747_/Y vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__nor2b_1
X_08679_ _09986_/A input17/X vssd1 vssd1 vccd1 vccd1 _08680_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08916__B _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10045__A2 _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08651__B _08651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07548__A _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10006_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08098__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05531__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06346__B _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06030_ _06030_/A _06030_/B vssd1 vssd1 vccd1 vccd1 _06035_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07981_ _08037_/B _08036_/B _07980_/Y vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09720_ _10050_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09721_/A sky130_fd_sc_hd__nand2_1
X_06932_ _06934_/A vssd1 vssd1 vccd1 vccd1 _06933_/B sky130_fd_sc_hd__inv_2
XANTENNA__08289__A _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10487__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09651_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__nand2_1
X_06863_ _06863_/A _06863_/B _06863_/C vssd1 vssd1 vccd1 vccd1 _07024_/B sky130_fd_sc_hd__nand3_1
X_09582_ _09582_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09911_/A sky130_fd_sc_hd__nand2_1
X_08602_ _08635_/A _08635_/B vssd1 vssd1 vccd1 vccd1 _08634_/A sky130_fd_sc_hd__nand2_1
X_06794_ _06796_/B _06795_/B _06795_/A vssd1 vssd1 vccd1 vccd1 _06797_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__05425__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05814_ _05814_/A _05814_/B _05814_/C vssd1 vssd1 vccd1 vccd1 _05815_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08533_ _08292_/B _08532_/Y _08290_/A vssd1 vssd1 vccd1 vccd1 _08802_/A sky130_fd_sc_hd__a21oi_2
X_05745_ _06205_/A _05745_/B vssd1 vssd1 vccd1 vccd1 _05891_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08464_ _08464_/A _08464_/B vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__nand2_1
X_05676_ _05675_/B _06126_/B _05676_/C vssd1 vssd1 vccd1 vccd1 _06126_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _08397_/B _08397_/A vssd1 vssd1 vccd1 vccd1 _08621_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07415_ _07415_/A _07415_/B _07415_/C vssd1 vssd1 vccd1 vccd1 _07419_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_18_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07346_ _07346_/A _07346_/B vssd1 vssd1 vccd1 vccd1 _07347_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ _09018_/A vssd1 vssd1 vccd1 vccd1 _09017_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07277_ _07259_/C _07259_/B _07253_/Y vssd1 vssd1 vccd1 vccd1 _07315_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06228_ _10043_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _06357_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06159_ _06604_/B _06159_/B vssd1 vssd1 vccd1 vccd1 _06162_/C sky130_fd_sc_hd__nand2_1
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09921_/C sky130_fd_sc_hd__nor2_1
X_09849_ _09925_/A _09925_/C vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07831__A _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06447__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05351__A _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10486_ _10494_/CLK _10486_/D fanout98/X vssd1 vssd1 vccd1 vccd1 _10486_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__05526__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05530_ _05534_/A _05534_/C vssd1 vssd1 vccd1 vccd1 _05532_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05461_ _05431_/Y _05461_/B _05461_/C vssd1 vssd1 vccd1 vccd1 _05826_/A sky130_fd_sc_hd__nand3b_1
X_08180_ _08180_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__nand2_1
X_07200_ _07227_/A _07228_/B vssd1 vssd1 vccd1 vccd1 _07203_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05392_ _05392_/A _05392_/B vssd1 vssd1 vccd1 vccd1 _05829_/B sky130_fd_sc_hd__nand2_1
X_07131_ _07125_/Y _07627_/B _07130_/Y vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07062_ _07088_/A vssd1 vssd1 vccd1 vccd1 _07079_/B sky130_fd_sc_hd__inv_2
X_06013_ _06451_/A _06013_/B _06013_/C vssd1 vssd1 vccd1 vccd1 _06014_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_2_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06820__A _06820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ _07964_/A _07971_/A vssd1 vssd1 vccd1 vccd1 _07988_/B sky130_fd_sc_hd__nand2_1
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06915_ _06890_/Y _07020_/B _06914_/Y vssd1 vssd1 vccd1 vccd1 _07008_/A sky130_fd_sc_hd__a21oi_2
X_07895_ _07902_/B _07902_/A vssd1 vssd1 vccd1 vccd1 _08055_/B sky130_fd_sc_hd__nand2_1
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09635_/B sky130_fd_sc_hd__nand2_1
X_06846_ _06768_/Y _06856_/B _06777_/Y vssd1 vssd1 vccd1 vccd1 _06847_/A sky130_fd_sc_hd__a21o_1
X_09565_ _09565_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09568_/B sky130_fd_sc_hd__xor2_1
X_06777_ _06854_/A _06853_/A vssd1 vssd1 vccd1 vccd1 _06777_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _09960_/A _09496_/B vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__nand2_1
X_08516_ _08517_/A _08672_/B _08516_/C vssd1 vssd1 vccd1 vccd1 _08672_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_65_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05728_ _05728_/A _05728_/B vssd1 vssd1 vccd1 vccd1 _06176_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08447_ _08449_/C _08449_/B vssd1 vssd1 vccd1 vccd1 _08448_/B sky130_fd_sc_hd__nand2_1
X_05659_ _09685_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _05662_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08482__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ _08378_/A _08378_/B _08604_/A vssd1 vssd1 vccd1 vccd1 _08382_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07329_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07329_/Y sky130_fd_sc_hd__inv_2
X_10340_ _10340_/A hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__xor2_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _10299_/B _10272_/A vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07561__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10476__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07736__A _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ _10495_/CLK _10469_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09951__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05256__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ _06703_/B _06703_/C vssd1 vssd1 vccd1 vccd1 _06702_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07680_ _07680_/A _07680_/B _07680_/C vssd1 vssd1 vccd1 vccd1 _07681_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08286__B _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06631_ _06631_/A _06637_/B vssd1 vssd1 vccd1 vccd1 _09188_/A sky130_fd_sc_hd__nand2_2
X_09350_ _09350_/A _09350_/B vssd1 vssd1 vccd1 vccd1 _09354_/C sky130_fd_sc_hd__nand2_1
X_06562_ input46/X _08337_/B vssd1 vssd1 vccd1 vccd1 _06564_/B sky130_fd_sc_hd__nand2_1
X_09281_ _09951_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _09286_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08301_ _08299_/Y _06458_/B _08300_/Y vssd1 vssd1 vccd1 vccd1 _08582_/A sky130_fd_sc_hd__a21oi_4
X_05513_ _05518_/C vssd1 vssd1 vccd1 vccd1 _05515_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08232_ _09951_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__nand2_1
X_06493_ _06493_/A _06493_/B vssd1 vssd1 vccd1 vccd1 _06495_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05444_ input29/X vssd1 vssd1 vccd1 vccd1 _08814_/B sky130_fd_sc_hd__clkbuf_8
X_08163_ _08163_/A _08189_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05375_ _05913_/A _05908_/A vssd1 vssd1 vccd1 vccd1 _05375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08094_ _08033_/B _08032_/B _08032_/C vssd1 vssd1 vccd1 vccd1 _08134_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07114_ _07114_/A _07114_/B vssd1 vssd1 vccd1 vccd1 _07116_/A sky130_fd_sc_hd__nand2_1
X_07045_ _08780_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _07060_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08996_ _10026_/A _10052_/A vssd1 vssd1 vccd1 vccd1 _08997_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07947_ _09854_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _07950_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08477__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _09392_/D _09953_/A _07877_/C vssd1 vssd1 vccd1 vccd1 _07878_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09617_ _09617_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _09619_/B sky130_fd_sc_hd__or2b_1
X_06829_ _06829_/A _06829_/B _06829_/C vssd1 vssd1 vccd1 vccd1 _07146_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_78_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09548_ _09548_/A vssd1 vssd1 vccd1 vccd1 _10044_/C sky130_fd_sc_hd__inv_2
XANTENNA__10499__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10323_ _10499_/Q hold107/X vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10254_ _10254_/A _10266_/A vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__nand2_1
XANTENNA__05820__A2 _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10185_ hold54/X _10381_/B vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05523__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08850_ _08850_/A vssd1 vssd1 vccd1 vccd1 _08851_/C sky130_fd_sc_hd__inv_2
X_07801_ _07801_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07804_/C sky130_fd_sc_hd__nand2_1
X_08781_ _10027_/A _09710_/D _08781_/C vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__or3_1
X_05993_ _09951_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _05995_/A sky130_fd_sc_hd__nand2_1
X_07732_ _07816_/B _07816_/C vssd1 vssd1 vccd1 vccd1 _07817_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05714__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _07667_/A _07667_/B _07666_/B vssd1 vssd1 vccd1 vccd1 _07664_/B sky130_fd_sc_hd__nand3_1
X_09402_ _09663_/A vssd1 vssd1 vccd1 vccd1 _09403_/B sky130_fd_sc_hd__inv_2
X_06614_ _06616_/A _06617_/A vssd1 vssd1 vccd1 vccd1 _06615_/C sky130_fd_sc_hd__nand2_1
X_09333_ _09575_/B _09334_/A vssd1 vssd1 vccd1 vccd1 _09339_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07594_ _07731_/C vssd1 vssd1 vccd1 vccd1 _07730_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ _06576_/B _06576_/C vssd1 vssd1 vccd1 vccd1 _06575_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09264_ _09264_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06476_ _06477_/A _06477_/B vssd1 vssd1 vccd1 vccd1 _08281_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09195_ _09190_/Y _09191_/Y _09194_/Y vssd1 vssd1 vccd1 vccd1 _09196_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08215_ _08215_/A vssd1 vssd1 vccd1 vccd1 _08223_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05427_ input35/X vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__clkbuf_8
X_08146_ _08147_/B _08147_/A vssd1 vssd1 vccd1 vccd1 _08148_/A sky130_fd_sc_hd__or2_1
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05358_ _05927_/A _05928_/A vssd1 vssd1 vccd1 vccd1 _05911_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05289_ _05338_/A vssd1 vssd1 vccd1 vccd1 _05337_/B sky130_fd_sc_hd__inv_2
X_08077_ _08077_/A _08077_/B vssd1 vssd1 vccd1 vccd1 _08202_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07028_ _07032_/A _07029_/A vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _08978_/B _08979_/B _08979_/C vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__08919__B input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08935__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09485__B _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06902__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10306_ hold115/X _10311_/A vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__and2_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ _10250_/B hold91/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__or2_1
X_10168_ _10168_/A _10168_/B vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__nand2_1
X_10099_ _10102_/B _10102_/C vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05253__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06330_ _06330_/A _06330_/B vssd1 vssd1 vccd1 vccd1 _06736_/B sky130_fd_sc_hd__nand2_1
X_06261_ _06264_/B _06264_/C vssd1 vssd1 vccd1 vccd1 _06263_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08000_ _08014_/B _08000_/B _08000_/C vssd1 vssd1 vccd1 vccd1 _08014_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05212_ input9/X vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06192_ _06199_/C vssd1 vssd1 vccd1 vccd1 _06196_/B sky130_fd_sc_hd__inv_2
XFILLER_0_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ _09951_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05709__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08902_ input20/X vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09882_ _09616_/C _09616_/B _09613_/Y vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__a21oi_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08833_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _08836_/B sky130_fd_sc_hd__nand2_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__nand2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05976_ _05977_/B _05977_/A vssd1 vssd1 vccd1 vccd1 _05976_/Y sky130_fd_sc_hd__nand2_1
X_07715_ _07715_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__nor2_1
X_08695_ _08933_/B _08695_/B _08695_/C vssd1 vssd1 vccd1 vccd1 _08933_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07646_ _07642_/Y _07410_/A _07643_/Y vssd1 vssd1 vccd1 vccd1 _07647_/A sky130_fd_sc_hd__a21oi_1
X_07577_ _07577_/A vssd1 vssd1 vccd1 vccd1 _07761_/A sky130_fd_sc_hd__inv_2
X_09316_ _09484_/B _09316_/B vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06528_ _06527_/B _08361_/B _06528_/C vssd1 vssd1 vccd1 vccd1 _08361_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _09641_/B _09247_/B vssd1 vssd1 vccd1 vccd1 _09252_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06459_ _06458_/B _06459_/B _06459_/C vssd1 vssd1 vccd1 vccd1 _06460_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_90_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09178_ _09178_/A _09178_/B vssd1 vssd1 vccd1 vccd1 _09182_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _08194_/A _08132_/A vssd1 vssd1 vccd1 vccd1 _08130_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06722__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput67 hold99/A vssd1 vssd1 vccd1 vccd1 y_o[10] sky130_fd_sc_hd__buf_12
Xoutput89 hold21/A vssd1 vssd1 vccd1 vccd1 y_o[30] sky130_fd_sc_hd__buf_12
Xoutput78 _10500_/Q vssd1 vssd1 vccd1 vccd1 y_o[20] sky130_fd_sc_hd__buf_12
X_10022_ _10039_/B _10039_/A vssd1 vssd1 vccd1 vccd1 _10022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05354__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09199__C _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09496__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05830_ _05830_/A _05830_/B vssd1 vssd1 vccd1 vccd1 _05920_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05761_ _05879_/C _05879_/B _05760_/Y vssd1 vssd1 vccd1 vccd1 _05772_/A sky130_fd_sc_hd__a21oi_2
X_07500_ _07556_/C _07496_/Y _07556_/A vssd1 vssd1 vccd1 vccd1 _07501_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08480_ _08480_/A vssd1 vssd1 vccd1 vccd1 _08737_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05692_ _05486_/C _05486_/B _05478_/Y vssd1 vssd1 vccd1 vccd1 _05694_/A sky130_fd_sc_hd__a21o_1
X_07431_ _07483_/C _07483_/B _07480_/A vssd1 vssd1 vccd1 vccd1 _07508_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07362_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07370_/A sky130_fd_sc_hd__nand2_1
X_09101_ _08882_/C _08882_/B _08878_/Y vssd1 vssd1 vccd1 vccd1 _09102_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06313_ _06313_/A _06313_/B _06313_/C vssd1 vssd1 vccd1 vccd1 _06314_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07293_ _07303_/A _07303_/B vssd1 vssd1 vccd1 vccd1 _07366_/B sky130_fd_sc_hd__nand2_1
X_09032_ _09042_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__nand2_1
X_06244_ _06366_/A _06365_/A vssd1 vssd1 vccd1 vccd1 _06244_/Y sky130_fd_sc_hd__nor2_1
X_06175_ _06175_/A _06175_/B vssd1 vssd1 vccd1 vccd1 _06176_/B sky130_fd_sc_hd__or2_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05439__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09934_ _09934_/A _09935_/A vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__nand2_1
X_09865_ _10091_/A _09867_/B _09868_/B vssd1 vssd1 vccd1 vccd1 _09866_/C sky130_fd_sc_hd__nand3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _08815_/B _09028_/B _08816_/C vssd1 vssd1 vccd1 vccd1 _09028_/A sky130_fd_sc_hd__nand3b_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _09796_/A _09796_/B _09796_/C vssd1 vssd1 vccd1 vccd1 _09800_/C sky130_fd_sc_hd__nand3_1
X_08747_ _09227_/A _09686_/D _08746_/C vssd1 vssd1 vccd1 vccd1 _08747_/Y sky130_fd_sc_hd__o21ai_1
X_05959_ _05959_/A _05959_/B vssd1 vssd1 vccd1 vccd1 _05963_/B sky130_fd_sc_hd__nand2_1
X_08678_ _08678_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08682_/C sky130_fd_sc_hd__nand2_1
X_07629_ _07635_/B _07635_/C vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05349__A _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10005_ _10006_/B _10006_/A vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__or2_1
XANTENNA__08098__C _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05531__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07739__A _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05259__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07980_ _08034_/A _07980_/B vssd1 vssd1 vccd1 vccd1 _07980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06931_ _06934_/B _06934_/C vssd1 vssd1 vccd1 vccd1 _06933_/A sky130_fd_sc_hd__nand2_1
X_09650_ _09652_/C vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__inv_2
XANTENNA__09392__C _09392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08601_ _09147_/A _08601_/B _08601_/C vssd1 vssd1 vccd1 vccd1 _08635_/B sky130_fd_sc_hd__nand3_1
X_06862_ _06864_/B _06862_/B vssd1 vssd1 vccd1 vccd1 _06863_/B sky130_fd_sc_hd__nand2_1
X_09581_ _09581_/A _09581_/B vssd1 vssd1 vccd1 vccd1 _09582_/B sky130_fd_sc_hd__nand2_1
X_06793_ _06793_/A _06793_/B vssd1 vssd1 vccd1 vccd1 _06795_/A sky130_fd_sc_hd__nand2_1
X_05813_ _05813_/A _05813_/B vssd1 vssd1 vccd1 vccd1 _05815_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08532_ _08532_/A vssd1 vssd1 vccd1 vccd1 _08532_/Y sky130_fd_sc_hd__inv_2
X_05744_ _05744_/A _05821_/A vssd1 vssd1 vccd1 vccd1 _05745_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08463_ _08463_/A _08757_/A _08719_/A vssd1 vssd1 vccd1 vccd1 _08467_/C sky130_fd_sc_hd__nand3_1
XANTENNA__05722__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05675_ _05675_/A _05675_/B vssd1 vssd1 vccd1 vccd1 _05686_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ _07416_/B _07417_/B _07417_/C vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__nand3_1
X_08394_ _06560_/A _06566_/B _06565_/A vssd1 vssd1 vccd1 vccd1 _08397_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07345_ _07345_/A _07345_/B _07345_/C vssd1 vssd1 vccd1 vccd1 _07350_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07276_ _07283_/A _07283_/C vssd1 vssd1 vccd1 vccd1 _07315_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _09013_/Y _08797_/B _09014_/Y vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06227_ _06353_/A _06354_/A vssd1 vssd1 vccd1 vccd1 _06358_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06158_ _06158_/A _06158_/B vssd1 vssd1 vccd1 vccd1 _06159_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06089_ _06579_/A vssd1 vssd1 vccd1 vccd1 _06090_/B sky130_fd_sc_hd__inv_2
X_09917_ _09917_/A vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__inv_2
X_09848_ _10078_/A _09848_/B _09848_/C vssd1 vssd1 vccd1 vccd1 _09925_/C sky130_fd_sc_hd__nand3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09777_/A _09777_/B _09777_/C vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__07831__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06447__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10485_ _10495_/CLK _10485_/D fanout98/X vssd1 vssd1 vccd1 vccd1 _10485_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07294__A _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05526__B _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05542__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05460_ _05493_/A _05493_/B vssd1 vssd1 vccd1 vccd1 _05491_/A sky130_fd_sc_hd__nand2_1
X_05391_ _05391_/A _05391_/B vssd1 vssd1 vccd1 vccd1 _05829_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07130_ _07623_/A _07625_/A vssd1 vssd1 vccd1 vccd1 _07130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07061_ _07054_/C _07054_/B _07060_/Y vssd1 vssd1 vccd1 vccd1 _07088_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_42_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09684__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06012_ _06012_/A vssd1 vssd1 vccd1 vccd1 _06013_/B sky130_fd_sc_hd__inv_2
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07963_ _07971_/B _07963_/B _07963_/C vssd1 vssd1 vccd1 vccd1 _07971_/A sky130_fd_sc_hd__nand3_1
X_09702_ _09702_/A vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__inv_2
X_06914_ _07013_/A _07018_/A vssd1 vssd1 vccd1 vccd1 _06914_/Y sky130_fd_sc_hd__nor2_1
X_07894_ _07796_/Y _07889_/B _07797_/Y vssd1 vssd1 vccd1 vccd1 _07902_/A sky130_fd_sc_hd__a21oi_1
X_09633_ _09634_/B _09634_/A vssd1 vssd1 vccd1 vccd1 _09903_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06845_ _06845_/A _06845_/B _06845_/C vssd1 vssd1 vccd1 vccd1 _06850_/A sky130_fd_sc_hd__nand3_1
X_09564_ _09564_/A _09563_/X vssd1 vssd1 vccd1 vccd1 _09565_/B sky130_fd_sc_hd__or2b_1
X_08515_ _08518_/B vssd1 vssd1 vccd1 vccd1 _08516_/C sky130_fd_sc_hd__inv_2
X_06776_ _06857_/C vssd1 vssd1 vccd1 vccd1 _06856_/B sky130_fd_sc_hd__inv_2
X_09495_ _09828_/A _09495_/B vssd1 vssd1 vccd1 vccd1 _09503_/C sky130_fd_sc_hd__nand2_1
X_05727_ _05729_/C vssd1 vssd1 vccd1 vccd1 _05728_/B sky130_fd_sc_hd__inv_2
XFILLER_0_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08446_ _08446_/A _08700_/A vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05658_ _05662_/A vssd1 vssd1 vccd1 vccd1 _05661_/A sky130_fd_sc_hd__inv_2
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08377_ _08377_/A vssd1 vssd1 vccd1 vccd1 _08604_/A sky130_fd_sc_hd__inv_2
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08482__B _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ _09951_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _07459_/A sky130_fd_sc_hd__nand2_1
X_05589_ _05610_/A _05610_/C vssd1 vssd1 vccd1 vccd1 _05609_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06283__A _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07259_ _07253_/Y _07259_/B _07259_/C vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__09023__B1 _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ _10267_/Y _10268_/Y hold104/X vssd1 vssd1 vccd1 vccd1 _10272_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08938__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__B _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10468_ _10494_/CLK _10468_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07736__B input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06640__B _06640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ _08200_/A _08200_/B _08086_/A vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09951__B _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05256__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ _06638_/A vssd1 vssd1 vccd1 vccd1 _06637_/B sky130_fd_sc_hd__inv_2
XANTENNA__05272__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ _10051_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _06564_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09280_ _09479_/B _09304_/B vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__nand2_1
X_06492_ _09960_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _06493_/B sky130_fd_sc_hd__nand2_1
X_08300_ _08300_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08300_/Y sky130_fd_sc_hd__nor2_1
X_05512_ _09963_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _05518_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08231_ _08231_/A vssd1 vssd1 vccd1 vccd1 _08237_/A sky130_fd_sc_hd__inv_2
X_05443_ _05448_/A _05448_/C vssd1 vssd1 vccd1 vccd1 _05446_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _08188_/B _08179_/A vssd1 vssd1 vccd1 vccd1 _08189_/A sky130_fd_sc_hd__nor2_1
X_05374_ _05911_/B _05911_/C _05373_/Y vssd1 vssd1 vccd1 vccd1 _05908_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06606__A2 _06173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ _08130_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08125_/A sky130_fd_sc_hd__nand2_1
X_07113_ _07113_/A _07114_/B _07114_/A vssd1 vssd1 vccd1 vccd1 _07356_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07044_ _07060_/A vssd1 vssd1 vccd1 vccd1 _07051_/A sky130_fd_sc_hd__inv_2
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08995_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _09011_/B sky130_fd_sc_hd__and2_1
X_07946_ _09601_/B _09986_/A vssd1 vssd1 vccd1 vccd1 _08003_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10471__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _09392_/D _09953_/A _07877_/C vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_97_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09616_ _09613_/Y _09616_/B _09616_/C vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06828_ _06828_/A vssd1 vssd1 vccd1 vccd1 _06829_/C sky130_fd_sc_hd__inv_2
X_09547_ _10043_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _09553_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06759_ _06759_/A _06759_/B _06759_/C vssd1 vssd1 vccd1 vccd1 _06854_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09478_ _09799_/A _09482_/C vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08429_ _08674_/A _08432_/C vssd1 vssd1 vccd1 vccd1 _08431_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10322_ _10499_/Q hold107/X vssd1 vssd1 vccd1 vccd1 _10322_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07837__A _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ _10266_/A _10254_/A vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__or2_1
XFILLER_0_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10184_ _10381_/B hold54/X vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09962__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08780_ _09685_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08781_/C sky130_fd_sc_hd__nand2_1
X_07800_ _07597_/Y _07721_/B _07604_/Y vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__a21o_1
X_05992_ _05996_/A _05996_/C vssd1 vssd1 vccd1 vccd1 _05994_/A sky130_fd_sc_hd__nand2_1
X_07731_ _07731_/A _07731_/B _07731_/C vssd1 vssd1 vccd1 vccd1 _07816_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05714__B input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ _07666_/A _07667_/C vssd1 vssd1 vccd1 vccd1 _07664_/A sky130_fd_sc_hd__nand2_1
X_09401_ _09401_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__nor2_2
X_06613_ _06401_/Y _06182_/B _06402_/Y vssd1 vssd1 vccd1 vccd1 _06617_/A sky130_fd_sc_hd__a21oi_1
X_07593_ _07593_/A _07600_/A vssd1 vssd1 vccd1 vccd1 _07731_/C sky130_fd_sc_hd__nand2_1
X_09332_ _09332_/A _09332_/B vssd1 vssd1 vccd1 vccd1 _09334_/A sky130_fd_sc_hd__nand2_1
X_06544_ _06544_/A _08365_/A _06544_/C vssd1 vssd1 vccd1 vccd1 _06576_/C sky130_fd_sc_hd__nand3_1
X_09263_ _09265_/B vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06475_ _10026_/B _08272_/B vssd1 vssd1 vccd1 vccd1 _06477_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09194_ _09194_/A _09194_/B vssd1 vssd1 vccd1 vccd1 _09194_/Y sky130_fd_sc_hd__nand2_1
X_08214_ _08214_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__nand2_1
X_05426_ _05462_/B _05463_/B vssd1 vssd1 vccd1 vccd1 _05461_/C sky130_fd_sc_hd__nand2_1
X_08145_ _08140_/Y _08144_/Y _08144_/A vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_43_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05357_ _05937_/C _05937_/B _05356_/Y vssd1 vssd1 vccd1 vccd1 _05928_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06561__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05288_ _05500_/A _05502_/A _05293_/B vssd1 vssd1 vccd1 vccd1 _05335_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _10400_/B _08086_/B vssd1 vssd1 vccd1 vccd1 _08077_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10083__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07027_ _07030_/B vssd1 vssd1 vccd1 vccd1 _07032_/A sky130_fd_sc_hd__inv_2
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _08978_/A _08978_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__nand2_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10466__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _08040_/B _07929_/B vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__nand2_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08935__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05640__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09485__C _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10305_ _10305_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__nand2_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10236_ _10226_/Y _10235_/Y hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__o21ai_2
X_10167_ _10169_/B _10169_/C vssd1 vssd1 vccd1 vccd1 _10168_/A sky130_fd_sc_hd__nand2_1
X_10098_ _10098_/A _10098_/B _10098_/C vssd1 vssd1 vccd1 vccd1 _10102_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_16_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09022__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06260_ _06260_/A _06260_/B _06260_/C vssd1 vssd1 vccd1 vccd1 _06264_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08861__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05211_ _05216_/B _05251_/A vssd1 vssd1 vccd1 vccd1 _05215_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06191_ _06635_/C _06191_/B vssd1 vssd1 vccd1 vccd1 _06199_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09950_ _09792_/A _09792_/C _09792_/B vssd1 vssd1 vccd1 vccd1 _09950_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__05709__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08901_ _08901_/A _08901_/B vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09881_ _09885_/A _09885_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__nand2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08832_ _08832_/A _08832_/B _08832_/C vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__nand3_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08763_ _08763_/A _08763_/B vssd1 vssd1 vccd1 vccd1 _08764_/B sky130_fd_sc_hd__nand2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05975_ _06394_/C _06394_/B _05974_/Y vssd1 vssd1 vccd1 vccd1 _06628_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07714_ _07714_/A _07716_/A vssd1 vssd1 vccd1 vccd1 _07715_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08694_ _08933_/B _08695_/C _08695_/B vssd1 vssd1 vccd1 vccd1 _08696_/A sky130_fd_sc_hd__a21o_1
X_07645_ _07645_/A _07645_/B vssd1 vssd1 vccd1 vccd1 _07697_/A sky130_fd_sc_hd__nand2_2
X_07576_ _07580_/B _07580_/C vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__nand2_1
X_09315_ _09963_/B _09485_/C _09962_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _09316_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06527_ _06527_/A _06527_/B vssd1 vssd1 vccd1 vccd1 _06537_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _09641_/A vssd1 vssd1 vccd1 vccd1 _09247_/B sky130_fd_sc_hd__inv_2
X_06458_ _06458_/A _06458_/B vssd1 vssd1 vccd1 vccd1 _06460_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05409_ _05590_/A vssd1 vssd1 vccd1 vccd1 _05413_/A sky130_fd_sc_hd__inv_2
XFILLER_0_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09177_ _09191_/B vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__inv_4
XFILLER_0_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06389_ _06276_/A _06277_/C _06314_/A vssd1 vssd1 vccd1 vccd1 _06812_/B sky130_fd_sc_hd__o21ai_2
X_08128_ _08128_/A _08128_/B vssd1 vssd1 vccd1 vccd1 _08132_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08059_ _08087_/B _08059_/B vssd1 vssd1 vccd1 vccd1 _08060_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10021_ _10075_/B _10075_/C vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__nand2_1
Xoutput79 _10501_/Q vssd1 vssd1 vccd1 vccd1 y_o[21] sky130_fd_sc_hd__buf_12
Xoutput68 _10491_/Q vssd1 vssd1 vccd1 vccd1 y_o[11] sky130_fd_sc_hd__buf_12
XANTENNA__05635__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05354__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__A _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09199__D _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09496__B _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07297__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ _10486_/Q hold35/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05760_ _05760_/A _05760_/B vssd1 vssd1 vccd1 vccd1 _05760_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05691_ _05749_/C vssd1 vssd1 vccd1 vccd1 _05748_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07430_ _07430_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07480_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_92_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07361_ _07363_/A vssd1 vssd1 vccd1 vccd1 _07362_/B sky130_fd_sc_hd__inv_2
X_09100_ _09104_/B _09385_/A vssd1 vssd1 vccd1 vccd1 _09102_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06312_ _06312_/A vssd1 vssd1 vccd1 vccd1 _06313_/B sky130_fd_sc_hd__inv_2
X_09031_ _09031_/A _09356_/A _09031_/C vssd1 vssd1 vccd1 vccd1 _09042_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07292_ _07104_/Y _07292_/B _07292_/C vssd1 vssd1 vccd1 vccd1 _07303_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06243_ _06782_/C _06243_/B vssd1 vssd1 vccd1 vccd1 _06368_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06174_ _06179_/A _06179_/B vssd1 vssd1 vccd1 vccd1 _06177_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05439__B _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09864_ _09867_/A _09868_/C vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _08815_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__nand2_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09795_/A vssd1 vssd1 vccd1 vccd1 _09796_/B sky130_fd_sc_hd__inv_2
X_08746_ _09227_/A _09686_/D _08746_/C vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__nor3_1
X_05958_ _05960_/A vssd1 vssd1 vccd1 vccd1 _05959_/B sky130_fd_sc_hd__inv_2
XFILLER_0_95_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10504__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _08678_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08911_/B sky130_fd_sc_hd__or2_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05889_ _05891_/A _05891_/B vssd1 vssd1 vccd1 vccd1 _05890_/A sky130_fd_sc_hd__nand2_1
X_07628_ _07627_/B _07628_/B _07628_/C vssd1 vssd1 vccd1 vccd1 _07635_/C sky130_fd_sc_hd__nand3b_1
XANTENNA__06286__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07559_ _09854_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09597__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09229_ _09229_/A _09230_/B _09230_/A vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07829__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10004_ _10004_/A vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__inv_2
XFILLER_0_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__D _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08676__A _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07739__B input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05259__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ _06930_/A _06930_/B _06930_/C vssd1 vssd1 vccd1 vccd1 _06934_/C sky130_fd_sc_hd__nand3_1
X_08600_ _09147_/B _08600_/B vssd1 vssd1 vccd1 vccd1 _08635_/A sky130_fd_sc_hd__nand2_1
X_06861_ _06861_/A vssd1 vssd1 vccd1 vccd1 _06864_/B sky130_fd_sc_hd__inv_2
X_09580_ _09583_/B _09583_/C vssd1 vssd1 vccd1 vccd1 _09582_/A sky130_fd_sc_hd__nand2_1
X_06792_ _06792_/A vssd1 vssd1 vccd1 vccd1 _06793_/A sky130_fd_sc_hd__inv_2
X_05812_ _05814_/C vssd1 vssd1 vccd1 vccd1 _05813_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08531_ _08796_/B _08531_/B _08531_/C vssd1 vssd1 vccd1 vccd1 _08800_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05743_ _05821_/A _05744_/A vssd1 vssd1 vccd1 vccd1 _06205_/A sky130_fd_sc_hd__or2_2
X_08462_ _08757_/B _08462_/B vssd1 vssd1 vccd1 vccd1 _08467_/A sky130_fd_sc_hd__nand2_1
X_05674_ _10026_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _05675_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06818__B _07709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07413_ _07264_/Y _07470_/B _07287_/Y vssd1 vssd1 vccd1 vccd1 _07416_/B sky130_fd_sc_hd__a21o_1
X_08393_ input49/X _10126_/B vssd1 vssd1 vccd1 vccd1 _08397_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07344_ _07202_/A _07225_/B _07203_/A vssd1 vssd1 vccd1 vccd1 _07386_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09210__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07275_ _07275_/A _07275_/B vssd1 vssd1 vccd1 vccd1 _07283_/C sky130_fd_sc_hd__nand2_1
X_09014_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09014_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06226_ _09684_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _06354_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06157_ _06157_/A vssd1 vssd1 vccd1 vccd1 _06604_/B sky130_fd_sc_hd__inv_2
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06088_ _05560_/A _05563_/A _06087_/Y vssd1 vssd1 vccd1 vccd1 _06579_/A sky130_fd_sc_hd__a21oi_2
X_09916_ _09916_/A _09916_/B vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__nand2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09778_/A vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__inv_2
X_08729_ _08729_/A _09953_/A _08729_/C vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_68_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07559__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10494_/CLK _10484_/D fanout98/X vssd1 vssd1 vccd1 vccd1 _10484_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07294__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05542__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05390_ _05392_/B vssd1 vssd1 vccd1 vccd1 _05391_/B sky130_fd_sc_hd__inv_2
XFILLER_0_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07060_ _07060_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07060_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06011_ _06011_/A _06012_/A vssd1 vssd1 vccd1 vccd1 _06014_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09684__B _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06820__C _06820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _09701_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09701_/Y sky130_fd_sc_hd__nand2_1
X_07962_ _07971_/B _07963_/C _07963_/B vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__a21o_1
X_06913_ _07021_/C vssd1 vssd1 vccd1 vccd1 _07020_/B sky130_fd_sc_hd__inv_2
X_07893_ _07893_/A _07893_/B vssd1 vssd1 vccd1 vccd1 _07902_/B sky130_fd_sc_hd__nand2_1
X_09632_ _09632_/A _09632_/B vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__xor2_1
X_06844_ _06999_/B _06999_/C vssd1 vssd1 vccd1 vccd1 _07001_/B sky130_fd_sc_hd__nand2_1
X_09563_ input46/X _10050_/B _10051_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09563_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ _08514_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__nand2_1
X_06775_ _06775_/A _06775_/B vssd1 vssd1 vccd1 vccd1 _06857_/C sky130_fd_sc_hd__nand2_1
X_09494_ _09495_/B _09828_/A vssd1 vssd1 vccd1 vccd1 _09503_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05726_ _05726_/A _06185_/A vssd1 vssd1 vccd1 vccd1 _05729_/C sky130_fd_sc_hd__nand2_1
X_08445_ _08445_/A _08445_/B _08700_/B vssd1 vssd1 vccd1 vccd1 _08700_/A sky130_fd_sc_hd__nand3_1
X_05657_ _09528_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _05662_/A sky130_fd_sc_hd__nand2_1
X_08376_ _08604_/B _08377_/A vssd1 vssd1 vccd1 vccd1 _08382_/B sky130_fd_sc_hd__nand2_1
X_05588_ _05588_/A _05588_/B _05588_/C vssd1 vssd1 vccd1 vccd1 _05610_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07327_ _07330_/A _07330_/B vssd1 vssd1 vccd1 vccd1 _07327_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09271__A1 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07258_ _07258_/A vssd1 vssd1 vccd1 vccd1 _07259_/B sky130_fd_sc_hd__inv_2
XANTENNA__09023__A1 _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__B2 _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06209_ _06211_/C vssd1 vssd1 vccd1 vccd1 _06209_/Y sky130_fd_sc_hd__inv_2
X_07189_ _07241_/C _07241_/B _07188_/Y vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06474__A _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10467_ _10495_/CLK _10467_/D fanout99/X vssd1 vssd1 vccd1 vccd1 _10467_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__05818__A _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ _10398_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10461_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06560_ _06560_/A vssd1 vssd1 vccd1 vccd1 _06566_/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05272__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06491_ _08356_/B _06494_/C vssd1 vssd1 vccd1 vccd1 _06493_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05511_ _05517_/A _05516_/A vssd1 vssd1 vccd1 vccd1 _05515_/A sky130_fd_sc_hd__nand2_1
X_08230_ _09963_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _08231_/A sky130_fd_sc_hd__nand2_1
X_05442_ _05678_/A _05678_/B vssd1 vssd1 vccd1 vccd1 _05448_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08161_ _08161_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _08179_/A sky130_fd_sc_hd__nand2_1
X_05373_ _05928_/A _05927_/A vssd1 vssd1 vccd1 vccd1 _05373_/Y sky130_fd_sc_hd__nor2_1
X_08092_ _08092_/A _08128_/A vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07112_ _07112_/A _07112_/B _07112_/C vssd1 vssd1 vccd1 vccd1 _07114_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_70_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07043_ _09022_/C _08688_/A vssd1 vssd1 vccd1 vccd1 _07060_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08994_ _08994_/A _09063_/A _09345_/A vssd1 vssd1 vccd1 vccd1 _09352_/B sky130_fd_sc_hd__nand3_2
X_07945_ _07966_/A _07966_/C vssd1 vssd1 vccd1 vccd1 _07954_/A sky130_fd_sc_hd__nand2_1
X_09615_ _09617_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _09616_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06559__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ _07862_/A _07861_/A _07862_/C vssd1 vssd1 vccd1 vccd1 _07877_/C sky130_fd_sc_hd__a21boi_1
X_06827_ _06827_/A _06828_/A vssd1 vssd1 vccd1 vccd1 _07146_/B sky130_fd_sc_hd__nand2_2
X_09546_ _09572_/A _09572_/C vssd1 vssd1 vccd1 vccd1 _09571_/A sky130_fd_sc_hd__nand2_1
X_06758_ _06758_/A _06758_/B vssd1 vssd1 vccd1 vccd1 _06759_/A sky130_fd_sc_hd__nand2_1
X_09477_ _09477_/A _09477_/B vssd1 vssd1 vccd1 vccd1 _09482_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_78_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05709_ _09199_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _05712_/B sky130_fd_sc_hd__nand2_1
X_08428_ _08428_/A _08428_/B vssd1 vssd1 vccd1 vccd1 _08432_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06689_ _09951_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _06928_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06294__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _08543_/A _08537_/A _08359_/C vssd1 vssd1 vccd1 vccd1 _08363_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ hold121/X vssd1 vssd1 vccd1 vccd1 _10498_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07837__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10252_ hold91/A _10267_/A _10251_/Y vssd1 vssd1 vccd1 vccd1 _10254_/A sky130_fd_sc_hd__a21o_1
X_10183_ hold53/X _10191_/B vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__nand2_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09962__B _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05991_ _06432_/A _06432_/B vssd1 vssd1 vccd1 vccd1 _05996_/C sky130_fd_sc_hd__nand2_1
X_07730_ _07730_/A _07730_/B vssd1 vssd1 vccd1 vccd1 _07816_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07661_ _07666_/B vssd1 vssd1 vccd1 vccd1 _07667_/C sky130_fd_sc_hd__inv_2
X_09400_ _09400_/A vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06612_ _08388_/A _06617_/C vssd1 vssd1 vccd1 vccd1 _06616_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ _07592_/A _07592_/B _07600_/B vssd1 vssd1 vccd1 vccd1 _07600_/A sky130_fd_sc_hd__nand3_1
X_09331_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06543_ _06543_/A _06543_/B vssd1 vssd1 vccd1 vccd1 _06576_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09265_/B sky130_fd_sc_hd__nand2_1
X_06474_ _09684_/B _09313_/D vssd1 vssd1 vccd1 vccd1 _06477_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09193_ _09193_/A _09193_/B _09194_/B vssd1 vssd1 vccd1 vccd1 _09194_/A sky130_fd_sc_hd__nand3_1
X_08213_ _08212_/Y _06438_/A _06438_/B vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05425_ _10051_/B _09313_/D vssd1 vssd1 vccd1 vccd1 _05463_/B sky130_fd_sc_hd__nand2_1
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08144_/Y sky130_fd_sc_hd__nand2_1
X_05356_ _05934_/B _05933_/A vssd1 vssd1 vccd1 vccd1 _05356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06561__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05287_ _05287_/A _05287_/B _05287_/C vssd1 vssd1 vccd1 vccd1 _05293_/B sky130_fd_sc_hd__nand3_1
X_08075_ _10402_/B _08075_/B _08075_/C vssd1 vssd1 vccd1 vccd1 _08086_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10083__B _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07026_ _07345_/B _07345_/C vssd1 vssd1 vccd1 vccd1 _07347_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _08735_/C _08735_/B _08730_/A vssd1 vssd1 vccd1 vccd1 _08978_/B sky130_fd_sc_hd__a21oi_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _07929_/B _07928_/B _07928_/C vssd1 vssd1 vccd1 vccd1 _08040_/B sky130_fd_sc_hd__nand3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07859_ _09392_/C _09777_/A _07859_/C vssd1 vssd1 vccd1 vccd1 _07861_/A sky130_fd_sc_hd__nor3_1
X_09529_ _09529_/A vssd1 vssd1 vccd1 vccd1 _09698_/B sky130_fd_sc_hd__inv_2
XFILLER_0_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05640__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09485__D _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ _10305_/B _10305_/A vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10235_ hold37/X vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08679__A _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ _10166_/A _10166_/B _10166_/C vssd1 vssd1 vccd1 vccd1 _10169_/C sky130_fd_sc_hd__nand3_1
X_10097_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09022__B _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05210_ _05251_/B vssd1 vssd1 vccd1 vccd1 _05216_/B sky130_fd_sc_hd__inv_2
XFILLER_0_32_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06190_ _06190_/A _06190_/B vssd1 vssd1 vccd1 vccd1 _06191_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05278__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _09876_/B _09880_/B _09880_/C vssd1 vssd1 vccd1 vccd1 _09885_/B sky130_fd_sc_hd__nand3b_1
X_08900_ _08900_/A _08900_/B vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__nand2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A vssd1 vssd1 vccd1 vccd1 _08832_/B sky130_fd_sc_hd__inv_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__A _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__nand2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05974_ _05974_/A _05974_/B vssd1 vssd1 vccd1 vccd1 _05974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08693_ _08693_/A vssd1 vssd1 vccd1 vccd1 _08695_/B sky130_fd_sc_hd__inv_2
X_07713_ _07713_/A _10427_/B vssd1 vssd1 vccd1 vccd1 _07716_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07644_ _07642_/Y _07410_/A _07643_/Y vssd1 vssd1 vccd1 vccd1 _07645_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ _07442_/B _07441_/C _07441_/B vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__a21o_1
X_09314_ _09314_/A vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__inv_2
X_06526_ _10026_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _06527_/B sky130_fd_sc_hd__nand2_1
X_09245_ _08986_/B _08983_/A _08991_/A vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06457_ _06457_/A _06457_/B vssd1 vssd1 vccd1 vccd1 _06458_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05408_ _08780_/B _09313_/D vssd1 vssd1 vccd1 vccd1 _05590_/A sky130_fd_sc_hd__nand2_1
X_09176_ _09193_/B _09194_/B vssd1 vssd1 vccd1 vccd1 _09191_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06388_ _06809_/A _06810_/A vssd1 vssd1 vccd1 vccd1 _06388_/Y sky130_fd_sc_hd__nand2_1
X_08127_ _08127_/A _08127_/B _08127_/C vssd1 vssd1 vccd1 vccd1 _08194_/A sky130_fd_sc_hd__nand3_2
X_05339_ _05339_/A _05339_/B _05339_/C vssd1 vssd1 vccd1 vccd1 _05908_/C sky130_fd_sc_hd__nand3_1
X_08058_ _08068_/B _08171_/B vssd1 vssd1 vccd1 vccd1 _08079_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07009_ _07011_/A _07011_/B vssd1 vssd1 vccd1 vccd1 _07010_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10020_ _10020_/A _10020_/B vssd1 vssd1 vccd1 vccd1 _10075_/C sky130_fd_sc_hd__nand2_1
Xoutput69 _10492_/Q vssd1 vssd1 vccd1 vccd1 y_o[12] sky130_fd_sc_hd__buf_12
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07161__A2 _06640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07297__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10218_ _10486_/Q hold35/X vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__or2_1
X_10149_ _10149_/A _10149_/B _10149_/C vssd1 vssd1 vccd1 vccd1 _10154_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08856__B _09141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05690_ _06133_/A _05690_/B vssd1 vssd1 vccd1 vccd1 _06175_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09033__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07360_ _07222_/B _07222_/C _07359_/Y vssd1 vssd1 vccd1 vccd1 _07363_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06311_ _06311_/A _06312_/A vssd1 vssd1 vccd1 vccd1 _06314_/A sky130_fd_sc_hd__nand2_1
X_09030_ _09030_/A vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__inv_2
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07291_ _07104_/Y _07290_/Y _07103_/A vssd1 vssd1 vccd1 vccd1 _07303_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06242_ _06243_/B _06242_/B _06242_/C vssd1 vssd1 vccd1 vccd1 _06782_/C sky130_fd_sc_hd__nand3_1
X_06173_ _06173_/A _06586_/A _06173_/C vssd1 vssd1 vccd1 vccd1 _06179_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _09932_/A vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__inv_2
XFILLER_0_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09863_ _09867_/B vssd1 vssd1 vccd1 vccd1 _09868_/C sky130_fd_sc_hd__inv_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09794_/A _09795_/A vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__nand2_1
X_08814_ _10043_/A _08814_/B vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__nand2_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ input37/X input5/X vssd1 vssd1 vccd1 vccd1 _08746_/C sky130_fd_sc_hd__nand2_1
X_05957_ _06318_/A _06316_/A vssd1 vssd1 vccd1 vccd1 _05957_/Y sky130_fd_sc_hd__nand2_1
X_08676_ _09988_/A input19/X vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__nand2_1
X_05888_ _05888_/A _05888_/B vssd1 vssd1 vccd1 vccd1 _05891_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07627_ _07627_/A _07627_/B vssd1 vssd1 vccd1 vccd1 _07635_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07558_ _07558_/A _07566_/B _07566_/A vssd1 vssd1 vccd1 vccd1 _07809_/A sky130_fd_sc_hd__nand3_2
XANTENNA__06286__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06509_ _08374_/A _08306_/A _06509_/C vssd1 vssd1 vccd1 vccd1 _06513_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09597__B input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ _07489_/A _07489_/B _07489_/C vssd1 vssd1 vccd1 vccd1 _07503_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09228_ _09228_/A vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__inv_2
XFILLER_0_51_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09159_ _09171_/C vssd1 vssd1 vccd1 vccd1 _09172_/C sky130_fd_sc_hd__inv_2
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10003_ _09764_/B _09980_/A input18/X _09762_/Y vssd1 vssd1 vccd1 vccd1 _10004_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_98_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10479__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08692__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06860_ _06864_/A _06861_/A vssd1 vssd1 vccd1 vccd1 _06863_/A sky130_fd_sc_hd__nand2_1
X_05811_ _05814_/A _05814_/B vssd1 vssd1 vccd1 vccd1 _05813_/A sky130_fd_sc_hd__nand2_1
X_06791_ _06792_/A _06791_/B _06791_/C vssd1 vssd1 vccd1 vccd1 _06795_/B sky130_fd_sc_hd__nand3_1
X_08530_ _08796_/B _08531_/C _08531_/B vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05742_ _05742_/A _05742_/B vssd1 vssd1 vccd1 vccd1 _05744_/A sky130_fd_sc_hd__xor2_1
X_08461_ _08757_/A vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__inv_2
X_05673_ _06126_/B _05676_/C vssd1 vssd1 vccd1 vccd1 _05675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07412_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08411_/B _08411_/C vssd1 vssd1 vccd1 vccd1 _08410_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07343_ _07415_/B _07415_/C _07342_/Y vssd1 vssd1 vccd1 vccd1 _07382_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09210__B _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ _07274_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07275_/A sky130_fd_sc_hd__nor2_1
X_09013_ _09014_/B _09014_/A vssd1 vssd1 vccd1 vccd1 _09013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06225_ _09533_/B _09981_/B vssd1 vssd1 vccd1 vccd1 _06353_/A sky130_fd_sc_hd__nand2_1
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06156_ _06158_/A _06158_/B vssd1 vssd1 vccd1 vccd1 _06157_/A sky130_fd_sc_hd__nor2_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06087_ _06087_/A _06087_/B vssd1 vssd1 vccd1 vccd1 _06087_/Y sky130_fd_sc_hd__nor2_1
X_09915_ _09921_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09920_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05466__A _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _09848_/C vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__inv_2
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09777_/A _09777_/B _09777_/C vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__nor3_1
X_06989_ _07000_/A _07001_/B vssd1 vssd1 vccd1 vccd1 _06989_/Y sky130_fd_sc_hd__nor2_1
X_08728_ _09816_/B _09313_/D vssd1 vssd1 vccd1 vccd1 _08729_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_68_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08659_ _08659_/A _08668_/C vssd1 vssd1 vccd1 vccd1 _09189_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10483_ _10495_/CLK hold20/X fanout98/X vssd1 vssd1 vccd1 vccd1 _10483_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09311__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06010_ _09960_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _06012_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07963_/B sky130_fd_sc_hd__inv_2
XANTENNA__09981__A _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09700_ _10023_/B _09700_/B _09700_/C vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06912_ _06912_/A _06912_/B vssd1 vssd1 vccd1 vccd1 _07021_/C sky130_fd_sc_hd__nand2_1
X_07892_ _08049_/B _08049_/A vssd1 vssd1 vccd1 vccd1 _07896_/B sky130_fd_sc_hd__nor2_1
X_09631_ _09629_/X _09631_/B vssd1 vssd1 vccd1 vccd1 _09632_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06843_ _06843_/A _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06999_/C sky130_fd_sc_hd__nand3_1
X_09562_ input46/X _10051_/A _10050_/B _09720_/B vssd1 vssd1 vccd1 vccd1 _09564_/A
+ sky130_fd_sc_hd__and4_1
X_06774_ _06774_/A _06774_/B _06774_/C vssd1 vssd1 vccd1 vccd1 _06775_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08513_ _08512_/B _08513_/B _08513_/C vssd1 vssd1 vccd1 vccd1 _08514_/B sky130_fd_sc_hd__nand3b_1
X_05725_ _05724_/B _06185_/B _05725_/C vssd1 vssd1 vccd1 vccd1 _06185_/A sky130_fd_sc_hd__nand3b_1
X_09493_ _09811_/A _09493_/B vssd1 vssd1 vccd1 vccd1 _09828_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08444_ _08444_/A vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__inv_2
X_05656_ _10026_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _05752_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08375_ _08375_/A _08375_/B vssd1 vssd1 vccd1 vccd1 _08377_/A sky130_fd_sc_hd__nand2_2
X_05587_ _05587_/A vssd1 vssd1 vccd1 vccd1 _05588_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07326_ _10112_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _07330_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07257_ _07253_/Y _07255_/Y _07258_/A vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09023__A2 _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07188_ _07188_/A _07188_/B vssd1 vssd1 vccd1 vccd1 _07188_/Y sky130_fd_sc_hd__nor2_1
X_06208_ _06208_/A _06208_/B _06208_/C vssd1 vssd1 vccd1 vccd1 _06641_/B sky130_fd_sc_hd__nand3_2
X_06139_ _09199_/A vssd1 vssd1 vccd1 vccd1 _10044_/A sky130_fd_sc_hd__inv_2
XANTENNA__08782__A1 _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _09829_/A _09829_/B vssd1 vssd1 vccd1 vccd1 _09830_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06474__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10466_ _10494_/CLK _10466_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10397_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05834__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06490_ _06490_/A _06490_/B vssd1 vssd1 vccd1 vccd1 _06494_/C sky130_fd_sc_hd__nand2_1
X_05510_ _05998_/B vssd1 vssd1 vccd1 vccd1 _05516_/A sky130_fd_sc_hd__inv_2
XANTENNA__06665__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05441_ _05441_/A _05441_/B vssd1 vssd1 vccd1 vccd1 _05448_/A sky130_fd_sc_hd__nand2_1
X_08160_ _08160_/A _08160_/B vssd1 vssd1 vccd1 vccd1 _08161_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05372_ _05929_/C vssd1 vssd1 vccd1 vccd1 _05911_/C sky130_fd_sc_hd__inv_2
X_07111_ _07111_/A _07111_/B vssd1 vssd1 vccd1 vccd1 _07112_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _08091_/A _08091_/B _08091_/C vssd1 vssd1 vccd1 vccd1 _08128_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07042_ _07196_/A _07197_/A vssd1 vssd1 vccd1 vccd1 _07195_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08993_ _08992_/B _09345_/B _08993_/C vssd1 vssd1 vccd1 vccd1 _09345_/A sky130_fd_sc_hd__nand3b_2
X_07944_ _07944_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _07966_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07875_ _08272_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__clkinv_4
X_09614_ _09372_/A _09360_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09616_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__06559__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ _06829_/A _06829_/B vssd1 vssd1 vccd1 vccd1 _06827_/A sky130_fd_sc_hd__nand2_1
X_09545_ _09740_/B _09545_/B vssd1 vssd1 vccd1 vccd1 _09572_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06757_ _06757_/A _06757_/B _06757_/C vssd1 vssd1 vccd1 vccd1 _06854_/B sky130_fd_sc_hd__nand3_1
X_09476_ _09476_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05708_ _09548_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _05712_/A sky130_fd_sc_hd__nand2_1
X_06688_ _06926_/A _06927_/B vssd1 vssd1 vccd1 vccd1 _06930_/C sky130_fd_sc_hd__nand2_1
X_05639_ input39/X vssd1 vssd1 vccd1 vccd1 _09528_/A sky130_fd_sc_hd__clkbuf_8
X_08427_ _08428_/B _08428_/A vssd1 vssd1 vccd1 vccd1 _08674_/A sky130_fd_sc_hd__or2_1
XFILLER_0_65_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06294__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__A _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ _08358_/A vssd1 vssd1 vccd1 vccd1 _08543_/A sky130_fd_sc_hd__inv_2
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08289_ _09227_/A _10044_/D _08289_/C vssd1 vssd1 vccd1 vccd1 _08290_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07309_ _09227_/A _09392_/C _07307_/C vssd1 vssd1 vccd1 vccd1 _07310_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10320_ hold120/X _10325_/A vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__and2_1
XFILLER_0_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10251_ hold40/A _10241_/Y _10243_/B vssd1 vssd1 vccd1 vccd1 _10251_/Y sky130_fd_sc_hd__o21ai_1
X_10182_ hold85/X hold52/X vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05654__A input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ _10449_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10475_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05990_ _05990_/A _05990_/B vssd1 vssd1 vccd1 vccd1 _05996_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07660_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__nand2_1
X_06611_ _06618_/C vssd1 vssd1 vccd1 vccd1 _06615_/B sky130_fd_sc_hd__inv_2
X_07591_ _07591_/A _07591_/B vssd1 vssd1 vccd1 vccd1 _07593_/A sky130_fd_sc_hd__nand2_1
X_09330_ _09320_/Y _09330_/B _09330_/C vssd1 vssd1 vccd1 vccd1 _09335_/B sky130_fd_sc_hd__nand3b_1
X_06542_ _06544_/A vssd1 vssd1 vccd1 vccd1 _06543_/B sky130_fd_sc_hd__inv_2
X_09261_ _09265_/A _09265_/C vssd1 vssd1 vccd1 vccd1 _09264_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08212_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08212_/Y sky130_fd_sc_hd__inv_2
X_06473_ _06517_/A _06518_/A vssd1 vssd1 vccd1 vccd1 _06516_/B sky130_fd_sc_hd__nand2_1
X_09192_ _10448_/B vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__inv_2
XFILLER_0_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05424_ _09022_/C vssd1 vssd1 vccd1 vccd1 _10051_/B sky130_fd_sc_hd__clkbuf_8
X_08143_ _09890_/D _09751_/A _08142_/C vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05355_ _05935_/C vssd1 vssd1 vccd1 vccd1 _05937_/B sky130_fd_sc_hd__inv_2
X_08074_ _08074_/A vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__inv_2
XANTENNA__05739__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07025_ _07025_/A _07025_/B _07025_/C vssd1 vssd1 vccd1 vccd1 _07345_/C sky130_fd_sc_hd__nand3_1
X_05286_ _05568_/A _05286_/B _05286_/C vssd1 vssd1 vccd1 vccd1 _05287_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _08979_/B _08979_/C vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__nand2_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _07927_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _07929_/B sky130_fd_sc_hd__nand2_1
X_07858_ _08866_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _07859_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07789_ _07789_/A _07790_/B _07789_/C vssd1 vssd1 vccd1 vccd1 _07807_/B sky130_fd_sc_hd__nand3_1
X_06809_ _06809_/A _06809_/B vssd1 vssd1 vccd1 vccd1 _06813_/B sky130_fd_sc_hd__nand2_1
X_09528_ _09528_/A _09685_/A _10026_/B _09684_/B vssd1 vssd1 vccd1 vccd1 _09529_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09459_ _09258_/B _09986_/A input19/X _09256_/X vssd1 vssd1 vccd1 vccd1 _09461_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10303_ _10267_/Y _10299_/Y _10268_/Y _10302_/X vssd1 vssd1 vccd1 vccd1 _10305_/A
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10234_ _10234_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _10250_/B sky130_fd_sc_hd__nor2_1
X_10165_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10169_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08679__B input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10096_ _10098_/A vssd1 vssd1 vccd1 vccd1 _10097_/B sky130_fd_sc_hd__inv_2
XFILLER_0_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09022__C _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05278__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07774__A _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ _08830_/A _08831_/A vssd1 vssd1 vccd1 vccd1 _08833_/A sky130_fd_sc_hd__nand2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08761_/A _08761_/B _09049_/A vssd1 vssd1 vccd1 vccd1 _08765_/C sky130_fd_sc_hd__nand3_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05973_ _06205_/A _06205_/B vssd1 vssd1 vccd1 vccd1 _06394_/B sky130_fd_sc_hd__xor2_2
X_08692_ _09980_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _08693_/A sky130_fd_sc_hd__nand2_1
X_07712_ _10418_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10427_/B sky130_fd_sc_hd__nor2_1
X_07643_ _07643_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07643_/Y sky130_fd_sc_hd__nor2_1
X_09313_ _09963_/B _09962_/B _09485_/C _09313_/D vssd1 vssd1 vccd1 vccd1 _09314_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07574_ _07725_/B _07728_/B vssd1 vssd1 vccd1 vccd1 _07574_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06525_ _08361_/B _06528_/C vssd1 vssd1 vccd1 vccd1 _06527_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09244_ _09581_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _09641_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06456_ _06459_/B _06459_/C vssd1 vssd1 vccd1 vccd1 _06458_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05407_ input34/X vssd1 vssd1 vccd1 vccd1 _09313_/D sky130_fd_sc_hd__buf_6
X_09175_ _09430_/A _09175_/B _09175_/C vssd1 vssd1 vccd1 vccd1 _09194_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08126_ _08164_/B vssd1 vssd1 vccd1 vccd1 _08127_/A sky130_fd_sc_hd__inv_2
XFILLER_0_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06387_ _06653_/B _06385_/Y _06386_/Y vssd1 vssd1 vccd1 vccd1 _06810_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__05469__A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05338_ _05338_/A _05338_/B _05338_/C vssd1 vssd1 vccd1 vccd1 _05339_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05269_ _05568_/B _05568_/A vssd1 vssd1 vccd1 vccd1 _05284_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08057_ _08060_/B _08065_/B vssd1 vssd1 vccd1 vccd1 _08068_/B sky130_fd_sc_hd__nand2_1
X_07008_ _07008_/A _07008_/B _07008_/C vssd1 vssd1 vccd1 vccd1 _07011_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08959_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07859__A _09392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10217_ hold79/X vssd1 vssd1 vccd1 vccd1 _10485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10148_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10154_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06003__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ _10079_/A _10079_/B vssd1 vssd1 vccd1 vccd1 _10149_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05842__A _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09033__B _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07290_ _07292_/C vssd1 vssd1 vccd1 vccd1 _07290_/Y sky130_fd_sc_hd__inv_2
X_06310_ _06302_/A _06305_/A _06716_/B vssd1 vssd1 vccd1 vccd1 _06312_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06241_ _06660_/B _06661_/B vssd1 vssd1 vccd1 vccd1 _06242_/C sky130_fd_sc_hd__nand2_1
X_06172_ _06172_/A _06172_/B vssd1 vssd1 vccd1 vccd1 _06179_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09931_ _09931_/A _09931_/B vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09862_ _09563_/X _09565_/A _09564_/A vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__a21oi_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09793_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__nand2_1
X_08813_ _09028_/B _08816_/C vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__nand2_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ input6/X vssd1 vssd1 vccd1 vccd1 _09686_/D sky130_fd_sc_hd__inv_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05956_ _06330_/B _05954_/Y _05955_/Y vssd1 vssd1 vccd1 vccd1 _06316_/A sky130_fd_sc_hd__a21oi_1
X_08675_ _09987_/A input18/X vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__nand2_1
X_05887_ _05887_/A vssd1 vssd1 vccd1 vccd1 _05888_/A sky130_fd_sc_hd__inv_2
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07626_ _07628_/B _07628_/C vssd1 vssd1 vccd1 vccd1 _07627_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07557_ _07556_/A _07556_/B _07556_/C vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06508_ _08374_/B _06508_/B vssd1 vssd1 vccd1 vccd1 _06513_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09597__C _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07488_ _07488_/A _07488_/B vssd1 vssd1 vccd1 vccd1 _07503_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09227_ _09227_/A _10027_/D _09227_/C vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06439_ _06439_/A _08212_/A vssd1 vssd1 vccd1 vccd1 _06467_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09158_ _09161_/B _09162_/B _09162_/C vssd1 vssd1 vccd1 vccd1 _09171_/A sky130_fd_sc_hd__nand3_1
X_09089_ _09089_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09090_/A sky130_fd_sc_hd__nand2_1
X_08109_ _08109_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _08109_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10002_ _10002_/A _10002_/B vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08692__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05810_ _06298_/A _06214_/C _06298_/B vssd1 vssd1 vccd1 vccd1 _06213_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06790_ _06841_/A _06842_/A vssd1 vssd1 vccd1 vccd1 _06834_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05741_ _05741_/A _05702_/Y vssd1 vssd1 vccd1 vccd1 _05742_/B sky130_fd_sc_hd__nor2b_1
XFILLER_0_77_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08460_ _08237_/A _08236_/B _08236_/A vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__a21boi_2
X_05672_ _05672_/A _05672_/B vssd1 vssd1 vccd1 vccd1 _05676_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08391_ _08391_/A _08638_/A _08391_/C vssd1 vssd1 vccd1 vccd1 _08411_/C sky130_fd_sc_hd__nand3_1
X_07411_ _07411_/A _07411_/B _07528_/A vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__nand3_1
X_07342_ _07417_/A _07416_/A vssd1 vssd1 vccd1 vccd1 _07342_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09283__B1 _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09210__C _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ _07274_/A _07274_/B _07217_/A vssd1 vssd1 vccd1 vccd1 _07283_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09012_ _09217_/A _09018_/C vssd1 vssd1 vccd1 vccd1 _09017_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06224_ _06366_/B _06366_/C vssd1 vssd1 vccd1 vccd1 _06365_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06155_ input46/X _08862_/B vssd1 vssd1 vccd1 vccd1 _06158_/B sky130_fd_sc_hd__nand2_1
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__B _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06086_ _06511_/A _06091_/C vssd1 vssd1 vccd1 vccd1 _06579_/B sky130_fd_sc_hd__nand2_1
X_09914_ _10156_/A _10141_/A _09914_/C vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05466__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _09845_/A _09845_/B vssd1 vssd1 vccd1 vccd1 _09848_/C sky130_fd_sc_hd__nand2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09999_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09777_/C sky130_fd_sc_hd__nand2_1
X_06988_ _07004_/C vssd1 vssd1 vccd1 vccd1 _07003_/B sky130_fd_sc_hd__inv_2
X_05939_ _09496_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _06340_/B sky130_fd_sc_hd__nand2_1
X_08727_ input9/X vssd1 vssd1 vccd1 vccd1 _08729_/A sky130_fd_sc_hd__inv_2
XANTENNA__09889__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ _08663_/A _08664_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08668_/C sky130_fd_sc_hd__nand3_2
X_07609_ _07609_/A _07609_/B vssd1 vssd1 vccd1 vccd1 _07611_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08589_ _08589_/A _08589_/B vssd1 vssd1 vccd1 vccd1 _08591_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10482_ _10494_/CLK _10482_/D fanout98/X vssd1 vssd1 vccd1 vccd1 _10482_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05657__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09311__B _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07960_ _08862_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _07961_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09981__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ _06910_/B _06911_/B _06911_/C vssd1 vssd1 vccd1 vccd1 _06912_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_4_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07891_ _08048_/B _08048_/C vssd1 vssd1 vccd1 vccd1 _08049_/A sky130_fd_sc_hd__nand2_1
X_09630_ input52/X _10112_/B input53/X _10111_/B vssd1 vssd1 vccd1 vccd1 _09631_/B
+ sky130_fd_sc_hd__a22o_1
X_06842_ _06842_/A _06842_/B _06842_/C vssd1 vssd1 vccd1 vccd1 _06843_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06398__A _06820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09561_ _09561_/A vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__inv_2
X_06773_ _06773_/A _06773_/B vssd1 vssd1 vccd1 vccd1 _06775_/A sky130_fd_sc_hd__nand2_1
X_08512_ _08512_/A _08512_/B vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__nand2_1
X_05724_ _05724_/A _05724_/B vssd1 vssd1 vccd1 vccd1 _05726_/A sky130_fd_sc_hd__nand2_1
X_09492_ _09492_/A _09492_/B vssd1 vssd1 vccd1 vccd1 _09493_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08443_ _08443_/A _08444_/A vssd1 vssd1 vccd1 vccd1 _08446_/A sky130_fd_sc_hd__nand2_1
X_05655_ _08337_/B vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08374_ _08374_/A _08374_/B vssd1 vssd1 vccd1 vccd1 _08375_/B sky130_fd_sc_hd__or2_1
XFILLER_0_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05586_ _05586_/A _05587_/A vssd1 vssd1 vccd1 vccd1 _05610_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07325_ _08862_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _07330_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07256_ _09560_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _07258_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06207_ _06207_/A vssd1 vssd1 vccd1 vccd1 _06208_/C sky130_fd_sc_hd__inv_2
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07187_ _07187_/A vssd1 vssd1 vccd1 vccd1 _07241_/B sky130_fd_sc_hd__inv_2
X_06138_ _06137_/Y _09199_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _06146_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__05477__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06069_ _06484_/A vssd1 vssd1 vccd1 vccd1 _06072_/A sky130_fd_sc_hd__inv_2
XANTENNA__08788__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ _09828_/A _09495_/B vssd1 vssd1 vccd1 vccd1 _09829_/B sky130_fd_sc_hd__or2b_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09768_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05940__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10465_ _10495_/CLK _10465_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10396_ _10396_/A vssd1 vssd1 vccd1 vccd1 _10460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05387__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05834__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06665__B _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05440_ _05678_/B vssd1 vssd1 vccd1 vccd1 _05441_/B sky130_fd_sc_hd__inv_2
XFILLER_0_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05371_ _05371_/A _05371_/B vssd1 vssd1 vccd1 vccd1 _05929_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_27_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ _07110_/A _07110_/B vssd1 vssd1 vccd1 vccd1 _07112_/A sky130_fd_sc_hd__nand2_1
X_08090_ _08120_/B _08120_/A vssd1 vssd1 vccd1 vccd1 _08091_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07041_ _07181_/C _07181_/B _07040_/Y vssd1 vssd1 vccd1 vccd1 _07197_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05297__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ _08992_/A _08992_/B vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07943_ _07944_/B _07944_/A vssd1 vssd1 vccd1 vccd1 _07966_/A sky130_fd_sc_hd__or2_1
X_07874_ _10126_/B vssd1 vssd1 vccd1 vccd1 _09392_/D sky130_fd_sc_hd__inv_2
X_09613_ _09615_/B _09617_/A vssd1 vssd1 vccd1 vccd1 _09613_/Y sky130_fd_sc_hd__nor2_1
X_06825_ _06825_/A _06825_/B vssd1 vssd1 vccd1 vccd1 _06829_/B sky130_fd_sc_hd__nand2_1
X_09544_ _09740_/B _09740_/A vssd1 vssd1 vccd1 vccd1 _09572_/A sky130_fd_sc_hd__nand2b_1
X_06756_ _06758_/B _06756_/B vssd1 vssd1 vccd1 vccd1 _06757_/B sky130_fd_sc_hd__nand2_1
X_09475_ _09477_/B _09476_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__nand3b_2
X_05707_ _05702_/Y _05705_/Y _05741_/A vssd1 vssd1 vccd1 vccd1 _05720_/B sky130_fd_sc_hd__a21oi_1
X_06687_ _09560_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _06927_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ _08674_/B _08426_/B vssd1 vssd1 vccd1 vccd1 _08428_/A sky130_fd_sc_hd__nand2_1
X_05638_ _05643_/A vssd1 vssd1 vccd1 vccd1 _05642_/A sky130_fd_sc_hd__inv_2
XFILLER_0_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08357_ _08543_/B _08358_/A vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05569_ _05284_/B _05284_/C _05568_/Y vssd1 vssd1 vccd1 vccd1 _05981_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_34_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08288_ _09962_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _08289_/C sky130_fd_sc_hd__nand2_1
X_07308_ _07308_/A vssd1 vssd1 vccd1 vccd1 _07380_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07239_ _07241_/C vssd1 vssd1 vccd1 vccd1 _07239_/Y sky130_fd_sc_hd__inv_2
X_10250_ _10250_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__and2_1
X_10181_ _10181_/A _10181_/B vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10448_ _10448_/A _10448_/B vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__nand2_1
X_10379_ hold3/X _10379_/B vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__xor2_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06610_ _08657_/C _06610_/B vssd1 vssd1 vccd1 vccd1 _06618_/C sky130_fd_sc_hd__nand2_2
X_07590_ _07592_/A vssd1 vssd1 vccd1 vccd1 _07591_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06541_ _06130_/A _06127_/A _06127_/B vssd1 vssd1 vccd1 vccd1 _06544_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05580__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ _09260_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _09265_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09987__A _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06472_ _06405_/Y _06048_/B _06406_/Y vssd1 vssd1 vccd1 vccd1 _06518_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _10437_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_28_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05423_ _10052_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _05462_/B sky130_fd_sc_hd__nand2_1
X_09191_ _09191_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09191_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ _09890_/D _09751_/A _08142_/C vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__or3_1
X_05354_ _09496_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _05935_/C sky130_fd_sc_hd__nand2_1
X_05285_ _05568_/B _05285_/B vssd1 vssd1 vccd1 vccd1 _05287_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ _08073_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _08074_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05739__B _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07024_ _07024_/A _07024_/B _07024_/C vssd1 vssd1 vccd1 vccd1 _07025_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08975_ _08975_/A _08975_/B vssd1 vssd1 vccd1 vccd1 _08979_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09227__A _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05755__A _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _07926_/A _07926_/B vssd1 vssd1 vccd1 vccd1 _07927_/B sky130_fd_sc_hd__nand2_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__buf_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10507__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ _08248_/B vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__inv_2
XFILLER_0_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06808_ _06810_/A vssd1 vssd1 vccd1 vccd1 _06809_/B sky130_fd_sc_hd__inv_2
X_07788_ _07788_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__nand2_1
X_09527_ _09326_/B _09960_/A _10026_/B _09324_/X vssd1 vssd1 vccd1 vccd1 _09702_/A
+ sky130_fd_sc_hd__a31o_1
X_06739_ _06739_/A _06739_/B _06739_/C vssd1 vssd1 vccd1 vccd1 _06747_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09458_ _09458_/A _09458_/B vssd1 vssd1 vccd1 vccd1 _09461_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09389_ _09397_/A _09397_/B vssd1 vssd1 vccd1 vccd1 _09396_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08409_ _08644_/B _08408_/Y vssd1 vssd1 vccd1 vccd1 _08410_/B sky130_fd_sc_hd__nor2b_1
XFILLER_0_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _10300_/X _10298_/Y _10299_/Y hold104/A _10301_/X vssd1 vssd1 vccd1 vccd1
+ _10302_/X sky130_fd_sc_hd__o221a_1
X_10233_ hold40/X vssd1 vssd1 vccd1 vccd1 _10234_/B sky130_fd_sc_hd__inv_2
XFILLER_0_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10164_ _10166_/B vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__inv_2
X_10095_ _09729_/C _09729_/B _09718_/Y vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09022__D _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08216__A _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07774__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08760_ _09049_/B _08760_/B vssd1 vssd1 vccd1 vccd1 _08765_/B sky130_fd_sc_hd__nand2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05972_ _05895_/A _05894_/A _05899_/B vssd1 vssd1 vccd1 vccd1 _06205_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08691_ _08691_/A _08691_/B vssd1 vssd1 vccd1 vccd1 _08695_/C sky130_fd_sc_hd__nand2_1
X_07711_ _10429_/B _07711_/B vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__nand2_1
X_07642_ _07643_/B _07643_/A vssd1 vssd1 vccd1 vccd1 _07642_/Y sky130_fd_sc_hd__nand2_1
X_09312_ _09312_/A vssd1 vssd1 vccd1 vccd1 _09318_/B sky130_fd_sc_hd__inv_2
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07573_ _07573_/A _07573_/B vssd1 vssd1 vccd1 vccd1 _07728_/B sky130_fd_sc_hd__nand2_2
X_06524_ _06524_/A _06524_/B vssd1 vssd1 vccd1 vccd1 _06528_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09243_ _09243_/A _09243_/B _09243_/C vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06455_ _08300_/A _06455_/B _08260_/A vssd1 vssd1 vccd1 vccd1 _06459_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _09178_/B _09178_/A vssd1 vssd1 vccd1 vccd1 _09175_/B sky130_fd_sc_hd__nor2_1
X_06386_ _06646_/A _06651_/A vssd1 vssd1 vccd1 vccd1 _06386_/Y sky130_fd_sc_hd__nor2_1
X_05406_ _05395_/A _05398_/A _05405_/Y vssd1 vssd1 vccd1 vccd1 _05732_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08125_ _08125_/A _08133_/A vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05337_ _05337_/A _05337_/B vssd1 vssd1 vccd1 vccd1 _05339_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05469__B _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05268_ _05219_/C _05219_/B _05251_/Y vssd1 vssd1 vccd1 vccd1 _05568_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ _08056_/A _08056_/B vssd1 vssd1 vccd1 vccd1 _08060_/B sky130_fd_sc_hd__nand2_1
X_07007_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07011_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08958_ _08959_/B _08959_/A vssd1 vssd1 vccd1 vccd1 _08958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08889_ _08857_/Y _08589_/B _08858_/Y vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__a21oi_1
X_07909_ _07909_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _08071_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07859__B _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07875__A _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10216_ hold78/X _10221_/A vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__and2_1
X_10147_ _10149_/B vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__inv_2
XFILLER_0_100_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06003__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _10078_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10079_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05842__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_06240_ _06662_/C vssd1 vssd1 vccd1 vccd1 _06242_/B sky130_fd_sc_hd__inv_2
XFILLER_0_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06171_ _06173_/A vssd1 vssd1 vccd1 vccd1 _06172_/B sky130_fd_sc_hd__inv_2
X_09930_ _09936_/A _09936_/C vssd1 vssd1 vccd1 vccd1 _09934_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09861_ _10091_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__nand2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09792_/A _09792_/B _09792_/C vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08812_ _10044_/A _08811_/B _08811_/C vssd1 vssd1 vccd1 vccd1 _08816_/C sky130_fd_sc_hd__o21ai_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08743_/A vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__inv_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05955_ _06328_/A _06327_/A vssd1 vssd1 vccd1 vccd1 _05955_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08674_ _08674_/A _08674_/B vssd1 vssd1 vccd1 vccd1 _08683_/A sky130_fd_sc_hd__nand2_1
X_05886_ _05887_/A _05886_/B _05886_/C vssd1 vssd1 vccd1 vccd1 _05891_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_88_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _07625_/A _07625_/B vssd1 vssd1 vccd1 vccd1 _07628_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07556_ _07556_/A _07556_/B _07556_/C vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06507_ _08374_/A vssd1 vssd1 vccd1 vccd1 _06508_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09597__D _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09226_ _09496_/B vssd1 vssd1 vccd1 vccd1 _10027_/D sky130_fd_sc_hd__inv_2
XFILLER_0_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07487_ _07489_/A _07489_/C vssd1 vssd1 vccd1 vccd1 _07488_/A sky130_fd_sc_hd__nand2_1
X_06438_ _06438_/A _06438_/B vssd1 vssd1 vccd1 vccd1 _06439_/A sky130_fd_sc_hd__nand2_1
X_09157_ _09146_/Y _08634_/B _09147_/Y vssd1 vssd1 vccd1 vccd1 _09161_/B sky130_fd_sc_hd__a21o_1
X_06369_ _06368_/B _06369_/B _06369_/C vssd1 vssd1 vccd1 vccd1 _06370_/B sky130_fd_sc_hd__nand3b_1
X_09088_ _09090_/B _09089_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ _08157_/B _08108_/B vssd1 vssd1 vccd1 vccd1 _08138_/A sky130_fd_sc_hd__and2_1
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08039_ _08039_/A _08088_/B _08088_/A vssd1 vssd1 vccd1 vccd1 _08127_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10001_ _10001_/A _10001_/B vssd1 vssd1 vccd1 vccd1 _10002_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10114__B1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05740_ _05740_/A vssd1 vssd1 vccd1 vccd1 _05821_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05671_ _05671_/A _05671_/B vssd1 vssd1 vccd1 vccd1 _06126_/B sky130_fd_sc_hd__nand2_1
X_08390_ _08390_/A vssd1 vssd1 vccd1 vccd1 _08638_/A sky130_fd_sc_hd__inv_2
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07410_ _07410_/A vssd1 vssd1 vccd1 vccd1 _07528_/A sky130_fd_sc_hd__inv_2
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07341_ _07418_/C vssd1 vssd1 vccd1 vccd1 _07415_/C sky130_fd_sc_hd__inv_2
XANTENNA__09283__B2 _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A1 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09210__D _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ _07272_/A vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__inv_2
X_09011_ _09011_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _09018_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06223_ _06223_/A _06223_/B _06223_/C vssd1 vssd1 vccd1 vccd1 _06366_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_26_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06154_ _10051_/A input1/X vssd1 vssd1 vccd1 vccd1 _06158_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09219__B _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06085_ _06085_/A _06085_/B _06085_/C vssd1 vssd1 vccd1 vccd1 _06091_/C sky130_fd_sc_hd__nand3_1
X_09913_ _09913_/A vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__inv_2
X_09844_ _10078_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05763__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ _09998_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _09782_/B sky130_fd_sc_hd__nand2_1
X_06987_ _06987_/A _06992_/A vssd1 vssd1 vccd1 vccd1 _07004_/C sky130_fd_sc_hd__nand2_1
X_08726_ _08726_/A _08769_/B _08901_/A vssd1 vssd1 vccd1 vccd1 _08900_/B sky130_fd_sc_hd__nand3_2
X_05938_ _06334_/B _06334_/C vssd1 vssd1 vccd1 vccd1 _06333_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09889__B _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ _08657_/A _08657_/B _08657_/C vssd1 vssd1 vccd1 vccd1 _08663_/B sky130_fd_sc_hd__nand3_1
X_05869_ _05871_/A _05871_/C vssd1 vssd1 vccd1 vccd1 _05870_/A sky130_fd_sc_hd__nand2_1
X_07608_ _07606_/Y _07803_/B _07607_/Y vssd1 vssd1 vccd1 vccd1 _07899_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08588_ _08368_/A _08366_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08589_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07539_ _07539_/A _07539_/B _07539_/C vssd1 vssd1 vccd1 vccd1 _07545_/A sky130_fd_sc_hd__nand3_1
X_09209_ _10050_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _09213_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10481_ _10494_/CLK _10481_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__05657__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__B _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06910_ _06910_/A _06910_/B vssd1 vssd1 vccd1 vccd1 _06912_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07890_ _07889_/B _07890_/B _07890_/C vssd1 vssd1 vccd1 vccd1 _08048_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06841_ _06841_/A _06841_/B vssd1 vssd1 vccd1 vccd1 _06843_/A sky130_fd_sc_hd__nand2_1
X_09560_ _10050_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _09561_/A sky130_fd_sc_hd__nand2_1
X_06772_ _06774_/A _06774_/C vssd1 vssd1 vccd1 vccd1 _06773_/A sky130_fd_sc_hd__nand2_1
X_09491_ _09492_/A _09490_/Y vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05723_ input46/X _08866_/B vssd1 vssd1 vccd1 vccd1 _05724_/B sky130_fd_sc_hd__nand2_1
X_08511_ _08511_/A _08511_/B vssd1 vssd1 vccd1 vccd1 _08512_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ _08442_/A _08714_/A vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__nand2_1
X_05654_ input23/X vssd1 vssd1 vccd1 vccd1 _08337_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _08378_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08604_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05585_ input35/X _08780_/B vssd1 vssd1 vccd1 vccd1 _05587_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07324_ _07448_/A _07448_/C vssd1 vssd1 vccd1 vccd1 _07447_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07255_ _07259_/C vssd1 vssd1 vccd1 vccd1 _07255_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05758__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06206_ _06206_/A _06207_/A vssd1 vssd1 vccd1 vccd1 _06641_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07186_ _10051_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _07187_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06137_ _09548_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _06137_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05477__B _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06068_ _09533_/B _09313_/D vssd1 vssd1 vccd1 vccd1 _06484_/A sky130_fd_sc_hd__nand2_1
X_09827_ _09831_/B _09831_/C vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__nand2_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ _09758_/A vssd1 vssd1 vccd1 vccd1 _09993_/B sky130_fd_sc_hd__inv_2
X_08709_ _08932_/B _08712_/C vssd1 vssd1 vccd1 vccd1 _08711_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09689_ _09690_/B _09690_/A vssd1 vssd1 vccd1 vccd1 _10034_/A sky130_fd_sc_hd__or2_1
XFILLER_0_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05940__B _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07213__A _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10464_ _10494_/CLK _10464_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__05387__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ _10395_/A _10397_/A vssd1 vssd1 vccd1 vccd1 _10396_/A sky130_fd_sc_hd__and2_1
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05370_ _05370_/A _05370_/B _05370_/C vssd1 vssd1 vccd1 vccd1 _05371_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07040_ _07178_/B _07177_/A vssd1 vssd1 vccd1 vccd1 _07040_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__05578__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05297__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08991_ _08991_/A _08991_/B vssd1 vssd1 vccd1 vccd1 _08992_/B sky130_fd_sc_hd__nand2_1
X_07942_ _07833_/Y _07942_/B vssd1 vssd1 vccd1 vccd1 _07944_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07873_ _07880_/B _07880_/A vssd1 vssd1 vccd1 vccd1 _07928_/B sky130_fd_sc_hd__nand2_1
X_09612_ _09612_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09617_/A sky130_fd_sc_hd__nand2_1
X_06824_ _06838_/B _06801_/Y _06802_/Y vssd1 vssd1 vccd1 vccd1 _06825_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09543_ _09545_/B vssd1 vssd1 vccd1 vccd1 _09740_/A sky130_fd_sc_hd__inv_2
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06755_ _06755_/A vssd1 vssd1 vccd1 vccd1 _06758_/B sky130_fd_sc_hd__inv_2
X_09474_ _09474_/A _09474_/B _09770_/A vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05706_ _05706_/A _05706_/B vssd1 vssd1 vccd1 vccd1 _05741_/A sky130_fd_sc_hd__nor2_1
X_06686_ _10083_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _06926_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ _08425_/A _08425_/B vssd1 vssd1 vccd1 vccd1 _08426_/B sky130_fd_sc_hd__nand2_1
X_05637_ _09685_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _05643_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _08356_/A _08356_/B vssd1 vssd1 vccd1 vccd1 _08358_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07307_ _09227_/A _09392_/C _07307_/C vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__nor3_1
X_05568_ _05568_/A _05568_/B vssd1 vssd1 vccd1 vccd1 _05568_/Y sky130_fd_sc_hd__nor2_1
X_08287_ _09533_/B vssd1 vssd1 vccd1 vccd1 _10044_/D sky130_fd_sc_hd__inv_2
XFILLER_0_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05499_ _05499_/A vssd1 vssd1 vccd1 vccd1 _05499_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07238_ _07466_/B _07466_/C vssd1 vssd1 vccd1 vccd1 _07468_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07169_ _07165_/Y _07169_/B _07169_/C vssd1 vssd1 vccd1 vccd1 _07173_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10180_ hold52/X vssd1 vssd1 vccd1 vccd1 _10181_/B sky130_fd_sc_hd__inv_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10447_ _10447_/A vssd1 vssd1 vccd1 vccd1 _10474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10378_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10379_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10506__RESET_B fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06540_ _08365_/A _06544_/C vssd1 vssd1 vccd1 vccd1 _06543_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05580__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06471_ _08268_/A _06518_/C vssd1 vssd1 vccd1 vccd1 _06517_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10459__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05422_ _08780_/B vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__buf_8
X_08210_ _08210_/A _10407_/B _08210_/C vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__nand3_1
X_09190_ _09190_/A _09190_/B vssd1 vssd1 vccd1 vccd1 _09190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08141_ _10111_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _08142_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05353_ _05934_/B _05933_/A vssd1 vssd1 vccd1 vccd1 _05937_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05284_ _05502_/B _05284_/B _05284_/C vssd1 vssd1 vccd1 vccd1 _05502_/A sky130_fd_sc_hd__nand3_1
X_08072_ _08072_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08073_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07023_ _07023_/A _07023_/B vssd1 vssd1 vccd1 vccd1 _07025_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05739__C _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ _08975_/B _08975_/A vssd1 vssd1 vccd1 vccd1 _08979_/B sky130_fd_sc_hd__or2_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _07925_/A _07925_/B _07925_/C vssd1 vssd1 vccd1 vccd1 _07926_/B sky130_fd_sc_hd__nand3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ _07862_/A _07862_/C vssd1 vssd1 vccd1 vccd1 _07860_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06867__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ _06804_/Y _06828_/A _06806_/Y vssd1 vssd1 vccd1 vccd1 _07148_/B sky130_fd_sc_hd__a21oi_2
X_07787_ _10111_/B _09485_/C _10126_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _07788_/B
+ sky130_fd_sc_hd__a22o_1
X_09526_ _09526_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09541_/A sky130_fd_sc_hd__nor2_1
X_06738_ _06831_/B _06831_/C vssd1 vssd1 vccd1 vccd1 _06836_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09457_ _09458_/B _09458_/A vssd1 vssd1 vccd1 vccd1 _09461_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08408_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08408_/Y sky130_fd_sc_hd__nand2_1
X_06669_ _06769_/A _06770_/A vssd1 vssd1 vccd1 vccd1 _06669_/Y sky130_fd_sc_hd__nor2_1
X_09388_ _09388_/A _09388_/B _09647_/A vssd1 vssd1 vccd1 vccd1 _09397_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08339_ _09083_/A _10113_/D _08338_/C vssd1 vssd1 vccd1 vccd1 _08340_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10301_ hold28/A _10290_/Y hold114/X vssd1 vssd1 vccd1 vccd1 _10301_/X sky130_fd_sc_hd__o21a_1
X_10232_ _10488_/Q hold39/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__nand2_1
X_10163_ _09936_/C _09936_/B _09928_/A vssd1 vssd1 vccd1 vccd1 _10166_/B sky130_fd_sc_hd__a21oi_1
X_10094_ _10098_/B _10098_/C vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08216__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08232__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05856__A _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _07710_/A _07710_/B vssd1 vssd1 vccd1 vccd1 _07711_/B sky130_fd_sc_hd__nand2_1
X_05971_ _05974_/B _05974_/A vssd1 vssd1 vccd1 vccd1 _06394_/C sky130_fd_sc_hd__nand2_1
X_08690_ _08691_/A _08691_/B vssd1 vssd1 vccd1 vccd1 _08933_/B sky130_fd_sc_hd__or2_1
XANTENNA__06687__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _07647_/B _07647_/C vssd1 vssd1 vccd1 vccd1 _07645_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09998__A _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ _07572_/A _07572_/B vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09311_ _09951_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09312_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06523_ _06524_/A _06524_/B vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ _09242_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06454_ _08300_/B _06454_/B vssd1 vssd1 vccd1 vccd1 _06459_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ _09173_/A _09173_/B vssd1 vssd1 vccd1 vccd1 _09178_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06385_ _06651_/A _06646_/A vssd1 vssd1 vccd1 vccd1 _06385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05405_ _05405_/A _05405_/B vssd1 vssd1 vccd1 vccd1 _05405_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ _08124_/A _08128_/A _08128_/B vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05336_ _05903_/B _05903_/C vssd1 vssd1 vccd1 vccd1 _05902_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05267_ _05286_/B _05286_/C vssd1 vssd1 vccd1 vccd1 _05568_/B sky130_fd_sc_hd__nand2_1
X_08055_ _08055_/A _08055_/B vssd1 vssd1 vccd1 vccd1 _08056_/A sky130_fd_sc_hd__nand2_1
X_07006_ _07008_/A vssd1 vssd1 vccd1 vccd1 _07007_/B sky130_fd_sc_hd__inv_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08957_ _09345_/B _08993_/C vssd1 vssd1 vccd1 vccd1 _08992_/A sky130_fd_sc_hd__nand2_1
X_08888_ _08888_/A _09118_/A vssd1 vssd1 vccd1 vccd1 _08890_/A sky130_fd_sc_hd__nand2_1
X_07908_ _07911_/B _07914_/B vssd1 vssd1 vccd1 vccd1 _07909_/A sky130_fd_sc_hd__nand2_1
X_07839_ _09854_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _07841_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09509_ _09511_/C vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__inv_2
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10215_ hold77/X _10215_/B vssd1 vssd1 vccd1 vccd1 _10221_/A sky130_fd_sc_hd__nand2_1
X_10146_ _10146_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__nand2_1
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06170_ _06168_/Y _05619_/A _06169_/Y vssd1 vssd1 vccd1 vccd1 _06173_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__06970__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _09860_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08897__A _09141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _09792_/A _09792_/C _09792_/B vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__a21o_1
X_08811_ _10044_/A _08811_/B _08811_/C vssd1 vssd1 vccd1 vccd1 _09028_/B sky130_fd_sc_hd__or3_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08742_ _09960_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__nand2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05954_ _06327_/A _06328_/A vssd1 vssd1 vccd1 vccd1 _05954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08673_ _08673_/A _08673_/B vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07306__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07624_ _07624_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _07625_/B sky130_fd_sc_hd__nand2_1
X_05885_ _05854_/Y _05962_/B _05884_/Y vssd1 vssd1 vccd1 vccd1 _05894_/A sky130_fd_sc_hd__a21oi_2
X_07555_ _07733_/B _07567_/C _07733_/A vssd1 vssd1 vccd1 vccd1 _07558_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06506_ _06504_/Y _06044_/B _06505_/Y vssd1 vssd1 vccd1 vccd1 _08374_/A sky130_fd_sc_hd__a21oi_2
X_07486_ _07486_/A vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__inv_2
X_09225_ _09525_/A _09231_/B vssd1 vssd1 vccd1 vccd1 _09229_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06437_ _08212_/A _06438_/A _06438_/B vssd1 vssd1 vccd1 vccd1 _06467_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _09430_/A _09175_/C vssd1 vssd1 vccd1 vccd1 _09170_/A sky130_fd_sc_hd__nand2_1
X_06368_ _06368_/A _06368_/B vssd1 vssd1 vccd1 vccd1 _06370_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ _09087_/A _09087_/B _09087_/C vssd1 vssd1 vccd1 vccd1 _09381_/B sky130_fd_sc_hd__nand3_1
X_08107_ _10111_/B _09981_/A _10126_/B _09981_/B vssd1 vssd1 vccd1 vccd1 _08108_/B
+ sky130_fd_sc_hd__a22o_1
X_05319_ _05324_/B vssd1 vssd1 vccd1 vccd1 _05320_/B sky130_fd_sc_hd__inv_2
X_06299_ _06299_/A _06299_/B vssd1 vssd1 vccd1 vccd1 _06300_/B sky130_fd_sc_hd__and2_1
X_08038_ _08038_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08088_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10000_ _10000_/A input18/X vssd1 vssd1 vccd1 vccd1 _10001_/B sky130_fd_sc_hd__nand2_1
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07216__A _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08004__B1 _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10129_ _10129_/A _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_89_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10114__B2 _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05670_ _05672_/B vssd1 vssd1 vccd1 vccd1 _05671_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07340_ _07378_/A _07340_/B vssd1 vssd1 vccd1 vccd1 _07418_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09283__A2 _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09010_ _09010_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09011_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07271_ _07423_/C _07423_/B _07270_/Y vssd1 vssd1 vccd1 vccd1 _07284_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06222_ _06222_/A _06222_/B vssd1 vssd1 vccd1 vccd1 _06223_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06153_ input47/X vssd1 vssd1 vccd1 vccd1 _10051_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ _06084_/A _06084_/B _06084_/C vssd1 vssd1 vccd1 vccd1 _06085_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09912_ _10156_/B _09913_/A vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__nand2_1
X_09843_ _09843_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08420__A _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05763__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _09796_/A _09796_/C vssd1 vssd1 vccd1 vccd1 _09794_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07036__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06986_ _07127_/A _06992_/B _06986_/C vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__nand3b_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _08725_/A _08901_/B _08725_/C vssd1 vssd1 vccd1 vccd1 _08901_/A sky130_fd_sc_hd__nand3_2
X_05937_ _05937_/A _05937_/B _05937_/C vssd1 vssd1 vccd1 vccd1 _06334_/C sky130_fd_sc_hd__nand3_1
XANTENNA__06875__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05868_ _05868_/A _05868_/B vssd1 vssd1 vccd1 vccd1 _05871_/A sky130_fd_sc_hd__nand2_1
X_08656_ _08656_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _08664_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ _08590_/B _08590_/C vssd1 vssd1 vccd1 vccd1 _08589_/A sky130_fd_sc_hd__nand2_1
X_07607_ _07799_/A _07801_/A vssd1 vssd1 vccd1 vccd1 _07607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07538_ _07799_/B _07799_/C vssd1 vssd1 vccd1 vccd1 _07801_/A sky130_fd_sc_hd__nand2_1
X_05799_ _10026_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _06280_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ _07471_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07470_/A sky130_fd_sc_hd__nand2_1
X_09208_ _09208_/A _09594_/A vssd1 vssd1 vccd1 vccd1 _09215_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_63_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10480_ _10494_/CLK _10480_/D fanout98/X vssd1 vssd1 vccd1 vccd1 _10480_/Q sky130_fd_sc_hd__dfrtp_1
X_09139_ _09141_/A vssd1 vssd1 vccd1 vccd1 _09140_/B sky130_fd_sc_hd__inv_2
XFILLER_0_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09982__B1 _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10494_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10492__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06025__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06840_ _07138_/B _07138_/C vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06771_ _06771_/A _06771_/B vssd1 vssd1 vccd1 vccd1 _06774_/A sky130_fd_sc_hd__nand2_1
X_09490_ _09492_/B vssd1 vssd1 vccd1 vccd1 _09490_/Y sky130_fd_sc_hd__inv_2
X_05722_ input1/X vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__clkbuf_8
X_08510_ _08510_/A _08510_/B vssd1 vssd1 vccd1 vccd1 _08511_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08441_ _08714_/B _08441_/B _08441_/C vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__nand3_1
X_05653_ _05665_/B _05665_/A vssd1 vssd1 vccd1 vccd1 _05749_/A sky130_fd_sc_hd__nand2_1
X_08372_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08378_/B sky130_fd_sc_hd__nand2_1
X_05584_ _05588_/A _05588_/C vssd1 vssd1 vccd1 vccd1 _05586_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07323_ _07323_/A _07323_/B _07323_/C vssd1 vssd1 vccd1 vccd1 _07448_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07254_ _07254_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07259_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06205_ _06205_/A _06205_/B vssd1 vssd1 vccd1 vccd1 _06207_/A sky130_fd_sc_hd__nor2_1
XANTENNA__05758__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ _07188_/A _07188_/B vssd1 vssd1 vccd1 vccd1 _07241_/C sky130_fd_sc_hd__nand2_2
X_06136_ _06166_/A _06166_/B vssd1 vssd1 vccd1 vccd1 _06165_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06067_ _06084_/B vssd1 vssd1 vccd1 vccd1 _06083_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09826_ _09826_/A _09975_/A _10063_/A vssd1 vssd1 vccd1 vccd1 _09831_/C sky130_fd_sc_hd__nand3_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09757_ _09759_/B _09759_/A vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__nor2_1
X_06969_ _06992_/B _06986_/C vssd1 vssd1 vccd1 vccd1 _06985_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08708_ _09805_/A _09777_/A _08707_/C vssd1 vssd1 vccd1 vccd1 _08712_/C sky130_fd_sc_hd__o21ai_1
X_09688_ _10034_/B _09688_/B vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08639_ _08637_/Y _08410_/B _08638_/Y vssd1 vssd1 vccd1 vccd1 _09166_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07213__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08325__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10463_ _10495_/CLK _10463_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfrtp_1
X_10394_ _10394_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05859__A _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05578__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08990_ _08989_/B _08990_/B _08990_/C vssd1 vssd1 vccd1 vccd1 _08991_/B sky130_fd_sc_hd__nand3b_1
X_07941_ _07941_/A _07941_/B vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__nand2_1
X_07872_ _07872_/A _07872_/B vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__nand2_1
X_09611_ _09611_/A _09611_/B _09611_/C vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__nand3_1
X_06823_ _06823_/A _06823_/B _06823_/C vssd1 vssd1 vccd1 vccd1 _06829_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09542_ _09542_/A _09542_/B vssd1 vssd1 vccd1 vccd1 _09545_/B sky130_fd_sc_hd__nand2_1
X_06754_ _06758_/A _06755_/A vssd1 vssd1 vccd1 vccd1 _06757_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05705_ _05742_/A vssd1 vssd1 vccd1 vccd1 _05705_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09473_ _09473_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__nand2_1
X_06685_ _08825_/B vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08674_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05636_ input27/X vssd1 vssd1 vccd1 vccd1 _09361_/C sky130_fd_sc_hd__buf_6
X_08355_ _08537_/A _08359_/C vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05567_ _06022_/A _05572_/C vssd1 vssd1 vccd1 vccd1 _05981_/B sky130_fd_sc_hd__nand2_1
X_07306_ _09962_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _07307_/C sky130_fd_sc_hd__nand2_1
X_08286_ _09960_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08532_/A sky130_fd_sc_hd__nand2_1
X_05498_ _05500_/B _05500_/A vssd1 vssd1 vccd1 vccd1 _05499_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07237_ _07237_/A _07237_/B _07237_/C vssd1 vssd1 vccd1 vccd1 _07466_/C sky130_fd_sc_hd__nand3_1
X_07168_ _07170_/A _07171_/A vssd1 vssd1 vccd1 vccd1 _07169_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06119_ _06534_/B _06119_/B _06119_/C vssd1 vssd1 vccd1 vccd1 _06534_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07099_ _09601_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _07104_/A sky130_fd_sc_hd__nand2_1
X_09809_ _09809_/A _09809_/B vssd1 vssd1 vccd1 vccd1 _09814_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10446_ _10446_/A _10448_/A vssd1 vssd1 vccd1 vccd1 _10447_/A sky130_fd_sc_hd__and2_1
X_10377_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__xor2_1
XFILLER_0_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09459__A2 _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06470_ _06517_/B _08268_/A _06518_/C vssd1 vssd1 vccd1 vccd1 _08317_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05421_ _05453_/A _05453_/C vssd1 vssd1 vccd1 vccd1 _05452_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ _10126_/B _09986_/A vssd1 vssd1 vccd1 vccd1 _08140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05352_ _09960_/B _09988_/A vssd1 vssd1 vccd1 vccd1 _05933_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05283_ _05287_/C vssd1 vssd1 vccd1 vccd1 _05284_/C sky130_fd_sc_hd__inv_2
X_08071_ _08071_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08072_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07022_ _07392_/B _07392_/C vssd1 vssd1 vccd1 vccd1 _07391_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05739__D input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08973_ _08973_/A _08973_/B vssd1 vssd1 vccd1 vccd1 _08975_/A sky130_fd_sc_hd__xor2_1
X_07924_ _07924_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07926_/A sky130_fd_sc_hd__nand2_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _07855_/A _07855_/B _07855_/C vssd1 vssd1 vccd1 vccd1 _07862_/C sky130_fd_sc_hd__nand3_1
XANTENNA__06867__B input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07786_ _07817_/A _07816_/A vssd1 vssd1 vccd1 vccd1 _07815_/C sky130_fd_sc_hd__nand2_1
X_06806_ _06823_/A _06825_/A vssd1 vssd1 vccd1 vccd1 _06806_/Y sky130_fd_sc_hd__nor2_1
X_09525_ _09525_/A vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__inv_2
X_06737_ _06737_/A _06737_/B _06737_/C vssd1 vssd1 vccd1 vccd1 _06831_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09456_ _09454_/X _09456_/B vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__nand2b_1
X_06668_ _06773_/B vssd1 vssd1 vccd1 vccd1 _06774_/B sky130_fd_sc_hd__inv_2
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _08408_/B _08408_/A vssd1 vssd1 vccd1 vccd1 _08644_/B sky130_fd_sc_hd__nor2_2
X_05619_ _05619_/A vssd1 vssd1 vccd1 vccd1 _05620_/C sky130_fd_sc_hd__inv_2
X_09387_ _09387_/A vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__inv_2
XFILLER_0_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06599_ _06599_/A _06599_/B vssd1 vssd1 vccd1 vccd1 _06600_/B sky130_fd_sc_hd__nand2_1
X_08338_ _09083_/A _10113_/D _08338_/C vssd1 vssd1 vccd1 vccd1 _08341_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08269_ _08313_/B vssd1 vssd1 vccd1 vccd1 _08314_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10300_ hold32/A hold81/A _10277_/B vssd1 vssd1 vccd1 vccd1 _10300_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10231_ _10488_/Q hold39/X vssd1 vssd1 vccd1 vccd1 _10234_/A sky130_fd_sc_hd__nor2_1
X_10162_ _10166_/A _10166_/C vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__nand2_1
X_10093_ _10092_/B _10093_/B _10093_/C vssd1 vssd1 vccd1 vccd1 _10098_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08232__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ _10429_/A _10429_/B _10429_/C vssd1 vssd1 vccd1 vccd1 _10431_/A sky130_fd_sc_hd__nand3_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06033__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05970_ _06211_/B _06211_/C _05969_/Y vssd1 vssd1 vccd1 vccd1 _05974_/A sky130_fd_sc_hd__a21oi_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06687__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ _07640_/A _07640_/B _07640_/C vssd1 vssd1 vccd1 vccd1 _07647_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09998__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ _07571_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07572_/A sky130_fd_sc_hd__nand2_1
X_09310_ _08973_/A _08973_/B _08979_/C vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__o21a_1
X_06522_ _09528_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _06524_/B sky130_fd_sc_hd__nand2_1
X_09241_ _09242_/B _09242_/A vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__or2_1
XFILLER_0_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06453_ _08300_/A vssd1 vssd1 vccd1 vccd1 _06454_/B sky130_fd_sc_hd__inv_2
X_09172_ _09172_/A _09172_/B _09172_/C vssd1 vssd1 vccd1 vccd1 _09173_/B sky130_fd_sc_hd__nand3_1
X_06384_ _06649_/C _06649_/B _06383_/Y vssd1 vssd1 vccd1 vccd1 _06646_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05404_ _05902_/A _05903_/A vssd1 vssd1 vccd1 vccd1 _05404_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _08123_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _08128_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05335_ _05335_/A _05335_/B _05335_/C vssd1 vssd1 vccd1 vccd1 _05903_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08054_ _08054_/A _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08176_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07005_ _07659_/B _07659_/C vssd1 vssd1 vccd1 vccd1 _07658_/A sky130_fd_sc_hd__nand2_1
X_05266_ _05285_/B _05286_/C _05286_/B vssd1 vssd1 vccd1 vccd1 _05502_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08142__B _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _08956_/A _08956_/B vssd1 vssd1 vccd1 vccd1 _08993_/C sky130_fd_sc_hd__nand2_1
X_08887_ _08887_/A _09118_/A _08888_/A vssd1 vssd1 vccd1 vccd1 _09132_/B sky130_fd_sc_hd__nand3_1
X_07907_ _07907_/A _07907_/B vssd1 vssd1 vccd1 vccd1 _07911_/B sky130_fd_sc_hd__nand2_1
X_07838_ _09361_/D _08688_/A vssd1 vssd1 vccd1 vccd1 _07841_/A sky130_fd_sc_hd__nand2_1
X_09508_ _09505_/Y _09506_/Y _09507_/Y vssd1 vssd1 vccd1 vccd1 _09511_/C sky130_fd_sc_hd__a21oi_2
X_07769_ _07769_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09439_/A vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__inv_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10214_ _10215_/B hold77/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__or2_1
X_10145_ _10145_/A _10145_/B _10145_/C vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__nand3_1
X_10076_ _10076_/A _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06970__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _09548_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _08811_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09790_/A vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__inv_2
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08741_ _08754_/A _08754_/B vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__nand2_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05953_ _06325_/B _06325_/C _05952_/Y vssd1 vssd1 vccd1 vccd1 _06328_/A sky130_fd_sc_hd__a21oi_1
X_08672_ _08672_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _08774_/A sky130_fd_sc_hd__nand2_1
X_05884_ _05960_/A _05959_/A vssd1 vssd1 vccd1 vccd1 _05884_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07306__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ _07623_/A _07623_/B _07623_/C vssd1 vssd1 vccd1 vccd1 _07628_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07554_ _07554_/A _10050_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07485_ _07572_/B vssd1 vssd1 vccd1 vccd1 _07540_/C sky130_fd_sc_hd__inv_2
X_06505_ _06505_/A _06505_/B vssd1 vssd1 vccd1 vccd1 _06505_/Y sky130_fd_sc_hd__nor2_1
X_09224_ _09224_/A _09224_/B vssd1 vssd1 vccd1 vccd1 _09231_/B sky130_fd_sc_hd__nand2_1
X_06436_ _06436_/A _08225_/A _06436_/C vssd1 vssd1 vccd1 vccd1 _06438_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_29_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09155_ _09155_/A _09155_/B _09155_/C vssd1 vssd1 vccd1 vccd1 _09175_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06367_ _06369_/B _06369_/C vssd1 vssd1 vccd1 vccd1 _06368_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _09086_/A vssd1 vssd1 vccd1 vccd1 _09087_/C sky130_fd_sc_hd__inv_2
X_08106_ _08158_/B vssd1 vssd1 vccd1 vccd1 _08157_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05318_ input4/X _08247_/B vssd1 vssd1 vccd1 vccd1 _05324_/B sky130_fd_sc_hd__nand2_1
X_06298_ _06298_/A _06298_/B vssd1 vssd1 vccd1 vccd1 _06300_/A sky130_fd_sc_hd__nand2_1
X_08037_ _08037_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05249_ _05338_/A _05337_/A vssd1 vssd1 vccd1 vccd1 _05249_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07992__A _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _09988_/A input25/X vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__nand2_1
X_08939_ _09296_/C _08939_/B vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07216__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08998__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A1 _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__B1 _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__B2 _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A1 _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ _10127_/B _10128_/B _10128_/C vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__nand3b_1
X_10059_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10067_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10114__A2 _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07270_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07270_/Y sky130_fd_sc_hd__nor2_1
X_06221_ _06221_/A _06221_/B vssd1 vssd1 vccd1 vccd1 _06223_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09440__B1 _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06152_ _06162_/A _06162_/B vssd1 vssd1 vccd1 vccd1 _06161_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05597__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06083_ _06083_/A _06083_/B vssd1 vssd1 vccd1 vccd1 _06085_/A sky130_fd_sc_hd__nand2_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _09911_/A _09911_/B vssd1 vssd1 vccd1 vccd1 _09913_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ _09842_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__nand2_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09796_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08420__B input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _08724_/A vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__inv_2
X_06985_ _06985_/A _07127_/A vssd1 vssd1 vccd1 vccd1 _06987_/A sky130_fd_sc_hd__nand2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07036__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05936_ _05936_/A _05936_/B vssd1 vssd1 vccd1 vccd1 _05937_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06875__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05867_ _05867_/A vssd1 vssd1 vccd1 vccd1 _05868_/B sky130_fd_sc_hd__inv_2
X_08655_ _08655_/A _08655_/B vssd1 vssd1 vccd1 vccd1 _08656_/B sky130_fd_sc_hd__or2_1
X_08586_ _08858_/A _08586_/B _08586_/C vssd1 vssd1 vccd1 vccd1 _08590_/C sky130_fd_sc_hd__nand3_1
X_07606_ _07801_/A _07799_/A vssd1 vssd1 vccd1 vccd1 _07606_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07537_ _07537_/A _07537_/B _07537_/C vssd1 vssd1 vccd1 vccd1 _07799_/C sky130_fd_sc_hd__nand3_1
X_05798_ _05798_/A _05808_/A vssd1 vssd1 vccd1 vccd1 _06298_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07468_ _07468_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__nand2_1
X_09207_ _09594_/A _09208_/A vssd1 vssd1 vccd1 vccd1 _09215_/A sky130_fd_sc_hd__or2_1
X_06419_ _06419_/A _08255_/A vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__nand2_1
X_07399_ _07399_/A _07399_/B vssd1 vssd1 vccd1 vccd1 _07400_/B sky130_fd_sc_hd__nand2_1
X_09138_ _09155_/B _09155_/C vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09982__A1 _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05300__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09069_ _09069_/A _09352_/A _09122_/A vssd1 vssd1 vccd1 vccd1 _09414_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_99_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06025__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _06770_/A vssd1 vssd1 vccd1 vccd1 _06771_/B sky130_fd_sc_hd__inv_2
X_05721_ _06185_/B _05725_/C vssd1 vssd1 vccd1 vccd1 _05724_/A sky130_fd_sc_hd__nand2_1
X_08440_ _08714_/B _08441_/C _08441_/B vssd1 vssd1 vccd1 vccd1 _08442_/A sky130_fd_sc_hd__a21o_1
X_05652_ _05486_/C _05486_/B _05478_/Y vssd1 vssd1 vccd1 vccd1 _05665_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _08371_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08372_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05583_ _06065_/A _06065_/B vssd1 vssd1 vccd1 vccd1 _05588_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07322_ _07323_/A _07323_/C _07323_/B vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07253_ _07254_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07253_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07184_ _10043_/B _09988_/A vssd1 vssd1 vccd1 vccd1 _07188_/B sky130_fd_sc_hd__nand2_1
X_06204_ _06208_/A _06208_/B vssd1 vssd1 vccd1 vccd1 _06206_/A sky130_fd_sc_hd__nand2_1
X_06135_ _06135_/A _06585_/B vssd1 vssd1 vccd1 vccd1 _06166_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06066_ _05588_/C _05588_/B _06065_/Y vssd1 vssd1 vccd1 vccd1 _06084_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09825_ _09825_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _10063_/A sky130_fd_sc_hd__nor2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _09756_/A vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__inv_2
X_06968_ _06968_/A _06968_/B vssd1 vssd1 vccd1 vccd1 _06986_/C sky130_fd_sc_hd__nand2_1
X_09687_ _09528_/A _09496_/B _09685_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _09688_/B
+ sky130_fd_sc_hd__a22o_1
X_08707_ _09805_/A _09777_/A _08707_/C vssd1 vssd1 vccd1 vccd1 _08932_/B sky130_fd_sc_hd__or3_1
X_05919_ _05950_/B _05919_/B vssd1 vssd1 vccd1 vccd1 _05920_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05790__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08638_ _08638_/A _08638_/B vssd1 vssd1 vccd1 vccd1 _08638_/Y sky130_fd_sc_hd__nor2_1
X_06899_ _06943_/A _06899_/B _06899_/C vssd1 vssd1 vccd1 vccd1 _06911_/C sky130_fd_sc_hd__nand3_1
X_08569_ _08567_/Y _08569_/B vssd1 vssd1 vccd1 vccd1 _08571_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08325__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10462_ _10494_/CLK _10462_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10393_ _10394_/B _10394_/A vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__or2_1
XANTENNA__09437__A _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10111__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__B1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07940_ _07940_/A _07940_/B vssd1 vssd1 vccd1 vccd1 _07941_/A sky130_fd_sc_hd__nand2_1
X_07871_ _07925_/A _07925_/B _07924_/B vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__nand3_1
X_09610_ _09611_/A _09611_/C _09611_/B vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__a21o_1
X_06822_ _10435_/A _10426_/A vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__nor2_1
X_09541_ _09541_/A _09541_/B vssd1 vssd1 vccd1 vccd1 _09740_/B sky130_fd_sc_hd__xor2_1
X_06753_ _06756_/B vssd1 vssd1 vccd1 vccd1 _06758_/A sky130_fd_sc_hd__inv_4
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05704_ _10043_/A input1/X vssd1 vssd1 vccd1 vccd1 _05742_/A sky130_fd_sc_hd__nand2_1
X_09472_ _09472_/A _09473_/B _09473_/A vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__nand3_1
X_06684_ _06793_/B _06792_/A vssd1 vssd1 vccd1 vccd1 _06684_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08423_ _08425_/B vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__inv_2
X_05635_ input40/X vssd1 vssd1 vccd1 vccd1 _09685_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08354_ _08354_/A _08354_/B vssd1 vssd1 vccd1 vccd1 _08359_/C sky130_fd_sc_hd__nand2_1
X_05566_ _05574_/C vssd1 vssd1 vccd1 vccd1 _05571_/B sky130_fd_sc_hd__inv_2
X_07305_ input36/X vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_73_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08285_ _08297_/B _08297_/C vssd1 vssd1 vccd1 vccd1 _08295_/A sky130_fd_sc_hd__nand2_1
X_05497_ _05404_/Y _05905_/B _05496_/Y vssd1 vssd1 vccd1 vccd1 _05977_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07236_ _07236_/A _07236_/B vssd1 vssd1 vccd1 vccd1 _07237_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ _07172_/C vssd1 vssd1 vccd1 vccd1 _07169_/B sky130_fd_sc_hd__inv_2
X_06118_ _06118_/A vssd1 vssd1 vccd1 vccd1 _06119_/B sky130_fd_sc_hd__inv_2
X_07098_ _07098_/A _07098_/B vssd1 vssd1 vccd1 vccd1 _07357_/B sky130_fd_sc_hd__nand2_1
X_06049_ _06049_/A _06049_/B _06049_/C vssd1 vssd1 vccd1 vccd1 _06100_/C sky130_fd_sc_hd__nand3_1
X_09808_ _09809_/B _09809_/A vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__or2_1
XANTENNA__10482__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _09745_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08336__A _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10448_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10376_ _10375_/Y _10376_/B _10376_/C vssd1 vssd1 vccd1 vccd1 _10378_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05420_ _05420_/A _05420_/B _05420_/C vssd1 vssd1 vccd1 vccd1 _05453_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08246__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05351_ _08422_/A vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__buf_12
XANTENNA__07150__A _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05282_ _05282_/A _05282_/B vssd1 vssd1 vccd1 vccd1 _05287_/C sky130_fd_sc_hd__nand2_1
X_08070_ _08062_/Y _08083_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _10400_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_3_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07021_ _07021_/A _07021_/B _07021_/C vssd1 vssd1 vccd1 vccd1 _07392_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ _09962_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _08973_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07923_ _08035_/B _07935_/A vssd1 vssd1 vccd1 vccd1 _07927_/A sky130_fd_sc_hd__nand2_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_07854_ _07854_/A vssd1 vssd1 vccd1 vccd1 _07855_/C sky130_fd_sc_hd__inv_2
X_06805_ _06805_/A _06805_/B vssd1 vssd1 vccd1 vccd1 _06828_/A sky130_fd_sc_hd__nand2_2
XANTENNA__07325__A _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__B1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ _07925_/A _07924_/B _07784_/Y vssd1 vssd1 vccd1 vccd1 _07816_/A sky130_fd_sc_hd__a21oi_1
X_09524_ _09587_/B _09845_/B vssd1 vssd1 vccd1 vccd1 _09585_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06736_ _06736_/A _06736_/B _06736_/C vssd1 vssd1 vccd1 vccd1 _06737_/B sky130_fd_sc_hd__nand3_1
X_09455_ _09988_/A input22/X _09987_/A input21/X vssd1 vssd1 vccd1 vccd1 _09456_/B
+ sky130_fd_sc_hd__a22o_1
X_06667_ _10052_/A _09980_/A vssd1 vssd1 vccd1 vccd1 _06773_/B sky130_fd_sc_hd__nand2_1
X_08406_ _06582_/A _06583_/B _06591_/A vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__o21a_1
X_05618_ _05618_/A _05619_/A vssd1 vssd1 vccd1 vccd1 _05621_/A sky130_fd_sc_hd__nand2_1
X_09386_ _09647_/B _09387_/A vssd1 vssd1 vccd1 vccd1 _09397_/A sky130_fd_sc_hd__nand2_1
X_06598_ _06598_/A _08317_/A _06598_/C vssd1 vssd1 vccd1 vccd1 _06600_/A sky130_fd_sc_hd__nand3_1
X_08337_ _10051_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _08338_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05549_ _09684_/B _07216_/B vssd1 vssd1 vccd1 vccd1 _05551_/A sky130_fd_sc_hd__nand2_1
X_08268_ _08268_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08313_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07219_ _07272_/A _07275_/B _07274_/A vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__a21oi_1
X_08199_ _08198_/Y _08177_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _08200_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_42_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10230_ _10230_/A hold37/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__xor2_1
X_10161_ _10161_/A _10161_/B _10161_/C vssd1 vssd1 vccd1 vccd1 _10166_/C sky130_fd_sc_hd__nand3_1
X_10092_ _10092_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ _10428_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10429_/C sky130_fd_sc_hd__or2_1
X_10359_ hold60/X _10360_/A vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__or2_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06033__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07570_ _07809_/A _07808_/B _07809_/B vssd1 vssd1 vccd1 vccd1 _07725_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_87_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06521_ _09685_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _06524_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09240_ _09243_/C _09581_/B _09240_/C vssd1 vssd1 vccd1 vccd1 _09581_/A sky130_fd_sc_hd__nand3b_1
X_06452_ _06013_/C _06013_/B _06451_/Y vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ _09171_/A _09171_/B _09171_/C vssd1 vssd1 vccd1 vccd1 _09173_/A sky130_fd_sc_hd__nand3_1
X_06383_ _06736_/A _06735_/A vssd1 vssd1 vccd1 vccd1 _06383_/Y sky130_fd_sc_hd__nor2_1
X_05403_ _05375_/Y _05915_/B _05402_/Y vssd1 vssd1 vccd1 vccd1 _05903_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ _08164_/B _08164_/A vssd1 vssd1 vccd1 vccd1 _08124_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05334_ _05334_/A _05334_/B vssd1 vssd1 vccd1 vccd1 _05903_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ _08053_/A _08056_/B _08053_/C vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07004_ _07004_/A _07004_/B _07004_/C vssd1 vssd1 vccd1 vccd1 _07659_/C sky130_fd_sc_hd__nand3_1
X_05265_ _05265_/A _05265_/B _05265_/C vssd1 vssd1 vccd1 vccd1 _05286_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08955_ _08955_/A _09306_/A vssd1 vssd1 vccd1 vccd1 _08956_/B sky130_fd_sc_hd__nand2_1
X_07906_ _07906_/A _07906_/B vssd1 vssd1 vccd1 vccd1 _07907_/A sky130_fd_sc_hd__nand2_1
X_08886_ _08886_/A _08886_/B _08886_/C vssd1 vssd1 vccd1 vccd1 _08888_/A sky130_fd_sc_hd__nand3_1
X_07837_ _08337_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _07851_/A sky130_fd_sc_hd__nand2_1
X_07768_ _07770_/B vssd1 vssd1 vccd1 vccd1 _07769_/B sky130_fd_sc_hd__inv_2
X_09507_ _09507_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09507_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09270__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06719_ _10027_/A _09392_/C _06295_/C vssd1 vssd1 vccd1 vccd1 _06719_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _07699_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07701_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09438_ _10000_/A _09999_/A _09775_/B _09998_/B vssd1 vssd1 vccd1 vccd1 _09439_/A
+ sky130_fd_sc_hd__and4_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ _09369_/A _09369_/B vssd1 vssd1 vccd1 vccd1 _09370_/B sky130_fd_sc_hd__nand2_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10213_ _10213_/A hold76/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__nand2_1
X_10144_ _10144_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__nand2_1
X_10075_ _10075_/A _10075_/B _10075_/C vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05213__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08524__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ _08740_/A _08740_/B _08740_/C vssd1 vssd1 vccd1 vccd1 _08754_/B sky130_fd_sc_hd__nand3_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05952_ _06334_/A _06333_/A vssd1 vssd1 vccd1 vccd1 _05952_/Y sky130_fd_sc_hd__nor2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08671_ _10441_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _10442_/A sky130_fd_sc_hd__nand2_1
X_05883_ _05875_/B _05874_/A _06377_/B vssd1 vssd1 vccd1 vccd1 _05962_/B sky130_fd_sc_hd__o21ai_2
X_07622_ _08206_/B vssd1 vssd1 vccd1 vccd1 _07652_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07553_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07554_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07484_ _07484_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07572_/B sky130_fd_sc_hd__nand2_1
X_06504_ _06505_/B _06505_/A vssd1 vssd1 vccd1 vccd1 _06504_/Y sky130_fd_sc_hd__nand2_1
X_09223_ _09224_/B _09224_/A vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__or2_1
X_06435_ _06435_/A _06435_/B vssd1 vssd1 vccd1 vccd1 _06438_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09154_ _09154_/A _09154_/B vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08434__A _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ _10111_/B _10126_/B _09981_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _08158_/B
+ sky130_fd_sc_hd__and4_1
X_06366_ _06366_/A _06366_/B _06366_/C vssd1 vssd1 vccd1 vccd1 _06369_/C sky130_fd_sc_hd__nand3_1
X_09085_ _09085_/A _09086_/A vssd1 vssd1 vccd1 vccd1 _09089_/A sky130_fd_sc_hd__nand2_1
X_05317_ _05324_/A vssd1 vssd1 vccd1 vccd1 _05320_/A sky130_fd_sc_hd__inv_2
X_06297_ _06303_/A _06720_/A _06304_/B vssd1 vssd1 vccd1 vccd1 _06302_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08036_ _08037_/A _08036_/B _08037_/B vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__nand3_1
X_05248_ _05339_/C vssd1 vssd1 vccd1 vccd1 _05291_/C sky130_fd_sc_hd__inv_2
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09987_ _09987_/A input24/X vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__nand2_1
X_08938_ _10000_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _08939_/B sky130_fd_sc_hd__nand2_1
X_08869_ _08873_/B _09071_/A vssd1 vssd1 vccd1 vccd1 _08872_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08998__B _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09201__B2 _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A1 _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A2 _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__nand2_1
X_10058_ _10060_/B vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__inv_2
XANTENNA__05208__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06220_ _06377_/B _06377_/C vssd1 vssd1 vccd1 vccd1 _06376_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09440__A1 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06151_ _06151_/A _06151_/B _06151_/C vssd1 vssd1 vccd1 vccd1 _06162_/B sky130_fd_sc_hd__nand3_1
XANTENNA__05597__B _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09440__B2 _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06082_ _06085_/C _06511_/B _06082_/C vssd1 vssd1 vccd1 vccd1 _06511_/A sky130_fd_sc_hd__nand3b_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _09910_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09911_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09841_ _09841_/A _09842_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_95_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09772_/A vssd1 vssd1 vccd1 vccd1 _09796_/A sky130_fd_sc_hd__inv_2
X_06984_ _07400_/A _07126_/A vssd1 vssd1 vccd1 vccd1 _07127_/A sky130_fd_sc_hd__or2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08723_/A _08724_/A vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__nand2_1
X_05935_ _05935_/A _05935_/B _05935_/C vssd1 vssd1 vccd1 vccd1 _06334_/B sky130_fd_sc_hd__nand3_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08654_ _08654_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _08663_/A sky130_fd_sc_hd__nand2_1
X_05866_ _05866_/A vssd1 vssd1 vccd1 vccd1 _05868_/A sky130_fd_sc_hd__inv_2
XFILLER_0_95_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08585_ _08858_/B _08585_/B vssd1 vssd1 vccd1 vccd1 _08590_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07333__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05797_ _06268_/C _06268_/B _05796_/Y vssd1 vssd1 vccd1 vccd1 _05808_/A sky130_fd_sc_hd__a21oi_1
X_07605_ _07597_/Y _07721_/B _07604_/Y vssd1 vssd1 vccd1 vccd1 _07799_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07536_ _07536_/A _07536_/B vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09206_ _09594_/B vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__inv_2
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07467_ _07467_/A vssd1 vssd1 vccd1 vccd1 _07468_/A sky130_fd_sc_hd__inv_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06418_ _08255_/B _06418_/B _06418_/C vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__nand3_1
X_07398_ _07404_/B _07404_/C vssd1 vssd1 vccd1 vccd1 _07403_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09137_ _09137_/A _09137_/B _09137_/C vssd1 vssd1 vccd1 vccd1 _09155_/C sky130_fd_sc_hd__nand3_1
X_06349_ _06757_/C vssd1 vssd1 vccd1 vccd1 _06759_/B sky130_fd_sc_hd__inv_2
X_09068_ _09068_/A _09068_/B vssd1 vssd1 vccd1 vccd1 _09122_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05300__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08019_ _08116_/B vssd1 vssd1 vccd1 vccd1 _08019_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06412__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07243__A _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05698__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05720_ _05720_/A _05720_/B vssd1 vssd1 vccd1 vccd1 _05725_/C sky130_fd_sc_hd__nand2_1
X_05651_ _05694_/C _05694_/B vssd1 vssd1 vccd1 vccd1 _05665_/B sky130_fd_sc_hd__nand2_1
X_08370_ _08370_/A vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__inv_2
XFILLER_0_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07321_ _07321_/A vssd1 vssd1 vccd1 vccd1 _07323_/A sky130_fd_sc_hd__inv_2
X_05582_ _05582_/A _05582_/B vssd1 vssd1 vccd1 vccd1 _05588_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ _10050_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _07254_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06203_ _06628_/B _06203_/B vssd1 vssd1 vccd1 vccd1 _06208_/B sky130_fd_sc_hd__nand2_1
X_07183_ _10052_/A _08420_/A vssd1 vssd1 vccd1 vccd1 _07188_/A sky130_fd_sc_hd__nand2_1
X_06134_ _06134_/A _06134_/B vssd1 vssd1 vccd1 vccd1 _06585_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06065_ _06065_/A _06065_/B vssd1 vssd1 vccd1 vccd1 _06065_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07328__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _09825_/A _09825_/B _10063_/B vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__o21ai_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09456_/B _09986_/A input20/X _09454_/X vssd1 vssd1 vccd1 vccd1 _09756_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06967_ _06967_/A _06967_/B vssd1 vssd1 vccd1 vccd1 _06992_/B sky130_fd_sc_hd__nand2_1
X_09686_ _10027_/A _10027_/C _10027_/D _09686_/D vssd1 vssd1 vccd1 vccd1 _10034_/B
+ sky130_fd_sc_hd__or4_1
X_08706_ _09963_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _08707_/C sky130_fd_sc_hd__nand2_1
X_05918_ _05919_/B _05918_/B _05918_/C vssd1 vssd1 vccd1 vccd1 _05950_/B sky130_fd_sc_hd__nand3_1
X_06898_ _06943_/B _06898_/B vssd1 vssd1 vccd1 vccd1 _06911_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05790__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08637_ _08638_/B _08638_/A vssd1 vssd1 vccd1 vccd1 _08637_/Y sky130_fd_sc_hd__nand2_1
X_05849_ _06222_/B _06221_/B vssd1 vssd1 vccd1 vccd1 _05850_/C sky130_fd_sc_hd__nand2_1
X_08568_ _09083_/A _10113_/B _08567_/C vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08499_ _08499_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08500_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07519_ _07609_/A _07610_/A vssd1 vssd1 vccd1 vccd1 _07524_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout98 fanout99/X vssd1 vssd1 vccd1 vccd1 fanout98/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10461_ _10495_/CLK _10461_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfrtp_1
X_10392_ _10391_/A _10390_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _10394_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09437__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__A _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10111__B _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__B2 _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05221__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07870_ _07924_/A _07925_/C vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06821_ _06821_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10426_/A sky130_fd_sc_hd__nand2_1
X_09540_ _09540_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09541_/B sky130_fd_sc_hd__nand2_1
X_06752_ _06845_/B _06845_/C vssd1 vssd1 vccd1 vccd1 _06847_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09471_ _09474_/A _09770_/A vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__nand2_1
X_05703_ input45/X vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__buf_4
X_08422_ _08422_/A input18/X vssd1 vssd1 vccd1 vccd1 _08425_/B sky130_fd_sc_hd__nand2_1
X_06683_ _06671_/Y _06784_/B _06682_/Y vssd1 vssd1 vccd1 vccd1 _06792_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05634_ _05785_/A _05785_/B vssd1 vssd1 vccd1 vccd1 _05784_/A sky130_fd_sc_hd__nand2_1
X_08353_ _08354_/B _08354_/A vssd1 vssd1 vccd1 vccd1 _08537_/A sky130_fd_sc_hd__or2_1
X_05565_ _05565_/A _05565_/B vssd1 vssd1 vccd1 vccd1 _05574_/C sky130_fd_sc_hd__nand2_1
X_08284_ _08510_/A _08489_/A _08284_/C vssd1 vssd1 vccd1 vccd1 _08297_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07304_ _07313_/A _07313_/B vssd1 vssd1 vccd1 vccd1 _07312_/A sky130_fd_sc_hd__nand2_1
X_07235_ _07235_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05496_ _05903_/A _05902_/A vssd1 vssd1 vccd1 vccd1 _05496_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07166_ _09720_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _07172_/C sky130_fd_sc_hd__nand2_1
X_06117_ _06117_/A _06118_/A vssd1 vssd1 vccd1 vccd1 _06129_/A sky130_fd_sc_hd__nand2_1
X_07097_ _07097_/A _07097_/B vssd1 vssd1 vccd1 vccd1 _07098_/A sky130_fd_sc_hd__nand2_1
X_06048_ _06048_/A _06048_/B vssd1 vssd1 vccd1 vccd1 _06100_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09807_ _09957_/B _09807_/B vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__nand2_1
X_07999_ _08014_/B _08000_/C _08000_/B vssd1 vssd1 vccd1 vccd1 _08001_/A sky130_fd_sc_hd__a21o_1
X_09738_ _09738_/A _09738_/B _10134_/A vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09669_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09672_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09720__B _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06137__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10444_ _10445_/B _10445_/A vssd1 vssd1 vccd1 vccd1 _10446_/A sky130_fd_sc_hd__or2_1
X_10375_ hold69/A hold1/X vssd1 vssd1 vccd1 vccd1 _10375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08246__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05350_ _09816_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _05934_/B sky130_fd_sc_hd__nand2_2
XANTENNA__07150__B _07150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05281_ _05281_/A _05281_/B _05281_/C vssd1 vssd1 vccd1 vccd1 _05282_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07020_ _07020_/A _07020_/B vssd1 vssd1 vccd1 vccd1 _07392_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _09960_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _08973_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09805__B _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ _07935_/A _07935_/B _07922_/C vssd1 vssd1 vccd1 vccd1 _08035_/B sky130_fd_sc_hd__nand3_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _07853_/A _07854_/A vssd1 vssd1 vccd1 vccd1 _07862_/A sky130_fd_sc_hd__nand2_1
X_06804_ _06825_/A _06823_/A vssd1 vssd1 vccd1 vccd1 _06804_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07325__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__A1 _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__B2 _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _07784_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07784_/Y sky130_fd_sc_hd__nor2_1
X_09523_ _09523_/A _09523_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _09845_/B sky130_fd_sc_hd__nand3_2
X_06735_ _06735_/A _06735_/B vssd1 vssd1 vccd1 vccd1 _06737_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _09988_/A _09987_/A input21/X input22/X vssd1 vssd1 vccd1 vccd1 _09454_/X
+ sky130_fd_sc_hd__and4_1
X_06666_ _06769_/A _06770_/A vssd1 vssd1 vccd1 vccd1 _06774_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09385_ _09385_/A _09385_/B vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__nand2_1
X_08405_ _08630_/B _08405_/B vssd1 vssd1 vccd1 vccd1 _08408_/B sky130_fd_sc_hd__nand2_1
X_05617_ _05617_/A _05617_/B vssd1 vssd1 vccd1 vccd1 _05619_/A sky130_fd_sc_hd__nand2_2
X_08336_ _09361_/D vssd1 vssd1 vccd1 vccd1 _10113_/D sky130_fd_sc_hd__inv_2
XFILLER_0_74_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06597_ _08388_/B _06597_/B _06597_/C vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05548_ _06043_/B _05552_/C vssd1 vssd1 vccd1 vccd1 _05550_/A sky130_fd_sc_hd__nand2_1
X_08267_ _08314_/A _08314_/C vssd1 vssd1 vccd1 vccd1 _08313_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05479_ _05479_/A _05479_/B vssd1 vssd1 vccd1 vccd1 _05486_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08198_ _10390_/B vssd1 vssd1 vccd1 vccd1 _08198_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07218_ _07218_/A _07218_/B vssd1 vssd1 vccd1 vccd1 _07274_/A sky130_fd_sc_hd__nor2_1
X_07149_ _07151_/B _07154_/B _07150_/B vssd1 vssd1 vccd1 vccd1 _07710_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10160_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10091_ _10091_/A _10091_/B vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06420__A _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08347__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__A _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10427_ _10427_/A _10427_/B vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10358_ _10360_/A hold50/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__nor2_1
XANTENNA__08810__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ hold84/X vssd1 vssd1 vccd1 vccd1 _10494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07426__A _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06520_ _06599_/B _08317_/A _06598_/C vssd1 vssd1 vccd1 vccd1 _08388_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_87_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06451_ _06451_/A vssd1 vssd1 vccd1 vccd1 _06451_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05402_ _05908_/A _05913_/A vssd1 vssd1 vccd1 vccd1 _05402_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09170_ _09170_/A _09182_/B vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__nand2_1
X_06382_ _06737_/C vssd1 vssd1 vccd1 vccd1 _06649_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08121_ _08127_/B _08127_/C vssd1 vssd1 vccd1 vccd1 _08164_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05333_ _05335_/C vssd1 vssd1 vccd1 vccd1 _05334_/B sky130_fd_sc_hd__inv_2
XANTENNA__10472__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ _08087_/B vssd1 vssd1 vccd1 vccd1 _08053_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05264_ _05264_/A _05503_/A vssd1 vssd1 vccd1 vccd1 _05265_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07003_ _07003_/A _07003_/B vssd1 vssd1 vccd1 vccd1 _07659_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10027__A _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08954_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08956_/A sky130_fd_sc_hd__inv_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07905_ _08065_/B _08065_/A vssd1 vssd1 vccd1 vccd1 _07912_/A sky130_fd_sc_hd__nor2_1
X_08885_ _08885_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _08886_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07836_ _07836_/A _07836_/B vssd1 vssd1 vccd1 vccd1 _07938_/A sky130_fd_sc_hd__nand2_1
X_07767_ _07767_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _07770_/B sky130_fd_sc_hd__nand2_1
X_09506_ _09506_/A vssd1 vssd1 vccd1 vccd1 _09506_/Y sky130_fd_sc_hd__inv_2
X_06718_ _06303_/A _06304_/B _06720_/A vssd1 vssd1 vccd1 vccd1 _06962_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07698_ _07700_/A vssd1 vssd1 vccd1 vccd1 _07699_/B sky130_fd_sc_hd__inv_2
X_09437_ _09998_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09443_/B sky130_fd_sc_hd__nand2_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06649_ _06650_/B _06649_/B _06649_/C vssd1 vssd1 vccd1 vccd1 _06831_/B sky130_fd_sc_hd__nand3_1
X_09368_ _09368_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _09608_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09299_ _09300_/A _09300_/C _09506_/A vssd1 vssd1 vccd1 vccd1 _09301_/A sky130_fd_sc_hd__a21o_1
X_08319_ _08319_/A vssd1 vssd1 vccd1 vccd1 _08597_/A sky130_fd_sc_hd__inv_2
XFILLER_0_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06415__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ _10212_/A hold71/X vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__and2_1
X_10143_ _10145_/C vssd1 vssd1 vccd1 vccd1 _10144_/B sky130_fd_sc_hd__inv_2
XANTENNA__07246__A _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10495__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08524__B _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06060__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05951_ _06335_/C vssd1 vssd1 vccd1 vccd1 _06325_/C sky130_fd_sc_hd__inv_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08670_ _08670_/A vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__inv_2
X_05882_ _05882_/A _05882_/B vssd1 vssd1 vccd1 vccd1 _06377_/B sky130_fd_sc_hd__nand2_1
X_07621_ _07913_/A _07621_/B _07913_/B vssd1 vssd1 vccd1 vccd1 _08206_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07552_ _07734_/B vssd1 vssd1 vccd1 vccd1 _07567_/C sky130_fd_sc_hd__inv_2
XFILLER_0_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06503_ _08306_/A _06509_/C vssd1 vssd1 vccd1 vccd1 _08374_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07483_ _07483_/A _07483_/B _07483_/C vssd1 vssd1 vccd1 vccd1 _07484_/B sky130_fd_sc_hd__nand3_1
X_09222_ _09526_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__nand2b_1
X_06434_ _06436_/A vssd1 vssd1 vccd1 vccd1 _06435_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _09155_/A vssd1 vssd1 vccd1 vccd1 _09154_/B sky130_fd_sc_hd__inv_2
X_06365_ _06365_/A _06365_/B vssd1 vssd1 vccd1 vccd1 _06369_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08434__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ _08109_/B _08109_/A vssd1 vssd1 vccd1 vccd1 _08137_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05316_ input5/X _08248_/B vssd1 vssd1 vccd1 vccd1 _05324_/A sky130_fd_sc_hd__nand2_1
X_09084_ _09082_/Y _08828_/B _09083_/Y vssd1 vssd1 vccd1 vccd1 _09086_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06296_ _06296_/A _06299_/A _06296_/C vssd1 vssd1 vccd1 vccd1 _06304_/B sky130_fd_sc_hd__nand3_2
X_08035_ _08035_/A _08035_/B _08035_/C vssd1 vssd1 vccd1 vccd1 _08037_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05247_ _05247_/A _05247_/B vssd1 vssd1 vccd1 vccd1 _05339_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09986_ _09986_/A input22/X vssd1 vssd1 vccd1 vccd1 _09990_/A sky130_fd_sc_hd__nand2_1
X_08937_ _09951_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _09296_/C sky130_fd_sc_hd__nand2_1
X_08868_ _08867_/B _09071_/B _08868_/C vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__09281__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__C1 _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07819_ _07819_/A _07819_/B _07819_/C vssd1 vssd1 vccd1 vccd1 _07921_/C sky130_fd_sc_hd__nand3_1
X_08799_ _08806_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09201__A2 _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ input57/X _10126_/B vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__nand2_1
X_10057_ _10057_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _10060_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05208__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05224__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09440__A2 _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06150_ _06150_/A _06150_/B vssd1 vssd1 vccd1 vccd1 _06162_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06055__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06081_ _06083_/A _06084_/B vssd1 vssd1 vccd1 vccd1 _06082_/C sky130_fd_sc_hd__nand2_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09366__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09840_ _09840_/A _10019_/A _09840_/C vssd1 vssd1 vccd1 vccd1 _10078_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09773_/B _09773_/A vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__nor2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _06983_/A _06983_/B vssd1 vssd1 vccd1 vccd1 _07126_/A sky130_fd_sc_hd__nand2_1
X_08722_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08724_/A sky130_fd_sc_hd__nand2_1
X_05934_ _05936_/B _05934_/B vssd1 vssd1 vccd1 vccd1 _05935_/B sky130_fd_sc_hd__nand2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08653_ _08657_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _08654_/A sky130_fd_sc_hd__nand2_1
X_05865_ _06260_/C _06260_/B _05864_/Y vssd1 vssd1 vccd1 vccd1 _05875_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_95_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08584_ _08858_/A vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07333__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05796_ _05796_/A _05796_/B vssd1 vssd1 vccd1 vccd1 _05796_/Y sky130_fd_sc_hd__nor2_1
X_07604_ _07717_/A _07719_/B vssd1 vssd1 vccd1 vccd1 _07604_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07535_ _07537_/A _07537_/B vssd1 vssd1 vccd1 vccd1 _07536_/A sky130_fd_sc_hd__nand2_1
X_07466_ _07467_/A _07466_/B _07466_/C vssd1 vssd1 vccd1 vccd1 _07471_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ _09555_/A _09205_/B vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06417_ _06417_/A vssd1 vssd1 vccd1 vccd1 _06418_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07397_ _07631_/B _07397_/B vssd1 vssd1 vccd1 vccd1 _07404_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09136_ _09136_/A _09136_/B _09414_/A vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__nand3_1
X_06348_ _09684_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _06757_/C sky130_fd_sc_hd__nand2_1
X_09067_ _09352_/B _09067_/B vssd1 vssd1 vccd1 vccd1 _09068_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06279_ _06299_/B _06279_/B vssd1 vssd1 vccd1 vccd1 _06280_/A sky130_fd_sc_hd__nand2_1
X_08018_ _08018_/A _08018_/B vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06412__B _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09969_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10492__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07243__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10509__RESET_B fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ _10117_/A _10109_/B _10109_/C vssd1 vssd1 vccd1 vccd1 _10109_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05650_ _05683_/B _05650_/B _05650_/C vssd1 vssd1 vccd1 vccd1 _05694_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05581_ _06065_/B vssd1 vssd1 vccd1 vccd1 _05582_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07320_ _07339_/A _07339_/B vssd1 vssd1 vccd1 vccd1 _07338_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07251_ _09720_/B _09981_/B vssd1 vssd1 vccd1 vccd1 _07254_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07182_ _07182_/A _07182_/B vssd1 vssd1 vccd1 vccd1 _07236_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06202_ _06394_/C _06394_/B _05974_/Y vssd1 vssd1 vccd1 vccd1 _06203_/B sky130_fd_sc_hd__a21o_1
X_06133_ _06133_/A _06133_/B vssd1 vssd1 vccd1 vccd1 _06135_/A sky130_fd_sc_hd__nand2_1
X_06064_ _06064_/A _06064_/B vssd1 vssd1 vccd1 vccd1 _06085_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07328__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _09826_/A _09975_/A vssd1 vssd1 vccd1 vccd1 _10063_/B sky130_fd_sc_hd__nand2_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _09754_/A _09754_/B vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__xor2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06966_ _06968_/B vssd1 vssd1 vccd1 vccd1 _06967_/B sky130_fd_sc_hd__inv_2
X_08705_ _09951_/B vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__inv_2
X_09685_ _09685_/A vssd1 vssd1 vccd1 vccd1 _10027_/C sky130_fd_sc_hd__inv_2
X_05917_ _06316_/B _06316_/C vssd1 vssd1 vccd1 vccd1 _06318_/A sky130_fd_sc_hd__nand2_1
X_06897_ _06943_/A vssd1 vssd1 vccd1 vccd1 _06898_/B sky130_fd_sc_hd__inv_2
X_08636_ _08642_/B _08642_/C vssd1 vssd1 vccd1 vccd1 _09166_/B sky130_fd_sc_hd__nand2_1
X_05848_ _06223_/C vssd1 vssd1 vccd1 vccd1 _05850_/B sky130_fd_sc_hd__inv_2
XFILLER_0_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08567_ _09083_/A _10113_/B _08567_/C vssd1 vssd1 vccd1 vccd1 _08567_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__05799__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05779_ _05781_/C vssd1 vssd1 vccd1 vccd1 _05780_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08498_ _08498_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08499_/B sky130_fd_sc_hd__nand2_1
X_07518_ _07536_/B _07516_/Y _07517_/Y vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout99 fanout99/A vssd1 vssd1 vccd1 vccd1 fanout99/X sky130_fd_sc_hd__clkbuf_8
X_07449_ _07451_/A _07451_/C vssd1 vssd1 vccd1 vccd1 _07450_/A sky130_fd_sc_hd__nand2_1
X_10460_ _10494_/CLK _10460_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfrtp_1
X_09119_ _09119_/A _09418_/B _09119_/C vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08903__A _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10391_ _10391_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10459_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06423__A _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08143__A2 _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__A2 _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05221__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09628__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08906__A1 _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _06820_/A _06820_/B _06820_/C vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06751_ _06751_/A _06751_/B _06751_/C vssd1 vssd1 vccd1 vccd1 _06845_/C sky130_fd_sc_hd__nand3_1
XANTENNA__07164__A _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _09469_/B _09470_/B _09770_/B vssd1 vssd1 vccd1 vccd1 _09770_/A sky130_fd_sc_hd__nand3b_2
X_05702_ _05706_/A _05706_/B vssd1 vssd1 vccd1 vccd1 _05702_/Y sky130_fd_sc_hd__nand2_1
X_06682_ _06782_/A _06781_/A vssd1 vssd1 vccd1 vccd1 _06682_/Y sky130_fd_sc_hd__nor2_1
X_08421_ _08425_/A vssd1 vssd1 vccd1 vccd1 _08424_/A sky130_fd_sc_hd__inv_2
XFILLER_0_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08707__B _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05633_ _05977_/B _05633_/B vssd1 vssd1 vccd1 vccd1 _05785_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08352_ _08537_/B _08352_/B vssd1 vssd1 vccd1 vccd1 _08354_/A sky130_fd_sc_hd__nand2_1
X_05564_ _05564_/A _05564_/B _05564_/C vssd1 vssd1 vccd1 vccd1 _05565_/B sky130_fd_sc_hd__nand3_1
X_08283_ _08283_/A vssd1 vssd1 vccd1 vccd1 _08510_/A sky130_fd_sc_hd__inv_2
X_07303_ _07303_/A _07303_/B _07366_/A vssd1 vssd1 vccd1 vccd1 _07313_/B sky130_fd_sc_hd__nand3_1
X_05495_ _05906_/C vssd1 vssd1 vccd1 vccd1 _05905_/B sky130_fd_sc_hd__inv_2
X_07234_ _07234_/A _07234_/B _07234_/C vssd1 vssd1 vccd1 vccd1 _07466_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07165_ _07170_/A _07171_/A vssd1 vssd1 vccd1 vccd1 _07165_/Y sky130_fd_sc_hd__nor2_1
X_06116_ _10026_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _06118_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07096_ _07096_/A _07096_/B vssd1 vssd1 vccd1 vccd1 _07097_/A sky130_fd_sc_hd__nand2_1
X_06047_ _06049_/C vssd1 vssd1 vccd1 vccd1 _06048_/B sky130_fd_sc_hd__inv_2
XFILLER_0_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09806_ _09951_/B _09804_/A _09485_/C _09437_/B vssd1 vssd1 vccd1 vccd1 _09807_/B
+ sky130_fd_sc_hd__a22o_1
X_07998_ _07998_/A vssd1 vssd1 vccd1 vccd1 _08000_/B sky130_fd_sc_hd__inv_2
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09737_ _10134_/B _09737_/B vssd1 vssd1 vccd1 vccd1 _09745_/A sky130_fd_sc_hd__nand2_1
X_06949_ _06959_/A _06949_/B _06949_/C vssd1 vssd1 vccd1 vccd1 _06951_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09668_ _09672_/B _09682_/A vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__nand2_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ input49/X _10083_/B input50/X _09854_/B vssd1 vssd1 vccd1 vccd1 _09600_/B
+ sky130_fd_sc_hd__a22o_1
X_08619_ _08886_/B _08621_/C vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__nand2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05322__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06137__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10443_ _10437_/A _10442_/Y _09190_/Y vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__a21o_1
X_10374_ hold21/X vssd1 vssd1 vccd1 vccd1 _10378_/A sky130_fd_sc_hd__inv_2
XFILLER_0_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09464__A _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05280_ _05280_/A vssd1 vssd1 vccd1 vccd1 _05281_/B sky130_fd_sc_hd__inv_2
XFILLER_0_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08970_ _08970_/A vssd1 vssd1 vccd1 vccd1 _08975_/B sky130_fd_sc_hd__inv_2
X_07921_ _07921_/A _07921_/B _07921_/C vssd1 vssd1 vccd1 vccd1 _07933_/B sky130_fd_sc_hd__nand3_1
X_07852_ _07841_/Y _07851_/Y _07842_/A vssd1 vssd1 vccd1 vccd1 _07854_/A sky130_fd_sc_hd__a21oi_1
X_06803_ _06838_/B _06801_/Y _06802_/Y vssd1 vssd1 vccd1 vccd1 _06823_/A sky130_fd_sc_hd__a21oi_1
Xinput1 a_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
X_09522_ _09522_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09587_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08107__A2 _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07783_ _07783_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06734_ _06839_/C vssd1 vssd1 vccd1 vccd1 _06838_/B sky130_fd_sc_hd__inv_2
XFILLER_0_78_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09453_ _09986_/A input20/X vssd1 vssd1 vccd1 vccd1 _09458_/B sky130_fd_sc_hd__nand2_1
X_06665_ _09533_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _06770_/A sky130_fd_sc_hd__nand2_1
X_09384_ _09388_/A _09388_/B vssd1 vssd1 vccd1 vccd1 _09647_/B sky130_fd_sc_hd__nand2_1
X_08404_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08405_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05616_ _05620_/A _05620_/B vssd1 vssd1 vccd1 vccd1 _05618_/A sky130_fd_sc_hd__nand2_1
X_08335_ input46/X vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__inv_2
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06596_ _06599_/A _06598_/A vssd1 vssd1 vccd1 vccd1 _06597_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05547_ _05547_/A _05547_/B vssd1 vssd1 vccd1 vccd1 _05552_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08291__A1 _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ _08266_/A _08266_/B _08266_/C vssd1 vssd1 vccd1 vccd1 _08314_/C sky130_fd_sc_hd__nand3_2
X_05478_ _05479_/A _05479_/B vssd1 vssd1 vccd1 vccd1 _05478_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08197_ _08197_/A _08197_/B vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07217_ _07217_/A vssd1 vssd1 vccd1 vccd1 _07275_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07148_ _07148_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07150_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07079_ _07088_/B _07079_/B vssd1 vssd1 vccd1 vccd1 _07082_/A sky130_fd_sc_hd__nand2_1
X_10090_ _10093_/B _10093_/C vssd1 vssd1 vccd1 vccd1 _10092_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06420__B _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__B _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10426_ _10426_/A vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10357_ _10357_/A _10357_/B vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__and2_1
XANTENNA__08810__B _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10293_/A hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__and2_1
XANTENNA__06611__A _06618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06450_ _06455_/B _08260_/A vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__nand2_1
X_05401_ _05916_/C vssd1 vssd1 vccd1 vccd1 _05915_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06381_ _06381_/A _06381_/B vssd1 vssd1 vccd1 vccd1 _06737_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08120_ _08120_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08127_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05332_ _05614_/A _05332_/B vssd1 vssd1 vccd1 vccd1 _05335_/C sky130_fd_sc_hd__nand2_1
X_08051_ _08059_/B _08087_/B vssd1 vssd1 vccd1 vccd1 _08171_/A sky130_fd_sc_hd__nand2_1
X_05263_ _05263_/A _05503_/B vssd1 vssd1 vccd1 vccd1 _05265_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07002_ _07004_/A _07004_/B vssd1 vssd1 vccd1 vccd1 _07003_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09816__B _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _08954_/A _08955_/A _09306_/A vssd1 vssd1 vccd1 vccd1 _09345_/B sky130_fd_sc_hd__nand3_2
XANTENNA__06521__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07904_ _08064_/C _08064_/B vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10043__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ _08885_/A _08885_/B _08884_/C vssd1 vssd1 vccd1 vccd1 _09118_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07835_ _07846_/B vssd1 vssd1 vccd1 vccd1 _07836_/B sky130_fd_sc_hd__inv_2
XFILLER_0_78_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07766_ _07770_/A _07770_/C vssd1 vssd1 vccd1 vccd1 _07769_/A sky130_fd_sc_hd__nand2_1
X_09505_ _09507_/B _09507_/A vssd1 vssd1 vccd1 vccd1 _09505_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ _06732_/A _06805_/B vssd1 vssd1 vccd1 vccd1 _06730_/A sky130_fd_sc_hd__nand2_1
X_09436_ _09802_/A vssd1 vssd1 vccd1 vccd1 _09446_/B sky130_fd_sc_hd__inv_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07697_ _07697_/A _07697_/B vssd1 vssd1 vccd1 vccd1 _07700_/A sky130_fd_sc_hd__nor2_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06648_ _06735_/B _06736_/B _06736_/C vssd1 vssd1 vccd1 vccd1 _06650_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09367_ _09369_/B vssd1 vssd1 vccd1 vccd1 _09368_/B sky130_fd_sc_hd__inv_2
X_06579_ _06579_/A _06579_/B vssd1 vssd1 vccd1 vccd1 _06579_/Y sky130_fd_sc_hd__nor2_1
X_09298_ _09298_/A _09298_/B vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08318_ _08597_/B _08319_/A vssd1 vssd1 vccd1 vccd1 _08386_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08249_ _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08464_/B sky130_fd_sc_hd__or2_1
XFILLER_0_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06415__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ _10485_/Q hold70/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10145_/C sky130_fd_sc_hd__nor2_1
X_10073_ _10075_/A vssd1 vssd1 vccd1 vccd1 _10074_/B sky130_fd_sc_hd__inv_2
XFILLER_0_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07246__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ _10409_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10465_/D sky130_fd_sc_hd__xor2_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06060__B _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05950_ _05950_/A _05950_/B vssd1 vssd1 vccd1 vccd1 _06335_/C sky130_fd_sc_hd__nand2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05881_ _06219_/C vssd1 vssd1 vccd1 vccd1 _05882_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _07620_/A _07620_/B _07620_/C vssd1 vssd1 vccd1 vccd1 _07913_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07551_ _09560_/B input55/X vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06502_ _06502_/A _06502_/B _06502_/C vssd1 vssd1 vccd1 vccd1 _06509_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07482_ _07482_/A _07482_/B vssd1 vssd1 vccd1 vccd1 _07484_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _09528_/A _09684_/B _09685_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _09222_/B
+ sky130_fd_sc_hd__a22o_1
X_06433_ _05996_/C _05996_/B _06432_/Y vssd1 vssd1 vccd1 vccd1 _06436_/A sky130_fd_sc_hd__a21o_1
X_09152_ _09171_/B _09171_/C _09151_/Y vssd1 vssd1 vccd1 vccd1 _09155_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06364_ _06366_/A vssd1 vssd1 vccd1 vccd1 _06365_/B sky130_fd_sc_hd__inv_2
X_08103_ _08103_/A _08103_/B vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__xor2_1
X_05315_ _05328_/B _05559_/A _05329_/A vssd1 vssd1 vccd1 vccd1 _05614_/B sky130_fd_sc_hd__nand3_1
X_09083_ _09083_/A _09856_/D _09083_/C vssd1 vssd1 vccd1 vccd1 _09083_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06295_ _10027_/A _09392_/C _06295_/C vssd1 vssd1 vccd1 vccd1 _06720_/A sky130_fd_sc_hd__nor3_1
X_08034_ _08034_/A vssd1 vssd1 vccd1 vccd1 _08035_/A sky130_fd_sc_hd__inv_2
X_05246_ _05246_/A _05246_/B _05246_/C vssd1 vssd1 vccd1 vccd1 _05247_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09985_ _09753_/B _09986_/A input21/X _09751_/Y vssd1 vssd1 vccd1 vccd1 _09991_/A
+ sky130_fd_sc_hd__a31oi_1
X_08936_ _08936_/A vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__inv_2
XANTENNA__09562__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _08867_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _08873_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09281__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _07889_/B _07818_/B vssd1 vssd1 vccd1 vccd1 _07819_/C sky130_fd_sc_hd__nand2b_1
X_08798_ _08797_/B _08798_/B _08798_/C vssd1 vssd1 vccd1 vccd1 _08806_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_67_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07749_ _07749_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07754_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09419_ _09421_/C vssd1 vssd1 vccd1 vccd1 _09420_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _10128_/B _10128_/C vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__nand2_1
X_10056_ _10056_/A _10055_/A vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__or2b_1
XANTENNA__10462__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05224__B input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06055__B _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
X_06080_ _06084_/A _06084_/C vssd1 vssd1 vccd1 vccd1 _06083_/A sky130_fd_sc_hd__nand2_1
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09366__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09770_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__and2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ _06982_/A _06982_/B vssd1 vssd1 vccd1 vccd1 _06983_/B sky130_fd_sc_hd__nand2_1
X_08721_ _08720_/B _08721_/B _08721_/C vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__nand3b_1
X_05933_ _05933_/A vssd1 vssd1 vccd1 vccd1 _05936_/B sky130_fd_sc_hd__inv_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _08652_/A _08652_/B _08652_/C vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__nand3_1
X_05864_ _06257_/B _06256_/A vssd1 vssd1 vccd1 vccd1 _05864_/Y sky130_fd_sc_hd__nor2_1
X_07603_ _07803_/B _07602_/Y vssd1 vssd1 vccd1 vccd1 _07721_/B sky130_fd_sc_hd__nor2b_1
XFILLER_0_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08583_ _08581_/Y _08307_/B _08582_/Y vssd1 vssd1 vccd1 vccd1 _08858_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05795_ _05795_/A vssd1 vssd1 vccd1 vccd1 _06268_/B sky130_fd_sc_hd__inv_2
XFILLER_0_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07534_ _07534_/A _07534_/B _07534_/C vssd1 vssd1 vccd1 vccd1 _07537_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07465_ _07537_/C vssd1 vssd1 vccd1 vccd1 _07536_/B sky130_fd_sc_hd__inv_2
X_09204_ _09204_/A _09204_/B vssd1 vssd1 vccd1 vccd1 _09205_/B sky130_fd_sc_hd__nand2_1
X_06416_ _06416_/A _06417_/A vssd1 vssd1 vccd1 vccd1 _06419_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07396_ _07385_/Y _07373_/B _07386_/Y vssd1 vssd1 vccd1 vccd1 _07397_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09135_ _09135_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09137_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06347_ _06756_/B _06755_/A vssd1 vssd1 vccd1 vccd1 _06759_/C sky130_fd_sc_hd__nand2_1
X_09066_ _09352_/B _09066_/B _09067_/B vssd1 vssd1 vccd1 vccd1 _09352_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06278_ _06313_/A _06313_/C vssd1 vssd1 vccd1 vccd1 _06311_/A sky130_fd_sc_hd__nand2_1
X_08017_ _08017_/A _08017_/B vssd1 vssd1 vccd1 vccd1 _08018_/B sky130_fd_sc_hd__nand2_1
X_05229_ input7/X vssd1 vssd1 vccd1 vccd1 _09496_/B sky130_fd_sc_hd__buf_8
X_09968_ _09958_/Y _09968_/B _09968_/C vssd1 vssd1 vccd1 vccd1 _09973_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__10485__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _09981_/A input17/X vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__nand2_1
X_09899_ _09897_/Y _09899_/B vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10108_ _10131_/B _10131_/C vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__nand2_1
X_10039_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05235__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05580_ input4/X _08272_/B vssd1 vssd1 vccd1 vccd1 _06065_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07250_ _07474_/A _07475_/C vssd1 vssd1 vccd1 vccd1 _07250_/Y sky130_fd_sc_hd__nand2_1
X_07181_ _07181_/A _07181_/B _07181_/C vssd1 vssd1 vccd1 vccd1 _07182_/B sky130_fd_sc_hd__nand3_1
X_06201_ _06201_/A _06201_/B vssd1 vssd1 vccd1 vccd1 _06628_/B sky130_fd_sc_hd__nand2_1
X_06132_ _06585_/A _06134_/A _06134_/B vssd1 vssd1 vccd1 vccd1 _06166_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06063_ _06063_/A _06063_/B _06063_/C vssd1 vssd1 vccd1 vccd1 _06064_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_39_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09822_ _09821_/B _09822_/B _09975_/B vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__nand3b_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _09751_/Y _09753_/B vssd1 vssd1 vccd1 vccd1 _09754_/B sky130_fd_sc_hd__and2b_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _08725_/C _08901_/B vssd1 vssd1 vccd1 vccd1 _08723_/A sky130_fd_sc_hd__nand2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _06965_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06968_/B sky130_fd_sc_hd__nand2_1
X_09684_ _10026_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10051__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05916_ _05916_/A _05916_/B _05916_/C vssd1 vssd1 vccd1 vccd1 _06316_/C sky130_fd_sc_hd__nand3_1
X_06896_ _06885_/C _06885_/B _06895_/Y vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08635_ _08635_/A _08635_/B _08635_/C vssd1 vssd1 vccd1 vccd1 _08642_/C sky130_fd_sc_hd__nand3_1
X_05847_ _10051_/B _07216_/B vssd1 vssd1 vccd1 vccd1 _06223_/C sky130_fd_sc_hd__nand2_1
X_08566_ _10051_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _08567_/C sky130_fd_sc_hd__nand2_1
X_07517_ _07534_/A _07533_/A vssd1 vssd1 vccd1 vccd1 _07517_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05778_ _05890_/B _05776_/Y _05777_/Y vssd1 vssd1 vccd1 vccd1 _05781_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ _08498_/B _08498_/A vssd1 vssd1 vccd1 vccd1 _08499_/A sky130_fd_sc_hd__or2_1
XANTENNA__05799__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07448_ _07448_/A _07448_/B _07448_/C vssd1 vssd1 vccd1 vccd1 _07451_/C sky130_fd_sc_hd__nand3_1
X_07379_ _07380_/B _07380_/A vssd1 vssd1 vccd1 vccd1 _07410_/A sky130_fd_sc_hd__nor2_2
X_09118_ _09118_/A vssd1 vssd1 vccd1 vccd1 _09119_/C sky130_fd_sc_hd__inv_2
X_10390_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__nand2_1
X_09049_ _09049_/A _09049_/B vssd1 vssd1 vccd1 vccd1 _09049_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06423__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09750__A _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10500__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06750_ _06750_/A _06750_/B _06750_/C vssd1 vssd1 vccd1 vccd1 _06751_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07164__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05701_ _09199_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _05706_/B sky130_fd_sc_hd__nand2_1
X_06681_ _06899_/C _06681_/B vssd1 vssd1 vccd1 vccd1 _06784_/B sky130_fd_sc_hd__nand2_1
X_08420_ _08420_/A input17/X vssd1 vssd1 vccd1 vccd1 _08425_/A sky130_fd_sc_hd__nand2_1
X_05632_ _05404_/Y _05905_/B _05496_/Y vssd1 vssd1 vccd1 vccd1 _05633_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08276__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05563_ _05563_/A vssd1 vssd1 vccd1 vccd1 _05564_/C sky130_fd_sc_hd__inv_2
X_08282_ _08510_/B _08283_/A vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05494_ _05494_/A _05494_/B vssd1 vssd1 vccd1 vccd1 _05906_/C sky130_fd_sc_hd__nand2_1
X_07302_ _07366_/B _07302_/B vssd1 vssd1 vccd1 vccd1 _07313_/A sky130_fd_sc_hd__nand2_1
X_07233_ _07235_/A _07236_/B vssd1 vssd1 vccd1 vccd1 _07234_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07164_ _09022_/C _08689_/A vssd1 vssd1 vccd1 vccd1 _07171_/A sky130_fd_sc_hd__nand2_1
X_06115_ _06534_/B _06119_/C vssd1 vssd1 vccd1 vccd1 _06117_/A sky130_fd_sc_hd__nand2_1
X_07095_ _07120_/B _07120_/C vssd1 vssd1 vccd1 vccd1 _07119_/A sky130_fd_sc_hd__nand2_1
X_06046_ _06046_/A _06046_/B vssd1 vssd1 vccd1 vccd1 _06049_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_10_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09805_ _09805_/A _09953_/A _09953_/B _09953_/C vssd1 vssd1 vccd1 vccd1 _09957_/B
+ sky130_fd_sc_hd__or4_1
X_07997_ _08866_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__nand2_1
X_09736_ _10134_/A vssd1 vssd1 vccd1 vccd1 _09737_/B sky130_fd_sc_hd__inv_2
X_06948_ _06948_/A _06959_/B vssd1 vssd1 vccd1 vccd1 _06951_/A sky130_fd_sc_hd__nand2_1
X_09667_ _09666_/B _09667_/B _09682_/B vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__nand3b_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08618_/A _08618_/B vssd1 vssd1 vccd1 vccd1 _08621_/C sky130_fd_sc_hd__nand2_1
X_06879_ _06879_/A _06879_/B vssd1 vssd1 vccd1 vccd1 _06885_/A sky130_fd_sc_hd__nand2_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09598_/A vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__inv_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08810_/B vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05322__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _10511_/CLK hold4/X fanout99/A vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ _10442_/A vssd1 vssd1 vccd1 vccd1 _10442_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10373_ hold1/X _10373_/B vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09464__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08824__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07920_ _10405_/B _10406_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08077_/A sky130_fd_sc_hd__o21ai_1
X_07851_ _07851_/A vssd1 vssd1 vccd1 vccd1 _07851_/Y sky130_fd_sc_hd__inv_2
X_07782_ _07789_/A _07806_/B _07790_/B vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__nand3_1
X_06802_ _06831_/A _06836_/B vssd1 vssd1 vccd1 vccd1 _06802_/Y sky130_fd_sc_hd__nor2_1
Xinput2 a_i[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_09521_ _09523_/A vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__inv_2
XANTENNA__09390__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06733_ _06733_/A _06805_/A vssd1 vssd1 vccd1 vccd1 _06839_/C sky130_fd_sc_hd__nand2_1
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09477_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06664_ _10043_/B _09981_/B vssd1 vssd1 vccd1 vccd1 _06769_/A sky130_fd_sc_hd__nand2_1
X_09383_ _09382_/B _09383_/B _09383_/C vssd1 vssd1 vccd1 vccd1 _09388_/B sky130_fd_sc_hd__nand3b_1
X_08403_ _08404_/B _08404_/A vssd1 vssd1 vccd1 vccd1 _08630_/B sky130_fd_sc_hd__or2_1
X_06595_ _06098_/B _06098_/C _06594_/Y vssd1 vssd1 vccd1 vccd1 _06598_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__05423__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05615_ _06169_/B _05615_/B vssd1 vssd1 vccd1 vccd1 _05620_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ _10050_/A _10111_/B vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__nand2_1
X_05546_ _05546_/A _05546_/B vssd1 vssd1 vccd1 vccd1 _06043_/B sky130_fd_sc_hd__nand2_1
X_08265_ _08265_/A vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05477_ input36/X _08810_/B vssd1 vssd1 vccd1 vccd1 _05479_/B sky130_fd_sc_hd__nand2_1
X_08196_ _08196_/A _08196_/B _08196_/C _08196_/D vssd1 vssd1 vccd1 vccd1 _08197_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07216_ _09361_/C _07216_/B vssd1 vssd1 vccd1 vccd1 _07217_/A sky130_fd_sc_hd__nand2_1
X_07147_ _07148_/B _07147_/B _07147_/C vssd1 vssd1 vccd1 vccd1 _07154_/B sky130_fd_sc_hd__nand3b_4
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07078_ _07092_/B _07078_/B _07081_/A vssd1 vssd1 vccd1 vccd1 _07092_/A sky130_fd_sc_hd__nand3_1
X_06029_ _06029_/A _06029_/B vssd1 vssd1 vccd1 vccd1 _06457_/B sky130_fd_sc_hd__nand2_1
X_09719_ _09728_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09719_/X sky130_fd_sc_hd__and2_1
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10425_ _10428_/B _10425_/B vssd1 vssd1 vccd1 vccd1 _10469_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10356_ _10357_/B _10357_/A vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__nor2_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ hold82/X _10287_/B vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05400_ _05400_/A _05400_/B vssd1 vssd1 vccd1 vccd1 _05916_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08554__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06380_ _06380_/A _06380_/B vssd1 vssd1 vccd1 vccd1 _06381_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05331_ _05331_/A _05331_/B _05331_/C vssd1 vssd1 vccd1 vccd1 _05332_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _08056_/B _08053_/C vssd1 vssd1 vccd1 vccd1 _08059_/B sky130_fd_sc_hd__nand2_1
X_05262_ _05262_/A _05262_/B _05262_/C vssd1 vssd1 vccd1 vccd1 _05286_/C sky130_fd_sc_hd__nand3_1
X_07001_ _07001_/A _07001_/B vssd1 vssd1 vccd1 vccd1 _07004_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08952_ _08952_/A _08952_/B _09306_/B vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__nand3_1
X_08883_ _08886_/C _08886_/B vssd1 vssd1 vccd1 vccd1 _08884_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06521__B _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ _07907_/B _07903_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10043__B _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _07942_/B _07832_/Y _07833_/Y vssd1 vssd1 vccd1 vccd1 _07846_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07765_ _07765_/A _07765_/B vssd1 vssd1 vccd1 vccd1 _07770_/C sky130_fd_sc_hd__nand2_1
X_09504_ _09829_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09510_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07696_ _07700_/C _07700_/B vssd1 vssd1 vccd1 vccd1 _07699_/A sky130_fd_sc_hd__nand2_1
X_06716_ _06716_/A _06716_/B _06716_/C vssd1 vssd1 vccd1 vccd1 _06805_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09435_ _09272_/B _09434_/Y _09270_/Y vssd1 vssd1 vccd1 vccd1 _09802_/A sky130_fd_sc_hd__a21oi_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06647_ _06363_/Y _06746_/B _06372_/Y vssd1 vssd1 vccd1 vccd1 _06735_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09366_ input51/X _10112_/B vssd1 vssd1 vccd1 vccd1 _09369_/B sky130_fd_sc_hd__nand2_1
X_06578_ _06579_/B _06579_/A vssd1 vssd1 vccd1 vccd1 _06578_/Y sky130_fd_sc_hd__nand2_1
X_09297_ _09297_/A vssd1 vssd1 vccd1 vccd1 _09298_/B sky130_fd_sc_hd__inv_2
X_08317_ _08317_/A _08317_/B vssd1 vssd1 vccd1 vccd1 _08319_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05529_ _06037_/A _06037_/B vssd1 vssd1 vccd1 vccd1 _05534_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08248_ _09962_/B _08248_/B vssd1 vssd1 vccd1 vccd1 _08250_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08179_ _08179_/A _08188_/B vssd1 vssd1 vccd1 vccd1 _08189_/B sky130_fd_sc_hd__and2_1
XFILLER_0_15_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10210_ _10485_/Q hold70/X vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__or2_1
XANTENNA__09295__A _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _10141_/A vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10072_ _10072_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09755__A2 _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ _10407_/B _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__a21bo_1
X_10339_ _10339_/A hold6/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__nand2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08549__A _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05880_ _05880_/A _05880_/B vssd1 vssd1 vccd1 vccd1 _06219_/C sky130_fd_sc_hd__nand2_1
X_07550_ _08811_/B _09751_/A _07553_/A vssd1 vssd1 vccd1 vccd1 _07733_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06501_ _06501_/A _08281_/A _06501_/C vssd1 vssd1 vccd1 vccd1 _06502_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09220_ _09528_/A _09685_/A _09684_/B _09533_/B vssd1 vssd1 vccd1 vccd1 _09526_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07481_ _07483_/A _07483_/C vssd1 vssd1 vccd1 vccd1 _07482_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06432_ _06432_/A _06432_/B vssd1 vssd1 vccd1 vccd1 _06432_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _09162_/A _09161_/A vssd1 vssd1 vccd1 vccd1 _09151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06363_ _06744_/A _06739_/A vssd1 vssd1 vccd1 vccd1 _06363_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05701__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ _09083_/A _09856_/D _09083_/C vssd1 vssd1 vccd1 vccd1 _09082_/Y sky130_fd_sc_hd__o21ai_1
X_08102_ _08102_/A _08004_/X vssd1 vssd1 vccd1 vccd1 _08103_/B sky130_fd_sc_hd__nor2b_1
X_05314_ _05246_/C _05246_/B _05311_/Y vssd1 vssd1 vccd1 vccd1 _05328_/B sky130_fd_sc_hd__a21o_1
X_08033_ _08134_/B _08033_/B vssd1 vssd1 vccd1 vccd1 _08039_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06294_ _09685_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _06295_/C sky130_fd_sc_hd__nand2_1
Xinput60 b_i[5] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
X_05245_ _05311_/A _05311_/B vssd1 vssd1 vccd1 vccd1 _05246_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__xor2_1
X_08935_ _09963_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09562__B _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ input51/X _08866_/B vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__nand2_1
X_08797_ _08797_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08806_/A sky130_fd_sc_hd__nand2_1
X_07817_ _07817_/A _07817_/B vssd1 vssd1 vccd1 vccd1 _07819_/B sky130_fd_sc_hd__nand2_1
X_07748_ _07748_/A vssd1 vssd1 vccd1 vccd1 _07767_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07679_ _07679_/A _07679_/B vssd1 vssd1 vccd1 vccd1 _07681_/A sky130_fd_sc_hd__nand2_1
X_09418_ _09418_/A _09418_/B vssd1 vssd1 vccd1 vccd1 _09421_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09349_ _09349_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09985__A2 _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06442__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ _10124_/A _10124_/B _10124_/C vssd1 vssd1 vccd1 vccd1 _10128_/C sky130_fd_sc_hd__nand3_1
X_10055_ _10055_/A _10056_/A vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _06981_/A vssd1 vssd1 vccd1 vccd1 _07400_/A sky130_fd_sc_hd__inv_2
X_08720_ _08720_/A _08720_/B vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__nand2_1
X_05932_ _05936_/A _05933_/A vssd1 vssd1 vccd1 vccd1 _05935_/A sky130_fd_sc_hd__nand2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _08651_/A _08651_/B vssd1 vssd1 vccd1 vccd1 _08657_/A sky130_fd_sc_hd__nand2_1
X_05863_ _06258_/C vssd1 vssd1 vccd1 vccd1 _06260_/B sky130_fd_sc_hd__inv_2
XANTENNA__07183__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _07602_/A _07602_/B vssd1 vssd1 vccd1 vccd1 _07602_/Y sky130_fd_sc_hd__nand2_1
X_08582_ _08582_/A _08582_/B vssd1 vssd1 vccd1 vccd1 _08582_/Y sky130_fd_sc_hd__nor2_1
X_05794_ _09960_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _05795_/A sky130_fd_sc_hd__nand2_1
X_07533_ _07533_/A _07533_/B vssd1 vssd1 vccd1 vccd1 _07537_/A sky130_fd_sc_hd__nand2_1
X_07464_ _07464_/A _07520_/A vssd1 vssd1 vccd1 vccd1 _07537_/C sky130_fd_sc_hd__nand2_1
X_09203_ _09204_/B _09204_/A vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06415_ _09962_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _06417_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09134_ _09424_/B _09134_/B _09134_/C vssd1 vssd1 vccd1 vccd1 _09155_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_60_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07395_ _07624_/A _07395_/B vssd1 vssd1 vccd1 vccd1 _07631_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08742__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06346_ _09496_/B _09988_/A vssd1 vssd1 vccd1 vccd1 _06755_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _09065_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _09067_/B sky130_fd_sc_hd__nand2_1
X_06277_ _06277_/A _06277_/B _06277_/C vssd1 vssd1 vccd1 vccd1 _06313_/C sky130_fd_sc_hd__nand3_1
X_08016_ _08032_/C vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__inv_2
X_05228_ _05337_/A _05338_/A vssd1 vssd1 vccd1 vccd1 _05291_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09968_/C sky130_fd_sc_hd__nand2_1
X_08918_ _09981_/B _09998_/B vssd1 vssd1 vccd1 vccd1 _09289_/C sky130_fd_sc_hd__nand2_1
X_09898_ _09898_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _09899_/B sky130_fd_sc_hd__nand2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _08849_/A _08850_/A vssd1 vssd1 vccd1 vccd1 _09141_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09748__A _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07969__A1 _09392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07268__A _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10107_ _10107_/A _10107_/B _10107_/C vssd1 vssd1 vccd1 vccd1 _10131_/C sky130_fd_sc_hd__nand3_1
X_10038_ _10022_/Y _10023_/X _10037_/Y vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05235__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06200_ _06628_/A _06201_/A _06201_/B vssd1 vssd1 vccd1 vccd1 _06208_/A sky130_fd_sc_hd__nand3_1
X_07180_ _07180_/A _07180_/B vssd1 vssd1 vccd1 vccd1 _07181_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06131_ _06131_/A _06131_/B _06131_/C vssd1 vssd1 vccd1 vccd1 _06134_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06062_ _06062_/A vssd1 vssd1 vccd1 vccd1 _06063_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09821_ _09821_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__nand2_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09752_ _09751_/A _09751_/B _09751_/C vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__o21ai_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _08703_/A _08703_/B _08927_/A vssd1 vssd1 vccd1 vccd1 _08901_/B sky130_fd_sc_hd__nand3_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _06964_/A _06983_/A vssd1 vssd1 vccd1 vccd1 _06965_/A sky130_fd_sc_hd__nand2_1
X_09683_ _09683_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09929_/B sky130_fd_sc_hd__and2_1
XANTENNA__10051__B _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05915_ _05915_/A _05915_/B vssd1 vssd1 vccd1 vccd1 _06316_/B sky130_fd_sc_hd__nand2_1
X_06895_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _06895_/Y sky130_fd_sc_hd__nor2_1
X_08634_ _08634_/A _08634_/B vssd1 vssd1 vccd1 vccd1 _08642_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05846_ _06221_/A _06222_/A vssd1 vssd1 vccd1 vccd1 _05851_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08565_ _10050_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _08870_/A sky130_fd_sc_hd__nand2_1
X_05777_ _05887_/A _05888_/B vssd1 vssd1 vccd1 vccd1 _05777_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07516_ _07533_/A _07534_/A vssd1 vssd1 vccd1 vccd1 _07516_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08496_ _08790_/C _08496_/B vssd1 vssd1 vccd1 vccd1 _08498_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ _07447_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07378_ _07378_/A _07378_/B vssd1 vssd1 vccd1 vccd1 _07380_/A sky130_fd_sc_hd__and2_1
X_09117_ _09117_/A _09118_/A vssd1 vssd1 vccd1 vccd1 _09120_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06329_ _06331_/A _06331_/B vssd1 vssd1 vccd1 vccd1 _06330_/A sky130_fd_sc_hd__nand2_1
X_09048_ _09049_/B _09049_/A vssd1 vssd1 vccd1 vccd1 _09048_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09325__B1 _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07551__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05700_ input42/X vssd1 vssd1 vccd1 vccd1 _09199_/A sky130_fd_sc_hd__buf_4
X_06680_ _06681_/B _06680_/B _06680_/C vssd1 vssd1 vccd1 vccd1 _06899_/C sky130_fd_sc_hd__nand3_1
X_05631_ _05631_/A _05631_/B vssd1 vssd1 vccd1 vccd1 _05977_/B sky130_fd_sc_hd__nand2_1
X_08350_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08537_/B sky130_fd_sc_hd__or2_1
XANTENNA__08276__B _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07301_ _07366_/A vssd1 vssd1 vccd1 vccd1 _07302_/B sky130_fd_sc_hd__inv_2
X_05562_ _05562_/A _06087_/A _06043_/A vssd1 vssd1 vccd1 vccd1 _05564_/B sky130_fd_sc_hd__nand3_1
X_08281_ _08281_/A _08281_/B vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05493_ _05493_/A _05493_/B _05493_/C vssd1 vssd1 vccd1 vccd1 _05494_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10475__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07232_ _07235_/B vssd1 vssd1 vccd1 vccd1 _07236_/B sky130_fd_sc_hd__inv_2
XFILLER_0_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07163_ _09022_/D _08688_/A vssd1 vssd1 vccd1 vccd1 _07170_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06114_ _06114_/A _06114_/B vssd1 vssd1 vccd1 vccd1 _06119_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07094_ _07094_/A _07094_/B vssd1 vssd1 vccd1 vccd1 _07120_/C sky130_fd_sc_hd__nand2_1
X_06045_ _06044_/B _06045_/B _06045_/C vssd1 vssd1 vccd1 vccd1 _06046_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09804_ _09804_/A vssd1 vssd1 vccd1 vccd1 _09953_/B sky130_fd_sc_hd__inv_2
XFILLER_0_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07996_ _09890_/D _09762_/A _07994_/C vssd1 vssd1 vccd1 vccd1 _08000_/C sky130_fd_sc_hd__o21ai_1
X_09735_ _09510_/A _09511_/C _09516_/A vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__o21a_1
X_06947_ _06949_/B _06949_/C vssd1 vssd1 vccd1 vccd1 _06959_/B sky130_fd_sc_hd__nand2_1
X_09666_ _09666_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _08618_/B _08618_/A vssd1 vssd1 vccd1 vccd1 _08886_/B sky130_fd_sc_hd__or2_1
X_06878_ _06895_/B vssd1 vssd1 vccd1 vccd1 _06879_/B sky130_fd_sc_hd__inv_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ input49/X input50/X _10083_/B _09854_/B vssd1 vssd1 vccd1 vccd1 _09598_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05829_ _05829_/A _05829_/B vssd1 vssd1 vccd1 vccd1 _05830_/A sky130_fd_sc_hd__nand2_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08548_ _08579_/A _08579_/B vssd1 vssd1 vccd1 vccd1 _08578_/A sky130_fd_sc_hd__nand2_1
X_08479_ _10027_/B _09953_/A _08479_/C vssd1 vssd1 vccd1 vccd1 _08480_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ _10511_/CLK hold22/X fanout99/A vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _10473_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _10372_/A vssd1 vssd1 vccd1 vccd1 _10508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07265__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09761__A _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08824__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07456__A _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _07855_/A _07855_/B vssd1 vssd1 vccd1 vccd1 _07853_/A sky130_fd_sc_hd__nand2_1
X_07781_ _07789_/C vssd1 vssd1 vccd1 vccd1 _07806_/B sky130_fd_sc_hd__inv_2
X_06801_ _06836_/B _06831_/A vssd1 vssd1 vccd1 vccd1 _06801_/Y sky130_fd_sc_hd__nand2_1
X_09520_ _09520_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__nand2_1
X_06732_ _06732_/A _06805_/B _06732_/C vssd1 vssd1 vccd1 vccd1 _06805_/A sky130_fd_sc_hd__nand3_1
Xinput3 a_i[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08287__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05704__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _09451_/A _09451_/B _09451_/C vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__nand3_1
X_06663_ _06782_/B _06782_/C vssd1 vssd1 vccd1 vccd1 _06781_/A sky130_fd_sc_hd__nand2_1
X_09382_ _09382_/A _09382_/B vssd1 vssd1 vccd1 vccd1 _09388_/A sky130_fd_sc_hd__nand2_1
X_08402_ _08623_/B _08402_/B vssd1 vssd1 vccd1 vccd1 _08404_/A sky130_fd_sc_hd__nand2_1
X_06594_ _06594_/A _06594_/B vssd1 vssd1 vccd1 vccd1 _06594_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05614_ _05614_/A _05614_/B vssd1 vssd1 vccd1 vccd1 _05615_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05423__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08333_ _08345_/C vssd1 vssd1 vccd1 vccd1 _08333_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05545_ _05547_/B vssd1 vssd1 vccd1 vccd1 _05546_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08264_ _08264_/A _08265_/A vssd1 vssd1 vccd1 vccd1 _08314_/A sky130_fd_sc_hd__nand2_1
X_05476_ input37/X _08814_/B vssd1 vssd1 vccd1 vccd1 _05479_/A sky130_fd_sc_hd__nand2_1
X_08195_ _10385_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08196_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_6_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07215_ _07218_/A _07218_/B vssd1 vssd1 vccd1 vccd1 _07272_/A sky130_fd_sc_hd__nand2_1
X_07146_ _07146_/A _07146_/B _07146_/C vssd1 vssd1 vccd1 vccd1 _07151_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07077_ _07209_/B _07077_/B vssd1 vssd1 vccd1 vccd1 _07081_/A sky130_fd_sc_hd__nand2_1
X_06028_ _06030_/B vssd1 vssd1 vccd1 vccd1 _06029_/B sky130_fd_sc_hd__inv_2
X_09718_ _09728_/B _09728_/A vssd1 vssd1 vccd1 vccd1 _09718_/Y sky130_fd_sc_hd__nor2_1
X_07979_ _07980_/B _08034_/A vssd1 vssd1 vccd1 vccd1 _08037_/B sky130_fd_sc_hd__nand2_1
X_09649_ _09649_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09652_/C sky130_fd_sc_hd__nor2_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10424_ _10424_/A _10428_/A vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10355_ hold49/X vssd1 vssd1 vccd1 vccd1 _10357_/B sky130_fd_sc_hd__inv_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10287_/B hold82/X vssd1 vssd1 vccd1 vccd1 _10293_/A sky130_fd_sc_hd__or2_1
XFILLER_0_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08554__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05330_ _05330_/A vssd1 vssd1 vccd1 vccd1 _05331_/C sky130_fd_sc_hd__inv_2
XFILLER_0_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05261_ _05503_/A _05503_/B vssd1 vssd1 vccd1 vccd1 _05262_/C sky130_fd_sc_hd__nand2_1
X_07000_ _07000_/A vssd1 vssd1 vccd1 vccd1 _07001_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08951_ _08951_/A vssd1 vssd1 vccd1 vccd1 _08952_/A sky130_fd_sc_hd__inv_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07186__A _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ _08878_/Y _08882_/B _08882_/C vssd1 vssd1 vccd1 vccd1 _08885_/B sky130_fd_sc_hd__nand3b_1
X_07902_ _07902_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _07903_/B sky130_fd_sc_hd__nor2_1
X_07833_ _07833_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _07833_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08729__B _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07764_ _07784_/B _07784_/A vssd1 vssd1 vccd1 vccd1 _07925_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _09503_/A _09503_/B _09503_/C vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07695_ _07695_/A _07695_/B vssd1 vssd1 vccd1 vccd1 _07700_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06715_ _06715_/A _06715_/B vssd1 vssd1 vccd1 vccd1 _06732_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _09434_/A vssd1 vssd1 vccd1 vccd1 _09434_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06646_ _06646_/A _06646_/B _06646_/C vssd1 vssd1 vccd1 vccd1 _06654_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08745__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09365_ _09369_/A vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06577_ _06583_/A _06583_/C vssd1 vssd1 vccd1 vccd1 _06582_/A sky130_fd_sc_hd__nand2_1
X_09296_ _09777_/A _09953_/C _09296_/C vssd1 vssd1 vccd1 vccd1 _09298_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08316_ _08521_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08597_/B sky130_fd_sc_hd__nand2_1
X_05528_ _05528_/A _05528_/B vssd1 vssd1 vccd1 vccd1 _05534_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08247_ _09960_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _08250_/A sky130_fd_sc_hd__nand2_1
X_05459_ _05732_/B _05459_/B vssd1 vssd1 vccd1 vccd1 _05493_/B sky130_fd_sc_hd__nand2_1
X_08178_ _10387_/B _10391_/A vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07129_ _07133_/A _07133_/B vssd1 vssd1 vccd1 vccd1 _07627_/B sky130_fd_sc_hd__xor2_2
X_10140_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__nor2_1
X_10071_ _10070_/B _10071_/B _10071_/C vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08390__A _08390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10407_ _10407_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10464_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10338_ _10336_/Y _10338_/B vssd1 vssd1 vccd1 vccd1 _10340_/A sky130_fd_sc_hd__and2b_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _10249_/B _10266_/B _10267_/B _10251_/Y _10260_/B vssd1 vssd1 vccd1 vccd1
+ hold104/A sky130_fd_sc_hd__a221oi_2
XFILLER_0_17_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06500_ _06500_/A _06500_/B vssd1 vssd1 vccd1 vccd1 _06502_/A sky130_fd_sc_hd__nand2_1
X_07480_ _07480_/A vssd1 vssd1 vccd1 vccd1 _07483_/A sky130_fd_sc_hd__inv_2
XANTENNA__08565__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06431_ _06436_/C _08225_/A vssd1 vssd1 vccd1 vccd1 _06435_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _09150_/A _09150_/B vssd1 vssd1 vccd1 vccd1 _09171_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05701__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06362_ _06742_/B _06742_/C _06361_/Y vssd1 vssd1 vccd1 vccd1 _06739_/A sky130_fd_sc_hd__a21oi_1
X_09081_ _10083_/B vssd1 vssd1 vccd1 vccd1 _09856_/D sky130_fd_sc_hd__inv_2
XFILLER_0_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06293_ _08862_/B vssd1 vssd1 vccd1 vccd1 _09392_/C sky130_fd_sc_hd__inv_2
X_08101_ _08147_/B _08147_/A _08098_/X vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05313_ _05576_/B _05576_/A vssd1 vssd1 vccd1 vccd1 _05327_/A sky130_fd_sc_hd__nand2_1
X_08032_ _08033_/B _08032_/B _08032_/C vssd1 vssd1 vccd1 vccd1 _08134_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_44_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05244_ _05244_/A vssd1 vssd1 vccd1 vccd1 _05246_/B sky130_fd_sc_hd__inv_2
Xinput50 b_i[25] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_4
XFILLER_0_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput61 b_i[6] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09983_ _09981_/X _09983_/B vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05429__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ _08947_/B vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__inv_2
XANTENNA__09562__C _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _09071_/B _08868_/C vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__nand2_1
X_08796_ _08800_/B _08796_/B vssd1 vssd1 vccd1 vccd1 _08797_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08182__A2 _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ _07816_/A _07816_/B _07816_/C vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07747_ _07749_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07748_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _08207_/B _07676_/Y _07677_/Y vssd1 vssd1 vccd1 vccd1 _07678_/Y sky130_fd_sc_hd__o21ai_1
X_09417_ _09421_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06629_ _06627_/Y _06207_/A _06628_/Y vssd1 vssd1 vccd1 vccd1 _06638_/A sky130_fd_sc_hd__a21oi_2
X_09348_ _09348_/A _09349_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_35_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09279_ _09278_/B _09279_/B vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07996__A2 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06723__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06442__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _10110_/A _09897_/Y _09899_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10054_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05802__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _07399_/B _07399_/A vssd1 vssd1 vccd1 vccd1 _06981_/A sky130_fd_sc_hd__nor2_1
X_05931_ _05934_/B vssd1 vssd1 vccd1 vccd1 _05936_/A sky130_fd_sc_hd__inv_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ _09180_/B _08660_/C vssd1 vssd1 vccd1 vccd1 _08659_/A sky130_fd_sc_hd__nand2_1
X_05862_ input35/X _09560_/B vssd1 vssd1 vccd1 vccd1 _06258_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07183__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ _07602_/B _07602_/A vssd1 vssd1 vccd1 vccd1 _07803_/B sky130_fd_sc_hd__nor2_1
X_08581_ _08582_/B _08582_/A vssd1 vssd1 vccd1 vccd1 _08581_/Y sky130_fd_sc_hd__nand2_1
X_05793_ _05796_/A _05796_/B vssd1 vssd1 vccd1 vccd1 _06268_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07532_ _07534_/A vssd1 vssd1 vccd1 vccd1 _07533_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07463_ _07520_/B _07463_/B _07463_/C vssd1 vssd1 vccd1 vccd1 _07520_/A sky130_fd_sc_hd__nand3_1
X_09202_ _09555_/B _09202_/B vssd1 vssd1 vccd1 vccd1 _09204_/A sky130_fd_sc_hd__nand2_1
X_06414_ _08255_/B _06418_/C vssd1 vssd1 vccd1 vccd1 _06416_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09133_ _09137_/C vssd1 vssd1 vccd1 vccd1 _09134_/C sky130_fd_sc_hd__inv_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ _07631_/A _07624_/A _07395_/B vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08742__B _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06345_ _10026_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _06756_/B sky130_fd_sc_hd__nand2_2
X_09064_ _08771_/B _08772_/B _08900_/B vssd1 vssd1 vccd1 vccd1 _09065_/B sky130_fd_sc_hd__a21boi_1
X_06276_ _06276_/A _06276_/B vssd1 vssd1 vccd1 vccd1 _06313_/A sky130_fd_sc_hd__nand2_1
X_08015_ _08017_/B _08017_/A vssd1 vssd1 vccd1 vccd1 _08032_/C sky130_fd_sc_hd__nor2_2
X_05227_ _05347_/C _05347_/B _05226_/Y vssd1 vssd1 vccd1 vccd1 _05338_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__09854__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09966_ _09958_/Y _09959_/X _09968_/B vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__o21bai_1
X_09897_ _10109_/B _09898_/A vssd1 vssd1 vccd1 vccd1 _09897_/Y sky130_fd_sc_hd__nor2_1
X_08917_ _08917_/A vssd1 vssd1 vccd1 vccd1 _08922_/B sky130_fd_sc_hd__inv_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08848_ _08848_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08850_/A sky130_fd_sc_hd__nand2_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08779_ input3/X vssd1 vssd1 vccd1 vccd1 _09710_/D sky130_fd_sc_hd__inv_2
XFILLER_0_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07969__A2 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__A _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07268__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10470__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__nand2_1
X_10037_ _10041_/A _10041_/B vssd1 vssd1 vccd1 vccd1 _10037_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06130_ _06130_/A vssd1 vssd1 vccd1 vccd1 _06131_/C sky130_fd_sc_hd__inv_2
XFILLER_0_14_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06061_ _06061_/A _06062_/A vssd1 vssd1 vccd1 vccd1 _06064_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__xor2_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09751_ _09751_/A _09751_/B _09751_/C vssd1 vssd1 vccd1 vccd1 _09751_/Y sky130_fd_sc_hd__nor3_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06963_ _06963_/A vssd1 vssd1 vccd1 vccd1 _06983_/A sky130_fd_sc_hd__inv_2
X_08702_ _08702_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _08725_/C sky130_fd_sc_hd__nand2_1
X_05914_ _05916_/A _05916_/B vssd1 vssd1 vccd1 vccd1 _05915_/A sky130_fd_sc_hd__nand2_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ _09682_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__and2_1
X_06894_ _06899_/B _06899_/C vssd1 vssd1 vccd1 vccd1 _06943_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08633_ _08635_/C vssd1 vssd1 vccd1 vccd1 _08634_/B sky130_fd_sc_hd__inv_2
XFILLER_0_55_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05845_ _06221_/B vssd1 vssd1 vccd1 vccd1 _06222_/A sky130_fd_sc_hd__inv_2
X_08564_ _08575_/B _08575_/C vssd1 vssd1 vccd1 vccd1 _08573_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05776_ _05888_/B _05887_/A vssd1 vssd1 vccd1 vccd1 _05776_/Y sky130_fd_sc_hd__nand2_1
X_07515_ _07505_/Y _07544_/B _07514_/Y vssd1 vssd1 vccd1 vccd1 _07534_/A sky130_fd_sc_hd__a21oi_2
X_08495_ _09963_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _08496_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07446_ _07448_/B vssd1 vssd1 vccd1 vccd1 _07447_/B sky130_fd_sc_hd__inv_2
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07377_ _07377_/A _07377_/B vssd1 vssd1 vccd1 vccd1 _07378_/B sky130_fd_sc_hd__or2_1
X_09116_ _09119_/A _09418_/B vssd1 vssd1 vccd1 vccd1 _09117_/A sky130_fd_sc_hd__nand2_1
X_06328_ _06328_/A _06328_/B _06328_/C vssd1 vssd1 vccd1 vccd1 _06331_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09047_ _09053_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _09399_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06259_ _06259_/A _06259_/B vssd1 vssd1 vccd1 vccd1 _06260_/A sky130_fd_sc_hd__nand2_1
X_09949_ _09971_/B _09971_/A vssd1 vssd1 vccd1 vccd1 _09949_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09325__B2 _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09325__A1 _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07551__B input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05352__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05630_ _05977_/A _05631_/A _05631_/B vssd1 vssd1 vccd1 vccd1 _05785_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07300_ _07323_/C _07323_/B _07321_/A vssd1 vssd1 vccd1 vccd1 _07366_/A sky130_fd_sc_hd__a21oi_2
X_05561_ _06087_/B _05561_/B vssd1 vssd1 vccd1 vccd1 _05564_/A sky130_fd_sc_hd__nand2_1
X_08280_ _08489_/A _08284_/C vssd1 vssd1 vccd1 vccd1 _08510_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05492_ _05492_/A vssd1 vssd1 vccd1 vccd1 _05493_/C sky130_fd_sc_hd__inv_2
X_07231_ _07236_/A vssd1 vssd1 vccd1 vccd1 _07235_/A sky130_fd_sc_hd__inv_2
X_07162_ _07162_/A _07162_/B vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__nand2_1
X_06113_ _06113_/A _06113_/B vssd1 vssd1 vccd1 vccd1 _06534_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07093_ _07093_/A _07093_/B vssd1 vssd1 vccd1 vccd1 _07094_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06044_ _06044_/A _06044_/B vssd1 vssd1 vccd1 vccd1 _06046_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09803_ _09951_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09809_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05437__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ _07995_/A vssd1 vssd1 vccd1 vccd1 _08014_/B sky130_fd_sc_hd__inv_2
X_09734_ _09738_/A _09738_/B vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06946_ _06946_/A _06946_/B _06946_/C vssd1 vssd1 vccd1 vccd1 _06949_/C sky130_fd_sc_hd__nand3_1
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__nor2_1
X_06877_ _10043_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _06895_/B sky130_fd_sc_hd__nand2_1
X_08616_ _08345_/C _08345_/B _08331_/Y vssd1 vssd1 vccd1 vccd1 _08618_/A sky130_fd_sc_hd__a21oi_1
X_05828_ _05960_/B _05960_/C vssd1 vssd1 vccd1 vccd1 _05959_/A sky130_fd_sc_hd__nand2_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09212_/B _10050_/A _10083_/B _09210_/X vssd1 vssd1 vccd1 vccd1 _09873_/A
+ sky130_fd_sc_hd__a31o_1
X_08547_ _08547_/A _08547_/B _08547_/C vssd1 vssd1 vccd1 vccd1 _08579_/B sky130_fd_sc_hd__nand3_1
X_05759_ _05759_/A vssd1 vssd1 vccd1 vccd1 _05879_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ input7/X _09313_/D vssd1 vssd1 vccd1 vccd1 _08479_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07429_ _07482_/B vssd1 vssd1 vccd1 vccd1 _07483_/B sky130_fd_sc_hd__inv_2
X_10440_ _10440_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10441_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07099__A _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ _10368_/Y _10373_/B vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09489__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08393__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07737__A _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ _07806_/A _07789_/C vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__nand2_1
X_06800_ _06834_/B _06834_/C _06799_/Y vssd1 vssd1 vccd1 vccd1 _06831_/A sky130_fd_sc_hd__a21oi_1
X_06731_ _06965_/B vssd1 vssd1 vccd1 vccd1 _06732_/C sky130_fd_sc_hd__inv_2
Xinput4 a_i[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
X_09450_ _09825_/B vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08401_ _08401_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _08402_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05704__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06662_ _06662_/A _06662_/B _06662_/C vssd1 vssd1 vccd1 vccd1 _06782_/B sky130_fd_sc_hd__nand3_1
Xclkbuf_2_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10495_/CLK sky130_fd_sc_hd__clkbuf_16
X_09381_ _09381_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09382_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06593_ _08317_/A _06598_/C vssd1 vssd1 vccd1 vccd1 _06599_/A sky130_fd_sc_hd__nand2_1
X_05613_ _06093_/A _05613_/B vssd1 vssd1 vccd1 vccd1 _06169_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08332_ _08332_/A _08332_/B vssd1 vssd1 vccd1 vccd1 _08345_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_46_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05544_ input7/X _08248_/B vssd1 vssd1 vccd1 vccd1 _05547_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08263_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07214_ _08814_/B _08248_/B vssd1 vssd1 vccd1 vccd1 _07218_/B sky130_fd_sc_hd__nand2_1
X_05475_ _05826_/A _05825_/B _05826_/B vssd1 vssd1 vccd1 vccd1 _05490_/B sky130_fd_sc_hd__nand3_1
X_08194_ _08194_/A _08194_/B vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__nand2_1
X_07145_ _07689_/A _07690_/A vssd1 vssd1 vccd1 vccd1 _07707_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06551__A _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07076_ _07077_/B _07076_/B _07076_/C vssd1 vssd1 vccd1 vccd1 _07209_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07787__B1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06027_ input8/X _08248_/B vssd1 vssd1 vccd1 vccd1 _06030_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07978_ _08027_/B _08026_/C _07977_/Y vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__a21oi_2
X_09717_ _09717_/A vssd1 vssd1 vccd1 vccd1 _09728_/A sky130_fd_sc_hd__inv_2
X_06929_ _06929_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _06930_/A sky130_fd_sc_hd__nand2_1
X_09648_ _09648_/A vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__inv_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09579_ _09741_/A _09579_/B _09910_/A vssd1 vssd1 vccd1 vccd1 _09583_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ _10423_/A vssd1 vssd1 vccd1 vccd1 _10468_/D sky130_fd_sc_hd__clkbuf_1
X_10354_ hold65/X vssd1 vssd1 vccd1 vccd1 _10504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ _10278_/A hold32/X _10277_/B hold81/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__a31o_1
XANTENNA__10465__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__A_N _10171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09455__B1 _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05260_ _05265_/C vssd1 vssd1 vccd1 vccd1 _05262_/B sky130_fd_sc_hd__inv_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08950_ _08950_/A _08951_/A vssd1 vssd1 vccd1 vccd1 _08955_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07186__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _08885_/A sky130_fd_sc_hd__nand2_1
X_07901_ _07910_/B _08055_/A vssd1 vssd1 vccd1 vccd1 _08064_/C sky130_fd_sc_hd__nand2_1
X_07832_ _07944_/B vssd1 vssd1 vccd1 vccd1 _07832_/Y sky130_fd_sc_hd__inv_2
X_09502_ _09503_/A _09503_/C _09503_/B vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07763_ _07763_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07694_ _07694_/A _07703_/A vssd1 vssd1 vccd1 vccd1 _10417_/A sky130_fd_sc_hd__nand2_1
X_06714_ _06716_/A vssd1 vssd1 vccd1 vccd1 _06715_/B sky130_fd_sc_hd__inv_2
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06645_ _06820_/A _06820_/C vssd1 vssd1 vccd1 vccd1 _06818_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09364_ _09608_/B _09364_/B vssd1 vssd1 vccd1 vccd1 _09369_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08745__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06546__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ _08315_/A _08315_/B _08315_/C vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__nand3_1
X_06576_ _06576_/A _06576_/B _06576_/C vssd1 vssd1 vccd1 vccd1 _06583_/C sky130_fd_sc_hd__nand3_1
X_09295_ _09437_/B vssd1 vssd1 vccd1 vccd1 _09953_/C sky130_fd_sc_hd__inv_2
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05527_ _06037_/B vssd1 vssd1 vccd1 vccd1 _05528_/B sky130_fd_sc_hd__inv_2
X_08246_ _09816_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__nand2_1
X_05458_ _05399_/C _05457_/Y _05395_/B vssd1 vssd1 vccd1 vccd1 _05459_/B sky130_fd_sc_hd__o21ai_1
X_08177_ _08177_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__nand2_1
X_07128_ _07094_/B _07091_/A _07121_/A vssd1 vssd1 vccd1 vccd1 _07133_/B sky130_fd_sc_hd__o21a_1
X_05389_ input4/X _08248_/B vssd1 vssd1 vccd1 vccd1 _05392_/B sky130_fd_sc_hd__nand2_1
X_07059_ _07347_/A _07345_/A vssd1 vssd1 vccd1 vccd1 _07059_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10488__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10072_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10495__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10406_ _10406_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10463_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10337_ _10501_/Q _10479_/Q vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ hold91/A vssd1 vssd1 vccd1 vccd1 _10268_/Y sky130_fd_sc_hd__inv_2
X_10199_ _10199_/A hold18/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08565__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06430_ _06429_/B _08225_/B _06430_/C vssd1 vssd1 vccd1 vccd1 _08225_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05270__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06361_ _06750_/A _06749_/A vssd1 vssd1 vccd1 vccd1 _06361_/Y sky130_fd_sc_hd__nor2_1
X_09080_ _09087_/A _09087_/B vssd1 vssd1 vccd1 vccd1 _09085_/A sky130_fd_sc_hd__nand2_1
X_08100_ _08098_/X _08100_/B vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05312_ _05246_/C _05246_/B _05311_/Y vssd1 vssd1 vccd1 vccd1 _05576_/A sky130_fd_sc_hd__a21oi_1
X_06292_ _09528_/A vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__inv_2
Xinput40 b_i[16] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_2
X_08031_ _08031_/A _08031_/B vssd1 vssd1 vccd1 vccd1 _08032_/B sky130_fd_sc_hd__nand2_1
X_05243_ _05243_/A _05243_/B vssd1 vssd1 vccd1 vccd1 _05246_/A sky130_fd_sc_hd__nand2_1
Xinput51 b_i[26] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_4
Xinput62 b_i[7] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09982_ _09981_/A input21/X _09981_/B input20/X vssd1 vssd1 vccd1 vccd1 _09983_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05429__B _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ _08933_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _08947_/B sky130_fd_sc_hd__nand2_2
XANTENNA__09562__D _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _10084_/A _09890_/D _08863_/C vssd1 vssd1 vccd1 vccd1 _08868_/C sky130_fd_sc_hd__o21ai_1
X_08795_ _08798_/B _08798_/C vssd1 vssd1 vccd1 vccd1 _08797_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05445__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ _07815_/A _07815_/B _07815_/C vssd1 vssd1 vccd1 vccd1 _07921_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_79_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07746_ _08825_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _07749_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _09415_/B _09416_/B _09658_/A vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__nand3b_1
X_07677_ _08203_/B _07677_/B vssd1 vssd1 vccd1 vccd1 _07677_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06628_ _06628_/A _06628_/B vssd1 vssd1 vccd1 vccd1 _06628_/Y sky130_fd_sc_hd__nor2_1
X_09347_ _09346_/B _09347_/B _09520_/A vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__nand3b_2
X_06559_ _10050_/A input1/X vssd1 vssd1 vccd1 vccd1 _06560_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09278_ _09279_/B _09278_/B vssd1 vssd1 vccd1 vccd1 _09479_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ _08240_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06723__B _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ _10109_/X _10110_/Y _10121_/Y vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10053_ _10053_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07554__B _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10503__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05802__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09497__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06633__B _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07745__A _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05930_ _06328_/B _06328_/C vssd1 vssd1 vccd1 vccd1 _06327_/A sky130_fd_sc_hd__nand2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09960__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05861_ _06257_/B _06256_/A vssd1 vssd1 vccd1 vccd1 _06260_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08580_ _08586_/B _08586_/C vssd1 vssd1 vccd1 vccd1 _08858_/B sky130_fd_sc_hd__nand2_1
X_07600_ _07600_/A _07600_/B vssd1 vssd1 vccd1 vccd1 _07602_/A sky130_fd_sc_hd__and2_1
XFILLER_0_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07531_ _07531_/A _07906_/A vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__nand2_1
X_05792_ _09963_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _05796_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ _07462_/A _07599_/A vssd1 vssd1 vccd1 vccd1 _07464_/A sky130_fd_sc_hd__nand2_1
X_09201_ _09199_/A _10052_/A _09548_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _09202_/B
+ sky130_fd_sc_hd__a22o_1
X_06413_ _06413_/A _06413_/B vssd1 vssd1 vccd1 vccd1 _06418_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_8_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07393_ _07393_/A _07393_/B _07393_/C vssd1 vssd1 vccd1 vccd1 _07395_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ _09132_/A _09132_/B vssd1 vssd1 vccd1 vccd1 _09137_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06344_ _06750_/B _06750_/C vssd1 vssd1 vccd1 vccd1 _06749_/A sky130_fd_sc_hd__nand2_1
X_09063_ _09063_/A _09345_/A vssd1 vssd1 vccd1 vccd1 _09065_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06275_ _06277_/C vssd1 vssd1 vccd1 vccd1 _06276_/B sky130_fd_sc_hd__inv_2
X_08014_ _08014_/A _08014_/B vssd1 vssd1 vccd1 vccd1 _08017_/A sky130_fd_sc_hd__and2_1
XFILLER_0_12_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05226_ _05344_/B _05343_/A vssd1 vssd1 vccd1 vccd1 _05226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09854__B _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09965_ _09965_/A _09965_/B vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__xor2_1
X_09896_ _09896_/A vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__inv_2
X_08916_ _09980_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__nand2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08847_ _08846_/B _08847_/B _08847_/C vssd1 vssd1 vccd1 vccd1 _08848_/B sky130_fd_sc_hd__nand3b_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08778_ _08899_/B _08851_/B vssd1 vssd1 vccd1 vccd1 _08849_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07729_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07730_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07549__B input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10105_ _10107_/C vssd1 vssd1 vccd1 vccd1 _10106_/B sky130_fd_sc_hd__inv_2
X_10036_ _10035_/B _10036_/B _10036_/C vssd1 vssd1 vccd1 vccd1 _10041_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_81_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09020__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06060_ _09960_/A _09022_/D vssd1 vssd1 vccd1 vccd1 _06062_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _09987_/A input22/X vssd1 vssd1 vccd1 vccd1 _09751_/C sky130_fd_sc_hd__nand2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06962_ _06962_/A _06962_/B vssd1 vssd1 vccd1 vccd1 _06964_/A sky130_fd_sc_hd__nand2_1
X_09681_ _09681_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _10457_/B sky130_fd_sc_hd__nand2_1
X_08701_ _08703_/A vssd1 vssd1 vccd1 vccd1 _08702_/B sky130_fd_sc_hd__inv_2
X_05913_ _05913_/A _05913_/B vssd1 vssd1 vccd1 vccd1 _05916_/B sky130_fd_sc_hd__nand2_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08632_ _08632_/A _09150_/A vssd1 vssd1 vccd1 vccd1 _08635_/C sky130_fd_sc_hd__nand2_1
X_06893_ _06893_/A _06893_/B _06893_/C vssd1 vssd1 vccd1 vccd1 _06899_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05844_ _10043_/B _08248_/B vssd1 vssd1 vccd1 vccd1 _06221_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06819__A _07709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08563_ _08563_/A _08563_/B vssd1 vssd1 vccd1 vccd1 _08575_/C sky130_fd_sc_hd__nand2_1
XANTENNA__05723__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05775_ _05814_/B _05814_/C _05774_/Y vssd1 vssd1 vccd1 vccd1 _05887_/A sky130_fd_sc_hd__a21oi_2
X_08494_ _09962_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _08790_/C sky130_fd_sc_hd__nand2_1
X_07514_ _07539_/A _07542_/A vssd1 vssd1 vccd1 vccd1 _07514_/Y sky130_fd_sc_hd__nor2_1
X_07445_ _07454_/B vssd1 vssd1 vccd1 vccd1 _07452_/A sky130_fd_sc_hd__inv_2
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07376_ _07382_/B _07382_/A vssd1 vssd1 vccd1 vccd1 _07527_/B sky130_fd_sc_hd__nand2_1
X_09115_ _09115_/A _09115_/B _09406_/A vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06327_ _06327_/A _06327_/B vssd1 vssd1 vccd1 vccd1 _06331_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09046_ _09046_/A _09046_/B _09046_/C vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__nand3_1
X_06258_ _06258_/A _06258_/B _06258_/C vssd1 vssd1 vccd1 vccd1 _06264_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05209_ _05216_/A _05251_/B vssd1 vssd1 vccd1 vccd1 _05215_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06189_ _06634_/B vssd1 vssd1 vccd1 vccd1 _06635_/C sky130_fd_sc_hd__inv_2
X_09948_ _09835_/A _09835_/B _10019_/B vssd1 vssd1 vccd1 vccd1 _10017_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09325__A2 _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09880_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_99_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05352__B _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09775__A _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07295__A _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ _10019_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10020_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07878__A2 _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05560_ _05560_/A _05560_/B _05563_/A vssd1 vssd1 vccd1 vccd1 _05565_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05491_ _05491_/A _05492_/A vssd1 vssd1 vccd1 vccd1 _05494_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07230_ _07417_/B _07417_/C vssd1 vssd1 vccd1 vccd1 _07416_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07161_ _07160_/Y _06640_/B _06640_/A vssd1 vssd1 vccd1 vccd1 _07162_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__09685__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06112_ _06114_/B vssd1 vssd1 vccd1 vccd1 _06113_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ _07092_/A _07092_/B vssd1 vssd1 vccd1 vccd1 _07094_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06043_ _06043_/A _06043_/B vssd1 vssd1 vccd1 vccd1 _06044_/B sky130_fd_sc_hd__nand2_1
X_09802_ _09802_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__nor2_1
XANTENNA__05437__B _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07994_ _09890_/D _09762_/A _07994_/C vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__nor3_1
X_09733_ _09733_/A _09733_/B _09733_/C vssd1 vssd1 vccd1 vccd1 _09738_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06945_ _06959_/A vssd1 vssd1 vccd1 vccd1 _06948_/A sky130_fd_sc_hd__inv_2
X_09664_ _09664_/A vssd1 vssd1 vccd1 vccd1 _09665_/B sky130_fd_sc_hd__inv_2
XFILLER_0_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06876_ _06895_/A vssd1 vssd1 vccd1 vccd1 _06879_/A sky130_fd_sc_hd__inv_2
XFILLER_0_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09595_ _09215_/B _09593_/X _09594_/Y vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__o21ba_1
X_08615_ _08881_/B _08615_/B vssd1 vssd1 vccd1 vccd1 _08618_/B sky130_fd_sc_hd__nand2_1
X_05827_ _05827_/A _05827_/B _05827_/C vssd1 vssd1 vccd1 vccd1 _05960_/C sky130_fd_sc_hd__nand3_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ _08546_/A _08546_/B vssd1 vssd1 vccd1 vccd1 _08579_/A sky130_fd_sc_hd__nand2_1
X_05758_ input38/X _09361_/C vssd1 vssd1 vccd1 vccd1 _05759_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08477_ input8/X vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__inv_2
X_05689_ _06175_/A _06133_/A _05690_/B vssd1 vssd1 vccd1 vccd1 _05729_/A sky130_fd_sc_hd__nand3_1
XANTENNA__06284__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07428_ _10083_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _07482_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07359_ _07359_/A _07359_/B vssd1 vssd1 vccd1 vccd1 _07359_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07099__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ _10376_/B hold69/X _10376_/C vssd1 vssd1 vccd1 vccd1 _10373_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ _09356_/B _09030_/A vssd1 vssd1 vccd1 vccd1 _09042_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07309__A1 _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09489__B _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ _10509_/CLK hold16/X fanout100/X vssd1 vssd1 vccd1 vccd1 _10499_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07737__B input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07456__C _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06730_ _06730_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06733_/A sky130_fd_sc_hd__nand2_1
Xinput5 a_i[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XFILLER_0_36_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06661_ _06661_/A _06661_/B vssd1 vssd1 vccd1 vccd1 _06662_/B sky130_fd_sc_hd__nand2_1
X_08400_ _08401_/B _08401_/A vssd1 vssd1 vccd1 vccd1 _08623_/B sky130_fd_sc_hd__or2_1
X_05612_ _06169_/A _06093_/A _05613_/B vssd1 vssd1 vccd1 vccd1 _05620_/A sky130_fd_sc_hd__nand3_1
X_09380_ _09383_/B _09383_/C vssd1 vssd1 vccd1 vccd1 _09382_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09549__D_N _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06592_ _06600_/C vssd1 vssd1 vccd1 vccd1 _06597_/B sky130_fd_sc_hd__inv_2
XFILLER_0_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ _08332_/B _08332_/A vssd1 vssd1 vccd1 vccd1 _08331_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05543_ _05547_/A vssd1 vssd1 vccd1 vccd1 _05546_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08262_ _08261_/B _08262_/B _08262_/C vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05474_ _05826_/C vssd1 vssd1 vccd1 vccd1 _05825_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07213_ _08825_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _07218_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08193_ _10385_/B vssd1 vssd1 vccd1 vccd1 _08196_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07144_ _07684_/B _07684_/A vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07787__A1 _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07075_ _07206_/B _07205_/B vssd1 vssd1 vccd1 vccd1 _07076_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07787__B2 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06026_ _06030_/A vssd1 vssd1 vccd1 vccd1 _06029_/A sky130_fd_sc_hd__inv_2
X_07977_ _08024_/A _08023_/A vssd1 vssd1 vccd1 vccd1 _07977_/Y sky130_fd_sc_hd__nor2_1
X_09716_ _09716_/A _09716_/B vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__nand2_1
X_06928_ _06928_/A _06928_/B _06928_/C vssd1 vssd1 vccd1 vccd1 _06934_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08478__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09649_/A sky130_fd_sc_hd__nor2_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ _06862_/B vssd1 vssd1 vccd1 vccd1 _06864_/A sky130_fd_sc_hd__inv_2
X_09578_ _09910_/B _09578_/B vssd1 vssd1 vccd1 vccd1 _09583_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08494__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08529_/A vssd1 vssd1 vccd1 vccd1 _08531_/B sky130_fd_sc_hd__inv_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07838__A _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ _10422_/A _10424_/A vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__and2_1
X_10353_ hold64/X _10357_/A vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__and2_1
XFILLER_0_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10284_ _10298_/B vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__inv_2
XFILLER_0_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06917__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09455__A1 _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09963__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08880_ _08878_/Y _08882_/C vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__nand2b_1
X_07900_ _07907_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__nand2_1
X_07831_ _09361_/C _08214_/A vssd1 vssd1 vccd1 vccd1 _07944_/B sky130_fd_sc_hd__nand2_1
X_09501_ _09501_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _09503_/B sky130_fd_sc_hd__xnor2_1
X_07762_ _07808_/A _07809_/C vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__nand2_1
X_07693_ _07693_/A _07693_/B _07700_/B vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06713_ _06684_/Y _06796_/B _06712_/Y vssd1 vssd1 vccd1 vccd1 _06716_/A sky130_fd_sc_hd__a21o_1
X_09432_ _09432_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _10450_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06644_ _06644_/A _07153_/A vssd1 vssd1 vccd1 vccd1 _06820_/A sky130_fd_sc_hd__nand2_2
X_09363_ input49/X _09854_/B input50/X _09601_/B vssd1 vssd1 vccd1 vccd1 _09364_/B
+ sky130_fd_sc_hd__a22o_1
X_06575_ _06575_/A _06575_/B vssd1 vssd1 vccd1 vccd1 _06583_/A sky130_fd_sc_hd__nand2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06546__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _08314_/A _08314_/B _08314_/C vssd1 vssd1 vccd1 vccd1 _08315_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05526_ _09962_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _06037_/B sky130_fd_sc_hd__nand2_1
X_09294_ _09447_/A _09294_/B _09507_/A vssd1 vssd1 vccd1 vccd1 _09300_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08245_ _08266_/A _08266_/C vssd1 vssd1 vccd1 vccd1 _08264_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05457_ _05397_/A _05397_/C _05396_/B vssd1 vssd1 vccd1 vccd1 _05457_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06562__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _08176_/A _08176_/B _08176_/C vssd1 vssd1 vccd1 vccd1 _08177_/B sky130_fd_sc_hd__nand3_1
X_05388_ _05392_/A vssd1 vssd1 vccd1 vccd1 _05391_/A sky130_fd_sc_hd__inv_2
XFILLER_0_27_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07127_ _07127_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _07133_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ _07195_/B _07195_/C _07057_/Y vssd1 vssd1 vccd1 vccd1 _07345_/A sky130_fd_sc_hd__a21oi_1
X_06009_ _06451_/A _06013_/C vssd1 vssd1 vccd1 vccd1 _06011_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_0__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ _10405_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10406_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10336_ _10501_/Q _10479_/Q vssd1 vssd1 vccd1 vccd1 _10336_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10267_/A _10267_/B vssd1 vssd1 vccd1 vccd1 _10267_/Y sky130_fd_sc_hd__nand2_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10198_ _10196_/Y hold95/A vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08862__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06360_ _06751_/C vssd1 vssd1 vccd1 vccd1 _06742_/C sky130_fd_sc_hd__inv_2
XANTENNA__05270__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05311_ _05311_/A _05311_/B vssd1 vssd1 vccd1 vccd1 _05311_/Y sky130_fd_sc_hd__nor2_1
X_06291_ _06291_/A _06291_/B vssd1 vssd1 vccd1 vccd1 _06303_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08030_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _08031_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 a_i[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
X_05242_ _05242_/A _05242_/B _05244_/A vssd1 vssd1 vccd1 vccd1 _05247_/A sky130_fd_sc_hd__nand3_1
Xinput52 b_i[27] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_4
Xinput41 b_i[17] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
Xinput63 b_i[8] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09981_ _09981_/A _09981_/B input20/X input21/X vssd1 vssd1 vccd1 vccd1 _09981_/X
+ sky130_fd_sc_hd__and4_1
X_08932_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _08948_/B sky130_fd_sc_hd__and2_1
X_08863_ _10084_/A _09890_/D _08863_/C vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__or3_1
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08794_ _08794_/A _08995_/A _09014_/A vssd1 vssd1 vccd1 vccd1 _08798_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_74_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05445__B _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07814_ _07817_/B _07816_/B _07816_/C vssd1 vssd1 vccd1 vccd1 _07815_/A sky130_fd_sc_hd__nand3_1
X_07745_ _09361_/C _08688_/A vssd1 vssd1 vccd1 vccd1 _07749_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09415_ _09415_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07676_ _07677_/B _08203_/B vssd1 vssd1 vccd1 vccd1 _07676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06627_ _06628_/B _06628_/A vssd1 vssd1 vccd1 vccd1 _06627_/Y sky130_fd_sc_hd__nand2_1
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09349_/A sky130_fd_sc_hd__nand2_1
X_06558_ input48/X vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__clkbuf_4
X_09277_ _09277_/A _09277_/B vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__nand2_1
X_06489_ _06490_/A _06490_/B vssd1 vssd1 vccd1 vccd1 _08356_/B sky130_fd_sc_hd__or2_1
XFILLER_0_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05509_ _09951_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _05998_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08228_/A _08228_/B _08228_/C vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06292__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08159_ _08186_/A _10383_/C _10383_/B vssd1 vssd1 vccd1 vccd1 _08188_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10121_ _10124_/A _10124_/C vssd1 vssd1 vccd1 vccd1 _10121_/Y sky130_fd_sc_hd__nand2_1
X_10052_ _10052_/A input46/X vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07554__C _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09497__B _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10436__B _10437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10319_ _10319_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10325_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07745__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__B _10171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09960__B _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05860_ _10050_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _06256_/A sky130_fd_sc_hd__nand2_2
X_05791_ input36/X vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__clkbuf_8
X_07530_ _07530_/A _07614_/B _07614_/A vssd1 vssd1 vccd1 vccd1 _07906_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_44_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07461_ _07463_/C vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__inv_2
X_09200_ _09200_/A vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__inv_2
XANTENNA__10478__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06412_ _09951_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _06413_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07392_ _07392_/A _07392_/B _07392_/C vssd1 vssd1 vccd1 vccd1 _07393_/B sky130_fd_sc_hd__nand3_1
X_09131_ _09135_/A _09136_/A vssd1 vssd1 vccd1 vccd1 _09134_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06343_ _06343_/A _06343_/B _06343_/C vssd1 vssd1 vccd1 vccd1 _06750_/C sky130_fd_sc_hd__nand3_1
X_09062_ _09068_/B vssd1 vssd1 vccd1 vccd1 _09066_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06274_ _06246_/Y _06380_/B _06273_/Y vssd1 vssd1 vccd1 vccd1 _06277_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08013_ _08866_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _08017_/B sky130_fd_sc_hd__nand2_1
X_05225_ _05345_/C vssd1 vssd1 vccd1 vccd1 _05347_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09964_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09965_/B sky130_fd_sc_hd__xnor2_1
X_09895_ _10117_/A _10109_/C vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__nand2_1
X_08915_ _08925_/B _09277_/B vssd1 vssd1 vccd1 vccd1 _08924_/A sky130_fd_sc_hd__nand2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _08846_/A _08846_/B vssd1 vssd1 vccd1 vccd1 _08848_/A sky130_fd_sc_hd__nand2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08851_/B sky130_fd_sc_hd__nand2_1
X_05989_ _06432_/B vssd1 vssd1 vccd1 vccd1 _05990_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07728_ _07728_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07731_/B sky130_fd_sc_hd__nand2_1
X_07659_ _07659_/A _07659_/B _07659_/C vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09329_ _09329_/A vssd1 vssd1 vccd1 vccd1 _09330_/B sky130_fd_sc_hd__inv_2
XFILLER_0_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08007__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10104_ _09876_/C _09876_/B _09872_/A vssd1 vssd1 vccd1 vccd1 _10107_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__05366__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ _10035_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09020__B _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06961_ _06968_/A vssd1 vssd1 vccd1 vccd1 _06967_/A sky130_fd_sc_hd__inv_2
X_09680_ _09676_/A _09679_/Y _09676_/B vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__a21boi_1
X_08700_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _08703_/A sky130_fd_sc_hd__nand2_1
X_05912_ _06328_/B _05912_/B vssd1 vssd1 vccd1 vccd1 _05913_/B sky130_fd_sc_hd__nand2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08631_ _08630_/B _09150_/B _08631_/C vssd1 vssd1 vccd1 vccd1 _09150_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__07491__A _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ _06892_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _06893_/B sky130_fd_sc_hd__nand2_1
X_05843_ _06222_/B vssd1 vssd1 vccd1 vccd1 _06221_/A sky130_fd_sc_hd__inv_2
X_08562_ _08563_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _08575_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__05723__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05774_ _05814_/A vssd1 vssd1 vccd1 vccd1 _05774_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08493_ _08493_/A vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__inv_2
X_07513_ _07545_/C vssd1 vssd1 vccd1 vccd1 _07544_/B sky130_fd_sc_hd__inv_2
X_07444_ _07432_/Y _07510_/B _07443_/Y vssd1 vssd1 vccd1 vccd1 _07454_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07375_ _07375_/A _07375_/B vssd1 vssd1 vccd1 vccd1 _07382_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09114_ _09114_/A _09114_/B vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06326_ _06739_/B _06326_/B vssd1 vssd1 vccd1 vccd1 _06327_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09045_ _09045_/A _09045_/B vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06257_ _06259_/B _06257_/B vssd1 vssd1 vccd1 vccd1 _06258_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05208_ _09963_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _05251_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06188_ _06190_/B _06190_/A vssd1 vssd1 vccd1 vccd1 _06634_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09947_ _09841_/A _09842_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10076_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09878_ _09878_/A vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__inv_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _08829_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09775__B _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07295__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _10018_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10020_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05490_ _05960_/B _05490_/B vssd1 vssd1 vccd1 vccd1 _05492_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07160_ _10434_/B vssd1 vssd1 vccd1 vccd1 _07160_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06111_ _09528_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _06114_/B sky130_fd_sc_hd__nand2_1
X_07091_ _07091_/A _07093_/A _07093_/B vssd1 vssd1 vccd1 vccd1 _07120_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06042_ _06045_/B _06045_/C vssd1 vssd1 vccd1 vccd1 _06044_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09801_ _09835_/B _10019_/B vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09732_ _09732_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09738_/A sky130_fd_sc_hd__nand2_1
X_07993_ _08862_/B _09981_/B vssd1 vssd1 vccd1 vccd1 _07994_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06944_ _06942_/Y _06910_/B _06943_/Y vssd1 vssd1 vccd1 vccd1 _06959_/A sky130_fd_sc_hd__a21oi_2
X_09663_ _09663_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__nor2_1
X_06875_ _10052_/A _08688_/A vssd1 vssd1 vccd1 vccd1 _06895_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09594_/Y sky130_fd_sc_hd__nor2_1
X_08614_ _08614_/A _08614_/B vssd1 vssd1 vccd1 vccd1 _08615_/B sky130_fd_sc_hd__nand2_1
X_05826_ _05826_/A _05826_/B _05826_/C vssd1 vssd1 vccd1 vccd1 _05827_/C sky130_fd_sc_hd__nand3_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _08547_/B vssd1 vssd1 vccd1 vccd1 _08546_/B sky130_fd_sc_hd__inv_2
XFILLER_0_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05757_ _05760_/A _05760_/B vssd1 vssd1 vccd1 vccd1 _05879_/C sky130_fd_sc_hd__nand2_1
X_08476_ _08476_/A _08476_/B _08673_/A vssd1 vssd1 vccd1 vccd1 _08672_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_64_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05688_ _05688_/A _05688_/B _05688_/C vssd1 vssd1 vccd1 vccd1 _05690_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06284__B _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07427_ _07430_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07483_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_45_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07358_ _07363_/B _07363_/C vssd1 vssd1 vccd1 vccd1 _07362_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06309_ _06309_/A _06309_/B vssd1 vssd1 vccd1 vccd1 _06716_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07289_ _07416_/A _07417_/A vssd1 vssd1 vccd1 vccd1 _07415_/B sky130_fd_sc_hd__nand2_1
X_09028_ _09028_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10489__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07309__A2 _09392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06475__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05819__A _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10498_ _10511_/CLK _10498_/D fanout100/X vssd1 vssd1 vccd1 vccd1 _10498_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07456__D _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 a_i[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06660_ _06660_/A _06660_/B vssd1 vssd1 vccd1 vccd1 _06662_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05611_ _05611_/A _05611_/B _05611_/C vssd1 vssd1 vccd1 vccd1 _05613_/B sky130_fd_sc_hd__nand3_1
X_06591_ _06591_/A _06591_/B vssd1 vssd1 vccd1 vccd1 _06600_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08330_ _08559_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08332_/A sky130_fd_sc_hd__xor2_1
X_05542_ _10026_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _05547_/A sky130_fd_sc_hd__nand2_1
X_08261_ _08261_/A _08261_/B vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05473_ _05825_/A _05826_/C vssd1 vssd1 vccd1 vccd1 _05489_/A sky130_fd_sc_hd__nand2_1
X_07212_ _07222_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07220_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08192_ _08192_/A vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__inv_2
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07143_ _07143_/A _07143_/B vssd1 vssd1 vccd1 vccd1 _07684_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08105__A _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _07207_/C vssd1 vssd1 vccd1 vccd1 _07076_/B sky130_fd_sc_hd__inv_2
XANTENNA__07787__A2 _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__RESET_B fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06025_ _09496_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _06030_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07976_ _08028_/B vssd1 vssd1 vccd1 vccd1 _08026_/C sky130_fd_sc_hd__inv_2
X_09715_ _10048_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09728_/B sky130_fd_sc_hd__nand2_1
X_06927_ _06929_/A _06927_/B vssd1 vssd1 vccd1 vccd1 _06928_/B sky130_fd_sc_hd__nand2_1
X_09646_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06858_ _07013_/B _07013_/C vssd1 vssd1 vccd1 vccd1 _07018_/A sky130_fd_sc_hd__nand2_1
X_09577_ _09910_/A vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08494__B _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _06779_/Y _06849_/B _06788_/Y vssd1 vssd1 vccd1 vccd1 _06842_/A sky130_fd_sc_hd__a21oi_1
X_05809_ _05809_/A _05809_/B _05809_/C vssd1 vssd1 vccd1 vccd1 _06298_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _10026_/A _09022_/D vssd1 vssd1 vccd1 vccd1 _08529_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06295__A _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08459_ _08463_/A _08719_/A vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07838__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _10427_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10424_/A sky130_fd_sc_hd__nand2_1
X_10352_ _10376_/B hold63/X vssd1 vssd1 vccd1 vccd1 _10357_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05639__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ _10283_/A _10283_/B vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06917__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05549__A _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__B _10175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__B _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07830_ _07833_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _07942_/B sky130_fd_sc_hd__nand2_1
X_07761_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07809_/C sky130_fd_sc_hd__xor2_1
X_09500_ _09500_/A _09692_/A vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__nand2_1
X_06712_ _06792_/A _06793_/B vssd1 vssd1 vccd1 vccd1 _06712_/Y sky130_fd_sc_hd__nor2_1
X_07692_ _07692_/A _07692_/B _07692_/C vssd1 vssd1 vccd1 vccd1 _07700_/B sky130_fd_sc_hd__nand3_1
X_09431_ _09431_/A _09431_/B _09674_/B vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06643_ _06643_/A _06643_/B _06643_/C vssd1 vssd1 vccd1 vccd1 _07153_/A sky130_fd_sc_hd__nand3_2
X_09362_ _09362_/A vssd1 vssd1 vccd1 vccd1 _09608_/B sky130_fd_sc_hd__inv_2
X_06574_ _06576_/A vssd1 vssd1 vccd1 vccd1 _06575_/B sky130_fd_sc_hd__inv_2
X_08313_ _08313_/A _08313_/B vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05525_ _08689_/A vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__buf_8
X_09293_ _09293_/A vssd1 vssd1 vccd1 vccd1 _09507_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08244_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08266_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05456_ _05617_/A _05456_/B vssd1 vssd1 vccd1 vccd1 _05732_/B sky130_fd_sc_hd__nand2_1
X_08175_ _08175_/A vssd1 vssd1 vccd1 vccd1 _08176_/A sky130_fd_sc_hd__inv_2
X_05387_ input3/X _08247_/B vssd1 vssd1 vccd1 vccd1 _05392_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06562__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07126_ _07126_/A _07400_/A vssd1 vssd1 vccd1 vccd1 _07127_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07057_ _07197_/A _07196_/A vssd1 vssd1 vccd1 vccd1 _07057_/Y sky130_fd_sc_hd__nor2_1
X_06008_ _06008_/A _06008_/B vssd1 vssd1 vccd1 vccd1 _06013_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07959_ _07959_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07963_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ input52/X input53/X _10112_/B _10111_/B vssd1 vssd1 vccd1 vccd1 _09629_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _10404_/A vssd1 vssd1 vccd1 vccd1 _10462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10335_ hold112/X vssd1 vssd1 vccd1 vccd1 _10500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07584__A _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10266_ _10266_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__and2_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10197_ _10483_/Q hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05832__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08862__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05310_ _05329_/A _05559_/A vssd1 vssd1 vccd1 vccd1 _05576_/B sky130_fd_sc_hd__nand2_1
X_06290_ _06296_/A vssd1 vssd1 vccd1 vccd1 _06291_/B sky130_fd_sc_hd__inv_2
Xinput20 a_i[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput31 a_i[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_1
X_05241_ _10026_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _05244_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput53 b_i[28] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_4
Xinput42 b_i[18] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_1
Xinput64 b_i[9] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09980_ _09980_/A input19/X vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__nand2_1
X_08931_ _08952_/B _09306_/B vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07494__A _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ input50/X _08862_/B vssd1 vssd1 vccd1 vccd1 _08863_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07813_ _07925_/C _07811_/Y _07925_/B vssd1 vssd1 vccd1 vccd1 _07817_/B sky130_fd_sc_hd__o21ai_1
X_08793_ _09014_/B _08793_/B vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07744_ _07743_/B _07744_/B _07744_/C vssd1 vssd1 vccd1 vccd1 _07821_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07675_ _07675_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _08203_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09414_ _09414_/A _09414_/B vssd1 vssd1 vccd1 vccd1 _09415_/B sky130_fd_sc_hd__and2_1
X_06626_ _06632_/B _06632_/C vssd1 vssd1 vccd1 vccd1 _06631_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09345_ _09345_/A _09345_/B vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__and2_1
X_06557_ _06571_/A _06570_/A vssd1 vssd1 vccd1 vccd1 _08399_/B sky130_fd_sc_hd__or2_1
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09276_ _09276_/A _09473_/A vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__nand2_1
X_06488_ _09963_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _06490_/B sky130_fd_sc_hd__nand2_1
X_05508_ _05998_/A vssd1 vssd1 vccd1 vccd1 _05517_/A sky130_fd_sc_hd__inv_2
X_08227_ _08227_/A _08227_/B vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__nand2_1
X_05439_ input36/X _09022_/D vssd1 vssd1 vccd1 vccd1 _05678_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08158_ _08112_/Y _08158_/B _08158_/C vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__nand3b_1
X_08089_ _08032_/C _08032_/B _08033_/B vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__a21boi_1
X_07109_ _07109_/A _07109_/B _07109_/C vssd1 vssd1 vccd1 vccd1 _07114_/B sky130_fd_sc_hd__nand3_1
X_10120_ _10120_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _10124_/C sky130_fd_sc_hd__nand2_1
XANTENNA_fanout99_A fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10051_ _10051_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _10053_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08963__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09497__C _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10318_ _10319_/B _10319_/A vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ _10249_/A _10249_/B vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__nor2_1
X_05790_ _09962_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _05796_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09034__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07460_ _07788_/A _07598_/A vssd1 vssd1 vccd1 vccd1 _07463_/C sky130_fd_sc_hd__nor2_1
XANTENNA__08609__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06411_ _06411_/A _09951_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__nand3_1
X_07391_ _07391_/A _07391_/B vssd1 vssd1 vccd1 vccd1 _07393_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ _08856_/Y _09143_/B _08897_/Y vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06342_ _06342_/A _06342_/B vssd1 vssd1 vccd1 vccd1 _06343_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ _09400_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _09068_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08012_ _08020_/B _08020_/A vssd1 vssd1 vccd1 vccd1 _08114_/B sky130_fd_sc_hd__nand2_1
X_06273_ _06377_/A _06376_/A vssd1 vssd1 vccd1 vccd1 _06273_/Y sky130_fd_sc_hd__nor2_1
X_05224_ input8/X input55/X vssd1 vssd1 vccd1 vccd1 _05345_/C sky130_fd_sc_hd__nand2_1
XANTENNA_fanout101_A input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09963_ _09963_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09964_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09209__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08914_ _08914_/A _08914_/B _09262_/A vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09888__A2 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ _09894_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _10109_/C sky130_fd_sc_hd__nand2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08547_/B _08546_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _08846_/B sky130_fd_sc_hd__o21ai_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _08517_/A _08516_/C _08672_/B vssd1 vssd1 vccd1 vccd1 _08777_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_79_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05988_ _08422_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _06432_/B sky130_fd_sc_hd__nand2_1
X_07727_ _07763_/B _07809_/B vssd1 vssd1 vccd1 vccd1 _07728_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07658_ _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__nand2_1
X_06609_ _06609_/A _06609_/B vssd1 vssd1 vccd1 vccd1 _06610_/B sky130_fd_sc_hd__nand2_1
X_07589_ _07770_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07592_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ _09320_/Y _09322_/Y _09329_/A vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _09260_/B _09260_/A vssd1 vssd1 vccd1 vccd1 _09265_/A sky130_fd_sc_hd__or2_1
XFILLER_0_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08007__B _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05647__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10103_ _10107_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10106_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10034_ _10034_/A _10034_/B vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07102__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06960_ _06958_/Y _06952_/B _06959_/Y vssd1 vssd1 vccd1 vccd1 _06968_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07772__A _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05911_ _05912_/B _05911_/B _05911_/C vssd1 vssd1 vccd1 vccd1 _06328_/B sky130_fd_sc_hd__nand3_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06891_ _06891_/A _06891_/B vssd1 vssd1 vccd1 vccd1 _06893_/A sky130_fd_sc_hd__nand2_1
X_08630_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _08632_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05842_ _08780_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _06222_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _08563_/B vssd1 vssd1 vccd1 vccd1 _08562_/B sky130_fd_sc_hd__inv_2
X_05773_ _05773_/A _05773_/B _05773_/C vssd1 vssd1 vccd1 vccd1 _05814_/A sky130_fd_sc_hd__nand3_1
X_08492_ input38/X input3/X vssd1 vssd1 vccd1 vccd1 _08493_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07512_ _07512_/A _07512_/B vssd1 vssd1 vccd1 vccd1 _07545_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07443_ _07508_/C _07507_/A vssd1 vssd1 vccd1 vccd1 _07443_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _09115_/A vssd1 vssd1 vccd1 vccd1 _09114_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07374_ _07374_/A _07374_/B _07374_/C vssd1 vssd1 vccd1 vccd1 _07375_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06325_ _06326_/B _06325_/B _06325_/C vssd1 vssd1 vccd1 vccd1 _06739_/B sky130_fd_sc_hd__nand3_1
X_09044_ _09046_/A vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__inv_2
XANTENNA__07947__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06256_ _06256_/A vssd1 vssd1 vccd1 vccd1 _06259_/B sky130_fd_sc_hd__inv_2
X_05207_ input33/X vssd1 vssd1 vccd1 vccd1 _08422_/A sky130_fd_sc_hd__buf_12
XFILLER_0_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05467__A _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06187_ _06187_/A _06187_/B vssd1 vssd1 vccd1 vccd1 _06190_/A sky130_fd_sc_hd__and2_1
X_09946_ _10176_/A _10176_/C vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09877_ _09878_/A _10100_/A _09877_/C vssd1 vssd1 vccd1 vccd1 _09880_/B sky130_fd_sc_hd__nand3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _08828_/A _08828_/B vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__nand2_1
X_08759_ _09049_/A vssd1 vssd1 vccd1 vccd1 _08760_/B sky130_fd_sc_hd__inv_2
XFILLER_0_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07857__A _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__A _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10468__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _10017_/A _10018_/B _10018_/A vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06639__C _06820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06110_ _06114_/A vssd1 vssd1 vccd1 vccd1 _06113_/A sky130_fd_sc_hd__inv_2
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07090_ _07090_/A _07090_/B _07090_/C vssd1 vssd1 vccd1 vccd1 _07093_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06041_ _06041_/A _06457_/A _06505_/A vssd1 vssd1 vccd1 vccd1 _06045_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ _09800_/A _09800_/B _09800_/C vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__nand3_2
X_07992_ _08689_/A vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__inv_2
X_09731_ _09733_/B vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__inv_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06943_ _06943_/A _06943_/B vssd1 vssd1 vccd1 vccd1 _06943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09662_ _09667_/B _09682_/B vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__nand2_1
X_06874_ _07023_/A _07024_/A vssd1 vssd1 vccd1 vccd1 _07016_/B sky130_fd_sc_hd__nand2_1
X_09593_ _09594_/B _09594_/A vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__and2_1
X_08613_ _08882_/B vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__inv_2
X_05825_ _05825_/A _05825_/B vssd1 vssd1 vccd1 vccd1 _05827_/A sky130_fd_sc_hd__nand2_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08544_ _08542_/Y _08362_/B _08543_/Y vssd1 vssd1 vccd1 vccd1 _08547_/B sky130_fd_sc_hd__a21oi_2
X_05756_ input36/X _09560_/B vssd1 vssd1 vccd1 vccd1 _05760_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08475_ _08475_/A _08475_/B vssd1 vssd1 vccd1 vccd1 _08517_/A sky130_fd_sc_hd__nand2_1
X_05687_ _05687_/A vssd1 vssd1 vccd1 vccd1 _05688_/C sky130_fd_sc_hd__inv_2
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07426_ _08810_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _07430_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09779__A1 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ _07357_/A _07357_/B vssd1 vssd1 vccd1 vccd1 _07363_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08780__B _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06308_ _06656_/C vssd1 vssd1 vccd1 vccd1 _06309_/B sky130_fd_sc_hd__inv_2
X_09027_ _09031_/A _09031_/C vssd1 vssd1 vccd1 vccd1 _09356_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07288_ _07264_/Y _07470_/B _07287_/Y vssd1 vssd1 vccd1 vccd1 _07417_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06239_ _10050_/B _07216_/B vssd1 vssd1 vccd1 vccd1 _06662_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09929_ _09929_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _09936_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06475__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08971__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10497_ _10509_/CLK hold12/X fanout100/X vssd1 vssd1 vccd1 vccd1 _10497_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05835__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 a_i[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05610_ _05610_/A _05610_/B _05610_/C vssd1 vssd1 vccd1 vccd1 _05611_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_86_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06590_ _06590_/A _06590_/B _06590_/C vssd1 vssd1 vccd1 vccd1 _06591_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05541_ _05573_/B _06022_/A _05572_/C vssd1 vssd1 vccd1 vccd1 _05571_/A sky130_fd_sc_hd__nand3_1
X_08260_ _08260_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08261_/B sky130_fd_sc_hd__nand2_1
X_05472_ _05871_/C _05871_/B _05471_/Y vssd1 vssd1 vccd1 vccd1 _05826_/C sky130_fd_sc_hd__a21oi_2
X_08191_ _08191_/A _10384_/B _08195_/B vssd1 vssd1 vccd1 vccd1 _08192_/A sky130_fd_sc_hd__nand3_1
X_07211_ _07359_/B _07359_/A vssd1 vssd1 vccd1 vccd1 _07222_/B sky130_fd_sc_hd__nand2_1
X_07142_ _07680_/A _07680_/B _07679_/B vssd1 vssd1 vccd1 vccd1 _07143_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09630__B1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07073_ _10083_/B _07216_/B vssd1 vssd1 vccd1 vccd1 _07207_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08105__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06024_ _06049_/A _06049_/B vssd1 vssd1 vccd1 vccd1 _06048_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07975_ _08038_/B _07975_/B vssd1 vssd1 vccd1 vccd1 _08028_/B sky130_fd_sc_hd__nand2_1
X_09714_ _09714_/A _09714_/B vssd1 vssd1 vccd1 vccd1 _09715_/B sky130_fd_sc_hd__nand2_1
X_06926_ _06926_/A vssd1 vssd1 vccd1 vccd1 _06929_/A sky130_fd_sc_hd__inv_2
X_09645_ _09917_/A _09931_/A _09645_/C vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_69_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07960__A _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06857_ _06857_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _07013_/C sky130_fd_sc_hd__nand3_1
X_05808_ _05808_/A vssd1 vssd1 vccd1 vccd1 _05809_/A sky130_fd_sc_hd__inv_2
X_09576_ _09574_/Y _09338_/B _09575_/Y vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__a21oi_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _06845_/A _06847_/B vssd1 vssd1 vccd1 vccd1 _06788_/Y sky130_fd_sc_hd__nor2_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08527_/A _08527_/B vssd1 vssd1 vccd1 vccd1 _08531_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06295__B _09392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05739_ _09199_/A _09548_/A _08862_/B input1/X vssd1 vssd1 vccd1 vccd1 _05740_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__09887__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08458_ _08719_/B _08458_/B _08458_/C vssd1 vssd1 vccd1 vccd1 _08719_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07409_ _07409_/A _07410_/A vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08389_ _08638_/B _08390_/A vssd1 vssd1 vccd1 vccd1 _08411_/B sky130_fd_sc_hd__nand2_1
X_10420_ _10421_/B _10427_/A vssd1 vssd1 vccd1 vccd1 _10422_/A sky130_fd_sc_hd__or2_1
XFILLER_0_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ hold63/X _10376_/B vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10282_ hold28/X vssd1 vssd1 vccd1 vccd1 _10283_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05655__A _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05549__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07760_ _07809_/A _07809_/B vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06711_ _06703_/A _06702_/A _06949_/B vssd1 vssd1 vccd1 vccd1 _06796_/B sky130_fd_sc_hd__o21ai_1
X_09430_ _09430_/A vssd1 vssd1 vccd1 vccd1 _09431_/B sky130_fd_sc_hd__inv_2
XFILLER_0_78_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07691_ _07691_/A _07691_/B vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06642_ _06816_/B vssd1 vssd1 vccd1 vccd1 _06643_/A sky130_fd_sc_hd__inv_2
X_09361_ input49/X input50/X _09361_/C _09361_/D vssd1 vssd1 vccd1 vccd1 _09362_/A
+ sky130_fd_sc_hd__and4_1
X_06573_ _08399_/A _06573_/B vssd1 vssd1 vccd1 vccd1 _06576_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09292_ _09507_/B _09293_/A vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__nand2_1
X_08312_ _08312_/A _08312_/B _08521_/B vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_59_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05524_ _06037_/A vssd1 vssd1 vccd1 vccd1 _05528_/A sky130_fd_sc_hd__inv_2
X_08243_ _08243_/A vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__inv_2
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05455_ _05732_/A _05617_/A _05456_/B vssd1 vssd1 vccd1 vccd1 _05493_/A sky130_fd_sc_hd__nand3_1
X_08174_ _08174_/A _08175_/A vssd1 vssd1 vccd1 vccd1 _08177_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05386_ _08780_/B _07216_/B vssd1 vssd1 vccd1 vccd1 _05830_/B sky130_fd_sc_hd__nand2_1
X_07125_ _07625_/A _07623_/A vssd1 vssd1 vccd1 vccd1 _07125_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07955__A _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _07198_/C vssd1 vssd1 vccd1 vccd1 _07195_/C sky130_fd_sc_hd__inv_2
XFILLER_0_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06007_ _06007_/A _06007_/B vssd1 vssd1 vccd1 vccd1 _06451_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07958_ _07958_/A vssd1 vssd1 vccd1 vccd1 _07971_/B sky130_fd_sc_hd__inv_2
XFILLER_0_97_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06909_ _07080_/B _07063_/A vssd1 vssd1 vccd1 vccd1 _06910_/B sky130_fd_sc_hd__nand2_1
X_07889_ _07889_/A _07889_/B vssd1 vssd1 vccd1 vccd1 _08048_/B sky130_fd_sc_hd__nand2_1
X_09628_ input54/X _10126_/B vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _09568_/A _09568_/C vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10403_ _10403_/A _10405_/A vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__and2_1
X_10334_ hold111/X _10339_/A vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__and2_1
XANTENNA__07584__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10263_/Y hold32/X vssd1 vssd1 vccd1 vccd1 _10299_/B sky130_fd_sc_hd__and2b_1
X_10196_ _10483_/Q hold94/X vssd1 vssd1 vccd1 vccd1 _10196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05832__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10443__A1 _10437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05240_ input60/X vssd1 vssd1 vccd1 vccd1 _07960_/B sky130_fd_sc_hd__buf_6
Xinput21 a_i[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput10 a_i[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput54 b_i[29] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_2
Xinput43 b_i[19] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput32 a_i[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput65 nrst vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
X_08930_ _08930_/A _08930_/B _09277_/A vssd1 vssd1 vccd1 vccd1 _09306_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07494__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08861_ input49/X vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__inv_2
X_07812_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _07925_/B sky130_fd_sc_hd__nand2_1
X_08792_ _09014_/A vssd1 vssd1 vccd1 vccd1 _08793_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ _07743_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__nand2_1
X_07674_ _07695_/B _07697_/A _07674_/C vssd1 vssd1 vccd1 vccd1 _07675_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09413_ _09416_/B _09658_/A vssd1 vssd1 vccd1 vccd1 _09415_/A sky130_fd_sc_hd__nand2_1
X_06625_ _06635_/A _06635_/B _06634_/B vssd1 vssd1 vccd1 vccd1 _06632_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09344_ _09347_/B _09520_/A vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06556_ _06146_/C _06146_/B _06146_/A vssd1 vssd1 vccd1 vccd1 _06570_/A sky130_fd_sc_hd__a21boi_2
X_09275_ _09274_/B _09275_/B _09473_/B vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__nand3b_1
X_06487_ _09962_/A _10052_/A vssd1 vssd1 vccd1 vccd1 _06490_/A sky130_fd_sc_hd__nand2_1
X_05507_ _09988_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _05998_/A sky130_fd_sc_hd__nand2_1
X_08226_ _08228_/B vssd1 vssd1 vccd1 vccd1 _08227_/B sky130_fd_sc_hd__inv_2
X_05438_ _05678_/A vssd1 vssd1 vccd1 vccd1 _05441_/A sky130_fd_sc_hd__inv_2
X_08157_ _08157_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _10383_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05369_ _05369_/A _05369_/B vssd1 vssd1 vccd1 vccd1 _05371_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ _07110_/A _07111_/A vssd1 vssd1 vccd1 vccd1 _07109_/A sky130_fd_sc_hd__nand2_1
X_08088_ _08088_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07039_ _07179_/C vssd1 vssd1 vccd1 vccd1 _07181_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _10050_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08963__B _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09497__D _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10317_ _10305_/A _10305_/B _10312_/A hold119/X vssd1 vssd1 vccd1 vccd1 _10319_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ hold24/X vssd1 vssd1 vccd1 vccd1 _10249_/B sky130_fd_sc_hd__inv_2
XFILLER_0_28_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10179_ hold85/A vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__inv_2
XFILLER_0_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09034__B _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06410_ _06413_/A vssd1 vssd1 vccd1 vccd1 _06411_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09806__B1 _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__B2 _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07390_ _07624_/B _07390_/B _07390_/C vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__nand3_2
XANTENNA__06674__A _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06341_ _06341_/A _06341_/B _06341_/C vssd1 vssd1 vccd1 vccd1 _06750_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _09060_/A _09060_/B _09060_/C vssd1 vssd1 vccd1 vccd1 _09061_/B sky130_fd_sc_hd__nand3_1
X_06272_ _06264_/A _06263_/A _06791_/B vssd1 vssd1 vccd1 vccd1 _06380_/B sky130_fd_sc_hd__o21ai_2
X_08011_ _08096_/A _08095_/B _08010_/Y vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__a21oi_1
X_05223_ _05344_/B _05343_/A vssd1 vssd1 vccd1 vccd1 _05347_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ _09962_/A _09962_/B vssd1 vssd1 vccd1 vccd1 _09964_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09209__B _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08913_ _08913_/A _08913_/B vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09888__A3 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _09894_/B _09894_/A vssd1 vssd1 vccd1 vccd1 _10117_/A sky130_fd_sc_hd__or2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08844_ _08847_/B _08847_/C vssd1 vssd1 vccd1 vccd1 _08846_/A sky130_fd_sc_hd__nand2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _08775_/A _08900_/A vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__nand2_1
X_05987_ input15/X vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__buf_4
XFILLER_0_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07726_ _07809_/A _07809_/B _07808_/B vssd1 vssd1 vccd1 vccd1 _07763_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07657_ _07659_/A vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__inv_2
XFILLER_0_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06608_ _08654_/B vssd1 vssd1 vccd1 vccd1 _08657_/C sky130_fd_sc_hd__inv_2
X_07588_ _07765_/B _07765_/A vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__or2_1
X_09327_ _09327_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__xor2_1
X_06539_ _06539_/A _06539_/B _06539_/C vssd1 vssd1 vccd1 vccd1 _06544_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09258_ _09256_/X _09258_/B vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08007__C _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09189_ _09189_/A _09190_/B _09189_/C vssd1 vssd1 vccd1 vccd1 _09190_/A sky130_fd_sc_hd__nand3_1
X_08209_ _10409_/A _08209_/B _10407_/A vssd1 vssd1 vccd1 vccd1 _08210_/C sky130_fd_sc_hd__and3_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05647__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10102_ _10101_/B _10102_/B _10102_/C vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__nand3b_1
X_10033_ _10036_/B _10036_/C vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07102__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08214__A _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07772__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05910_ _05927_/B _05928_/C _05928_/B vssd1 vssd1 vccd1 vccd1 _05912_/B sky130_fd_sc_hd__nand3_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06890_ _07018_/A _07013_/A vssd1 vssd1 vccd1 vccd1 _06890_/Y sky130_fd_sc_hd__nand2_1
X_05841_ _05852_/B _05852_/A vssd1 vssd1 vccd1 vccd1 _05924_/B sky130_fd_sc_hd__nand2_1
X_08560_ _08328_/A _08559_/Y _08329_/A vssd1 vssd1 vccd1 vccd1 _08563_/B sky130_fd_sc_hd__a21oi_1
X_05772_ _05772_/A vssd1 vssd1 vccd1 vccd1 _05773_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08491_ _08501_/B _08763_/B vssd1 vssd1 vccd1 vccd1 _08500_/A sky130_fd_sc_hd__nand2_1
X_07511_ _07510_/B _07511_/B _07511_/C vssd1 vssd1 vccd1 vccd1 _07512_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_71_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07442_ _07580_/C _07442_/B vssd1 vssd1 vccd1 vccd1 _07510_/B sky130_fd_sc_hd__nand2_1
X_07373_ _07373_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10505__RESET_B fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ _09110_/Y _08846_/B _09111_/Y vssd1 vssd1 vccd1 vccd1 _09115_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_57_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06324_ _06333_/B _06334_/C _06334_/B vssd1 vssd1 vccd1 vccd1 _06326_/B sky130_fd_sc_hd__nand3_1
X_09043_ _09357_/A _09043_/B vssd1 vssd1 vccd1 vccd1 _09046_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07947__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06255_ _06259_/A _06256_/A vssd1 vssd1 vccd1 vccd1 _06258_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05206_ input11/X vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__buf_4
X_06186_ _06186_/A _06186_/B vssd1 vssd1 vccd1 vccd1 _06187_/B sky130_fd_sc_hd__or2_1
XFILLER_0_96_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05467__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _10457_/B _10457_/A vssd1 vssd1 vccd1 vccd1 _10176_/A sky130_fd_sc_hd__nand2_1
X_09876_ _09876_/A _09876_/B _09876_/C vssd1 vssd1 vccd1 vccd1 _09885_/A sky130_fd_sc_hd__nand3_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08828_/B _08828_/A vssd1 vssd1 vccd1 vccd1 _08829_/A sky130_fd_sc_hd__or2_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05483__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ _08756_/Y _08465_/A _08757_/Y vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08689_ _08689_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _08691_/B sky130_fd_sc_hd__nand2_1
X_07709_ _07709_/A _07709_/B vssd1 vssd1 vccd1 vccd1 _07710_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06761__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08969__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08688__B _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _10016_/A _10016_/B _10016_/C vssd1 vssd1 vccd1 vccd1 _10018_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06040_ _06505_/B _06040_/B vssd1 vssd1 vccd1 vccd1 _06045_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07991_ _08337_/B vssd1 vssd1 vccd1 vccd1 _09890_/D sky130_fd_sc_hd__inv_2
XFILLER_0_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09730_ _09730_/A _09730_/B vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06942_ _06943_/B _06943_/A vssd1 vssd1 vccd1 vccd1 _06942_/Y sky130_fd_sc_hd__nand2_1
X_09661_ _09661_/A _09661_/B _09683_/A vssd1 vssd1 vccd1 vccd1 _09682_/B sky130_fd_sc_hd__nand3_1
X_06873_ _07033_/C _07033_/B _06872_/Y vssd1 vssd1 vccd1 vccd1 _07024_/A sky130_fd_sc_hd__a21oi_2
X_09592_ _09683_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09654_/A sky130_fd_sc_hd__nand2_1
X_08612_ _08614_/B _08614_/A vssd1 vssd1 vccd1 vccd1 _08882_/B sky130_fd_sc_hd__nor2_1
X_05824_ _06277_/B _05824_/B vssd1 vssd1 vccd1 vccd1 _05898_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05755_ _08814_/B vssd1 vssd1 vccd1 vccd1 _09560_/B sky130_fd_sc_hd__clkbuf_8
X_08543_ _08543_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08543_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08474_ _08476_/A vssd1 vssd1 vccd1 vccd1 _08475_/B sky130_fd_sc_hd__inv_2
X_05686_ _05686_/A _06126_/A _06107_/A vssd1 vssd1 vccd1 vccd1 _05688_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_45_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07425_ _08814_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _07430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07356_ _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07357_/A sky130_fd_sc_hd__nand2_1
X_07287_ _07467_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _07287_/Y sky130_fd_sc_hd__nor2_1
X_06307_ _09199_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _06656_/C sky130_fd_sc_hd__nand2_1
X_09026_ _09026_/A _09026_/B vssd1 vssd1 vccd1 vccd1 _09031_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06238_ _06661_/A _06660_/A vssd1 vssd1 vccd1 vccd1 _06243_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06169_ _06169_/A _06169_/B vssd1 vssd1 vccd1 vccd1 _06169_/Y sky130_fd_sc_hd__nor2_1
X_09928_ _09928_/A vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__inv_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09859_ _09860_/B _09860_/A vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__or2_1
XFILLER_0_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08971__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10496_ _10511_/CLK _10496_/D fanout100/X vssd1 vssd1 vccd1 vccd1 _10496_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05835__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 a_i[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09323__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05540_ _05540_/A _05540_/B _05540_/C vssd1 vssd1 vccd1 vccd1 _05572_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05471_ _05866_/A _05867_/A vssd1 vssd1 vccd1 vccd1 _05471_/Y sky130_fd_sc_hd__nor2_1
X_08190_ _08163_/A _08164_/B _08189_/A vssd1 vssd1 vccd1 vccd1 _10384_/B sky130_fd_sc_hd__a21o_1
X_07210_ _07169_/C _07169_/B _07165_/Y vssd1 vssd1 vccd1 vccd1 _07359_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07141_ _07680_/C vssd1 vssd1 vccd1 vccd1 _07679_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09630__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__B2 _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07072_ _07205_/A _07206_/A vssd1 vssd1 vccd1 vccd1 _07077_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08105__C _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06023_ _06406_/B _06023_/B vssd1 vssd1 vccd1 vccd1 _06049_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07974_ _07974_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07975_/B sky130_fd_sc_hd__nand2_1
X_09713_ _09714_/B _09714_/A vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__or2_1
X_06925_ _06929_/B _06926_/A vssd1 vssd1 vccd1 vccd1 _06928_/A sky130_fd_sc_hd__nand2_1
X_09644_ _09931_/B _09644_/B vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07960__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06856_ _06856_/A _06856_/B vssd1 vssd1 vccd1 vccd1 _07013_/B sky130_fd_sc_hd__nand2_1
X_05807_ _06299_/A _06299_/B vssd1 vssd1 vccd1 vccd1 _06214_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ _09575_/A _09575_/B vssd1 vssd1 vccd1 vccd1 _09575_/Y sky130_fd_sc_hd__nor2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ _06850_/C vssd1 vssd1 vccd1 vccd1 _06849_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08526_ _08527_/A _08527_/B vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05738_ input12/X vssd1 vssd1 vccd1 vccd1 _08862_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__09887__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08457_ _08719_/B _08458_/C _08458_/B vssd1 vssd1 vccd1 vccd1 _08463_/A sky130_fd_sc_hd__a21o_1
X_05669_ input39/X _08814_/B vssd1 vssd1 vccd1 vccd1 _05672_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10458__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07408_ _07411_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__nand2_1
X_08388_ _08388_/A _08388_/B vssd1 vssd1 vccd1 vccd1 _08390_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07339_ _07339_/A _07339_/B _07339_/C vssd1 vssd1 vccd1 vccd1 _07340_/B sky130_fd_sc_hd__nand3_1
X_10350_ _10376_/B hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__nor2_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09009_ _09011_/B _09010_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__nand3b_1
X_10281_ _10494_/Q hold27/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10479_ _10509_/CLK _10479_/D fanout100/X vssd1 vssd1 vccd1 vccd1 _10479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06710_ _06710_/A _06710_/B vssd1 vssd1 vccd1 vccd1 _06949_/B sky130_fd_sc_hd__nand2_1
X_07690_ _07690_/A _07690_/B _07690_/C vssd1 vssd1 vccd1 vccd1 _07693_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06677__A _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ _06641_/A _06641_/B vssd1 vssd1 vccd1 vccd1 _06644_/A sky130_fd_sc_hd__nand2_1
X_09360_ _09360_/A vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__inv_2
X_06572_ _06572_/A _06572_/B _06572_/C vssd1 vssd1 vccd1 vccd1 _06573_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09988__A _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09291_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08311_ _08314_/A _08313_/B _08314_/C vssd1 vssd1 vccd1 vccd1 _08521_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_47_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05523_ _09960_/B _09981_/B vssd1 vssd1 vccd1 vccd1 _06037_/A sky130_fd_sc_hd__nand2_1
X_08242_ _08244_/B _08244_/A vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__nor2_1
X_05454_ _05454_/A _05454_/B _05454_/C vssd1 vssd1 vccd1 vccd1 _05456_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08173_ _08176_/B _08176_/C vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05385_ input2/X vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__buf_6
X_07124_ _07390_/C _07390_/B _07123_/Y vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07955__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ _07055_/A _07055_/B vssd1 vssd1 vccd1 vccd1 _07198_/C sky130_fd_sc_hd__nand2_1
X_06006_ _06008_/B vssd1 vssd1 vccd1 vccd1 _06007_/B sky130_fd_sc_hd__inv_2
XANTENNA__05756__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07957_ _07959_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07958_/A sky130_fd_sc_hd__nor2_1
X_06908_ _07064_/B _07063_/A _07063_/B vssd1 vssd1 vccd1 vccd1 _07080_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_97_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07888_ _07890_/B _07890_/C vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__nand2_1
X_09627_ _09638_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09637_/A sky130_fd_sc_hd__nand2_1
X_06839_ _06839_/A _06839_/B _06839_/C vssd1 vssd1 vccd1 vccd1 _07138_/C sky130_fd_sc_hd__nand3_1
X_09558_ _09716_/A _09851_/A _09558_/C vssd1 vssd1 vccd1 vccd1 _09568_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08509_ _08513_/B _08513_/C vssd1 vssd1 vccd1 vccd1 _08512_/A sky130_fd_sc_hd__nand2_1
X_09489_ _09951_/A _09962_/B vssd1 vssd1 vccd1 vccd1 _09492_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ _10402_/A _10402_/B vssd1 vssd1 vccd1 vccd1 _10405_/A sky130_fd_sc_hd__nand2_1
X_10333_ hold110/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10339_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10264_ _10492_/Q hold31/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__nand2_1
X_10195_ hold88/X vssd1 vssd1 vccd1 vccd1 _10482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09530__B1 _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08217__A _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput22 a_i[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
Xinput11 a_i[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput55 b_i[2] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_4
Xinput44 b_i[1] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_4
Xinput33 b_i[0] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08860_ _08575_/A _08575_/C _08575_/B vssd1 vssd1 vccd1 vccd1 _08879_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_20_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07811_ _07812_/B _07812_/A vssd1 vssd1 vccd1 vccd1 _07811_/Y sky130_fd_sc_hd__nor2_1
X_08791_ _08789_/Y _08498_/B _08790_/Y vssd1 vssd1 vccd1 vccd1 _09014_/A sky130_fd_sc_hd__a21oi_2
X_07742_ _07824_/B _07826_/B _07741_/Y vssd1 vssd1 vccd1 vccd1 _07743_/B sky130_fd_sc_hd__a21oi_1
X_07673_ _07697_/B _07673_/B vssd1 vssd1 vccd1 vccd1 _07675_/A sky130_fd_sc_hd__nand2_1
X_09412_ _09412_/A _09412_/B _09658_/B vssd1 vssd1 vccd1 vccd1 _09658_/A sky130_fd_sc_hd__nand3_2
X_06624_ _06634_/A _06635_/C vssd1 vssd1 vccd1 vccd1 _06632_/B sky130_fd_sc_hd__nand2_1
X_09343_ _09343_/A _09343_/B _09520_/B vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06555_ _06555_/A _08322_/A vssd1 vssd1 vccd1 vccd1 _06571_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _09274_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09276_/A sky130_fd_sc_hd__nand2_1
X_06486_ _06500_/A _06501_/C vssd1 vssd1 vccd1 vccd1 _06499_/A sky130_fd_sc_hd__nand2_1
X_05506_ input14/X vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__buf_4
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08225_ _08225_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08228_/B sky130_fd_sc_hd__nand2_1
X_05437_ input37/X _08810_/B vssd1 vssd1 vccd1 vccd1 _05678_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08156_ _08112_/Y _08158_/C vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_43_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05368_ _05370_/C vssd1 vssd1 vccd1 vccd1 _05369_/B sky130_fd_sc_hd__inv_2
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06870__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _07110_/B vssd1 vssd1 vccd1 vccd1 _07111_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05299_ input61/X vssd1 vssd1 vccd1 vccd1 _08248_/B sky130_fd_sc_hd__clkbuf_8
X_08087_ _08087_/A _08087_/B vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07038_ _10052_/A _08214_/A vssd1 vssd1 vccd1 vccd1 _07179_/C sky130_fd_sc_hd__nand2_1
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06764__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10316_ hold10/X _10308_/Y hold118/X vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ hold99/A hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__nand2_1
X_10178_ _10480_/Q hold43/X vssd1 vssd1 vccd1 vccd1 _10381_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09806__A1 _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__B2 _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__A2 _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06674__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06340_ _06342_/B _06340_/B vssd1 vssd1 vccd1 vccd1 _06341_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06271_ _06271_/A _06271_/B vssd1 vssd1 vccd1 vccd1 _06791_/B sky130_fd_sc_hd__nand2_1
X_08010_ _08010_/A _08010_/B vssd1 vssd1 vccd1 vccd1 _08010_/Y sky130_fd_sc_hd__nor2_1
X_05222_ _09962_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _05343_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _09961_/A vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__inv_2
XFILLER_0_12_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08912_ _08914_/B vssd1 vssd1 vccd1 vccd1 _08913_/B sky130_fd_sc_hd__inv_2
X_09892_ _10117_/B _09892_/B vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__nand2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _09111_/A _09056_/A _08843_/C vssd1 vssd1 vccd1 vccd1 _08847_/C sky130_fd_sc_hd__nand3_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ _08774_/A _08900_/A _08775_/A vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__nand3_2
X_05986_ _06432_/A vssd1 vssd1 vccd1 vccd1 _05990_/A sky130_fd_sc_hd__inv_2
X_07725_ _07725_/A _07725_/B vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07656_ _07654_/Y _07640_/C _07655_/Y vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06607_ _06609_/B _06609_/A vssd1 vssd1 vccd1 vccd1 _08654_/B sky130_fd_sc_hd__nor2_2
X_07587_ _07589_/B _07587_/B vssd1 vssd1 vccd1 vccd1 _07765_/A sky130_fd_sc_hd__nand2_1
X_09326_ _09324_/X _09326_/B vssd1 vssd1 vccd1 vccd1 _09327_/B sky130_fd_sc_hd__and2b_1
X_06538_ _06538_/A vssd1 vssd1 vccd1 vccd1 _06539_/C sky130_fd_sc_hd__inv_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09257_ _09988_/A input21/X _09987_/A input20/X vssd1 vssd1 vccd1 vccd1 _09258_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08481__B1 _08479_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06469_ _06469_/A _06469_/B _06469_/C vssd1 vssd1 vccd1 vccd1 _06518_/C sky130_fd_sc_hd__nand3_1
X_08208_ _08208_/A vssd1 vssd1 vccd1 vccd1 _10407_/A sky130_fd_sc_hd__inv_2
X_09188_ _09188_/A _09188_/B vssd1 vssd1 vccd1 vccd1 _09189_/C sky130_fd_sc_hd__nor2_1
XANTENNA__08007__D _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08139_ _10126_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__nand2_1
X_10101_ _10101_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__nand2_1
X_10032_ _10032_/A _10032_/B vssd1 vssd1 vccd1 vccd1 _10036_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_98_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08214__B _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08230__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05840_ _05918_/B _05918_/C _05919_/B vssd1 vssd1 vccd1 vccd1 _05852_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _07510_/A _07510_/B vssd1 vssd1 vccd1 vccd1 _07512_/A sky130_fd_sc_hd__nand2_1
X_05771_ _05766_/B _05765_/B _05809_/B vssd1 vssd1 vccd1 vccd1 _05814_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08490_ _08490_/A _08490_/B _08737_/A vssd1 vssd1 vccd1 vccd1 _08763_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06685__A _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07441_ _07442_/B _07441_/B _07441_/C vssd1 vssd1 vccd1 vccd1 _07580_/C sky130_fd_sc_hd__nand3_1
XANTENNA__10000__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ _07374_/C vssd1 vssd1 vccd1 vccd1 _07373_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _09111_/A _09111_/B vssd1 vssd1 vccd1 vccd1 _09111_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06323_ _06334_/A vssd1 vssd1 vccd1 vccd1 _06333_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10491__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ _09042_/A _09042_/B _09042_/C vssd1 vssd1 vccd1 vccd1 _09043_/B sky130_fd_sc_hd__nand3_1
X_06254_ _06257_/B vssd1 vssd1 vccd1 vccd1 _06259_/A sky130_fd_sc_hd__inv_2
X_06185_ _06185_/A _06185_/B vssd1 vssd1 vccd1 vccd1 _06190_/B sky130_fd_sc_hd__and2_1
XFILLER_0_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05205_ _05251_/A vssd1 vssd1 vccd1 vccd1 _05216_/A sky130_fd_sc_hd__inv_2
XFILLER_0_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09944_ _09944_/A vssd1 vssd1 vccd1 vccd1 _10457_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09875_ _09879_/B _09878_/A vssd1 vssd1 vccd1 vccd1 _09876_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08140__A _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05764__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08826_ _09083_/C _08826_/B vssd1 vssd1 vccd1 vccd1 _08828_/A sky130_fd_sc_hd__xor2_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05483__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ _08757_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _08757_/Y sky130_fd_sc_hd__nor2_1
X_05969_ _05969_/A _05969_/B vssd1 vssd1 vccd1 vccd1 _05969_/Y sky130_fd_sc_hd__nor2_1
X_08688_ _08688_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _08691_/A sky130_fd_sc_hd__nand2_1
X_07708_ _07708_/A _10428_/A vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__nand2_1
X_07639_ _07639_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _07647_/B sky130_fd_sc_hd__nand2_1
X_09309_ _09343_/B _09520_/B vssd1 vssd1 vccd1 vccd1 _09341_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05939__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__B1 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08969__B _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05674__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07990_ _07990_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _08020_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06941_ _06934_/A _06933_/A _07093_/A vssd1 vssd1 vccd1 vccd1 _06952_/B sky130_fd_sc_hd__o21ai_1
X_09660_ _09660_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09667_/B sky130_fd_sc_hd__nand2_1
X_08611_ _08342_/A _08341_/B _08341_/A vssd1 vssd1 vccd1 vccd1 _08614_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06872_ _07030_/B _07029_/A vssd1 vssd1 vccd1 vccd1 _06872_/Y sky130_fd_sc_hd__nor2_1
X_09591_ _09591_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09656_/C sky130_fd_sc_hd__nand2_1
X_05823_ _05824_/B _05823_/B _05823_/C vssd1 vssd1 vccd1 vccd1 _06277_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_89_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08542_ _08543_/B _08543_/A vssd1 vssd1 vccd1 vccd1 _08542_/Y sky130_fd_sc_hd__nand2_1
X_05754_ input37/X _08825_/B vssd1 vssd1 vccd1 vccd1 _05760_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08473_ _08266_/B _08266_/C _08243_/A vssd1 vssd1 vccd1 vccd1 _08476_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05685_ _06107_/B _05685_/B vssd1 vssd1 vccd1 vccd1 _05688_/A sky130_fd_sc_hd__nand2_1
X_07424_ _07508_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07507_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07355_ _07374_/A _07374_/B vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ _07471_/C vssd1 vssd1 vccd1 vccd1 _07470_/B sky130_fd_sc_hd__inv_2
X_06306_ _06656_/A _06656_/B vssd1 vssd1 vccd1 vccd1 _06309_/A sky130_fd_sc_hd__nand2_1
X_09025_ _09026_/B _09026_/A vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06237_ _06661_/B vssd1 vssd1 vccd1 vccd1 _06660_/A sky130_fd_sc_hd__inv_2
XFILLER_0_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06168_ _06169_/B _06169_/A vssd1 vssd1 vccd1 vccd1 _06168_/Y sky130_fd_sc_hd__nand2_1
X_06099_ _06594_/B _06099_/B vssd1 vssd1 vccd1 vccd1 _06101_/A sky130_fd_sc_hd__nand2_1
X_09927_ _09929_/B _09929_/A vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__nor2_1
X_09858_ _10091_/B _09858_/B vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__nand2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09789_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09790_/A sky130_fd_sc_hd__nand2_1
X_08809_ _08809_/A vssd1 vssd1 vccd1 vccd1 _08820_/B sky130_fd_sc_hd__inv_2
XANTENNA__07214__A _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_3__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05669__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10495_ _10495_/CLK hold30/X fanout99/X vssd1 vssd1 vccd1 vccd1 _10495_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 a_i[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09323__B _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05470_ _05870_/B vssd1 vssd1 vccd1 vccd1 _05871_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ _07679_/A _07680_/C vssd1 vssd1 vccd1 vccd1 _07143_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09630__A2 _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07071_ _07205_/B vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__inv_2
XANTENNA__08105__D _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06022_ _06022_/A _06022_/B vssd1 vssd1 vccd1 vccd1 _06023_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09712_ _10048_/B _09712_/B vssd1 vssd1 vccd1 vccd1 _09714_/A sky130_fd_sc_hd__nand2_1
X_07973_ _08036_/B vssd1 vssd1 vccd1 vccd1 _08038_/B sky130_fd_sc_hd__inv_2
X_06924_ _06927_/B vssd1 vssd1 vccd1 vccd1 _06929_/B sky130_fd_sc_hd__inv_2
X_09643_ _09931_/A vssd1 vssd1 vccd1 vccd1 _09644_/B sky130_fd_sc_hd__inv_2
X_06855_ _06857_/A _06857_/B vssd1 vssd1 vccd1 vccd1 _06856_/A sky130_fd_sc_hd__nand2_1
X_09574_ _09575_/B _09575_/A vssd1 vssd1 vccd1 vccd1 _09574_/Y sky130_fd_sc_hd__nand2_1
X_05806_ _06280_/B _06299_/B _06279_/B vssd1 vssd1 vccd1 vccd1 _06299_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _09528_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08527_/B sky130_fd_sc_hd__nand2_1
X_06786_ _06786_/A _06786_/B vssd1 vssd1 vccd1 vccd1 _06850_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05737_ _05781_/A _05781_/B vssd1 vssd1 vccd1 vccd1 _05780_/A sky130_fd_sc_hd__nand2_1
X_08456_ _08456_/A vssd1 vssd1 vccd1 vccd1 _08458_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05668_ _05672_/A vssd1 vssd1 vccd1 vccd1 _05671_/A sky130_fd_sc_hd__inv_2
XFILLER_0_92_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08387_ _08391_/A _08391_/C vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__nand2_1
X_07407_ _07643_/A _07407_/B _07407_/C vssd1 vssd1 vccd1 vccd1 _07411_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05599_ _05599_/A _05599_/B vssd1 vssd1 vccd1 vccd1 _05605_/A sky130_fd_sc_hd__nand2_1
X_07338_ _07338_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07378_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07269_ _07269_/A vssd1 vssd1 vccd1 vccd1 _07423_/B sky130_fd_sc_hd__inv_2
X_09008_ _09008_/A _09233_/A _09008_/C vssd1 vssd1 vccd1 vccd1 _09217_/B sky130_fd_sc_hd__nand3_1
X_10280_ _10494_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_20_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10478_ _10511_/CLK _10478_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__05862__A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06677__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ _06640_/A _06640_/B vssd1 vssd1 vccd1 vccd1 _10435_/A sky130_fd_sc_hd__nand2_1
X_06571_ _06571_/A _06570_/A vssd1 vssd1 vccd1 vccd1 _06572_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09290_ _09290_/A vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__inv_2
X_08310_ _08315_/B vssd1 vssd1 vccd1 vccd1 _08312_/B sky130_fd_sc_hd__inv_2
X_05522_ _08688_/A vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__buf_8
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08241_ _08241_/A _08449_/C vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__nand2_1
X_05453_ _05453_/A _05453_/B _05453_/C vssd1 vssd1 vccd1 vccd1 _05454_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08172_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08176_/B sky130_fd_sc_hd__nand2_1
X_05384_ _05396_/B _05397_/C _05397_/A vssd1 vssd1 vccd1 vccd1 _05395_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ _07392_/A _07391_/A vssd1 vssd1 vccd1 vccd1 _07123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07054_ _07054_/A _07054_/B _07054_/C vssd1 vssd1 vccd1 vccd1 _07055_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06005_ _09963_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _06008_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05756__B _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07956_ _09361_/D _08689_/A vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06868__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ _06907_/A _06907_/B vssd1 vssd1 vccd1 vccd1 _07063_/B sky130_fd_sc_hd__nand2_1
X_07887_ _07887_/A _07887_/B _07887_/C vssd1 vssd1 vccd1 vccd1 _07890_/C sky130_fd_sc_hd__nand3_1
X_09626_ _09626_/A _09626_/B _09916_/A vssd1 vssd1 vccd1 vccd1 _09638_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06838_ _06838_/A _06838_/B vssd1 vssd1 vccd1 vccd1 _07138_/B sky130_fd_sc_hd__nand2_1
X_09557_ _09557_/A vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__inv_2
X_06769_ _06769_/A vssd1 vssd1 vccd1 vccd1 _06771_/A sky130_fd_sc_hd__inv_2
XFILLER_0_93_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ _09811_/B _09488_/B vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08508_ _08508_/A _08763_/A _08839_/A vssd1 vssd1 vccd1 vccd1 _08513_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08439_ _08439_/A vssd1 vssd1 vccd1 vccd1 _08441_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _10402_/B _10402_/A vssd1 vssd1 vccd1 vccd1 _10403_/A sky130_fd_sc_hd__or2_1
XFILLER_0_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ _10333_/B hold110/X vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08323__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _10492_/Q hold31/X vssd1 vssd1 vccd1 vccd1 _10263_/Y sky130_fd_sc_hd__nor2_1
X_10194_ hold87/X _10199_/A vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__and2_1
XANTENNA__09530__A1 _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__B2 _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__B _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08217__B input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 a_i[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
Xinput45 b_i[20] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
Xinput34 b_i[10] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput23 a_i[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput56 b_i[30] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05857__A _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__A _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08790_ _09227_/A _10044_/B _08790_/C vssd1 vssd1 vccd1 vccd1 _08790_/Y sky130_fd_sc_hd__nor3_1
X_07810_ _07810_/A _07810_/B vssd1 vssd1 vccd1 vccd1 _07812_/A sky130_fd_sc_hd__nand2_1
X_07741_ _07741_/A _07741_/B vssd1 vssd1 vccd1 vccd1 _07741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09999__A _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ _07697_/A vssd1 vssd1 vccd1 vccd1 _07673_/B sky130_fd_sc_hd__inv_2
X_09411_ _09411_/A vssd1 vssd1 vccd1 vccd1 _09412_/A sky130_fd_sc_hd__inv_2
X_06623_ _06635_/A _06635_/B vssd1 vssd1 vccd1 vccd1 _06634_/A sky130_fd_sc_hd__nand2_1
X_09342_ _09342_/A vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__inv_2
X_06554_ _06553_/B _08322_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05505_ _05983_/A vssd1 vssd1 vccd1 vccd1 _05538_/B sky130_fd_sc_hd__inv_2
X_09273_ _09434_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06485_ _06077_/B _06076_/B _06484_/Y vssd1 vssd1 vccd1 vccd1 _06501_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08224_ _08228_/A _08228_/C vssd1 vssd1 vccd1 vccd1 _08227_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05436_ input30/X vssd1 vssd1 vccd1 vccd1 _08810_/B sky130_fd_sc_hd__clkbuf_8
X_08155_ _08180_/B _08180_/A vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05367_ _09684_/B _07960_/B vssd1 vssd1 vccd1 vccd1 _05370_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06870__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ _07111_/B vssd1 vssd1 vccd1 vccd1 _07110_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05298_ _05303_/A vssd1 vssd1 vccd1 vccd1 _05302_/A sky130_fd_sc_hd__inv_2
X_08086_ _08086_/A _08086_/B vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__nor2_1
X_07037_ _07178_/B _07177_/A vssd1 vssd1 vccd1 vccd1 _07181_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08988_ _08740_/A _08738_/A _08761_/A vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__o21ai_1
X_07939_ _07939_/A vssd1 vssd1 vccd1 vccd1 _07940_/B sky130_fd_sc_hd__inv_2
XFILLER_0_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _09609_/A vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__inv_2
XFILLER_0_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10315_ _10313_/Y hold14/X vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ hold99/X hold23/X vssd1 vssd1 vccd1 vccd1 _10249_/A sky130_fd_sc_hd__nor2_1
X_10177_ _10177_/A _10177_/B vssd1 vssd1 vccd1 vccd1 _10479_/D sky130_fd_sc_hd__nand2_1
XANTENNA__09806__A2 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06270_ _06658_/C vssd1 vssd1 vccd1 vccd1 _06271_/B sky130_fd_sc_hd__inv_2
XANTENNA__06971__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05221_ _09960_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _05344_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09960_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08911_ _08911_/A _08911_/B vssd1 vssd1 vccd1 vccd1 _08914_/B sky130_fd_sc_hd__nand2_1
X_09891_ input52/X _09601_/B input53/X _10112_/B vssd1 vssd1 vccd1 vccd1 _09892_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08842_ _09111_/B _08842_/B vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__nand2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08773_ _08773_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08775_/A sky130_fd_sc_hd__nand2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05985_ _08420_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _06432_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07307__A _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07724_ _07728_/B vssd1 vssd1 vccd1 vccd1 _07725_/A sky130_fd_sc_hd__inv_2
XFILLER_0_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07655_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07655_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06606_ _06172_/A _06173_/A _06180_/A vssd1 vssd1 vccd1 vccd1 _06609_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07586_ _07586_/A _07586_/B vssd1 vssd1 vccd1 vccd1 _07587_/B sky130_fd_sc_hd__nand2_1
X_09325_ _09963_/A _09816_/B _09962_/A _09496_/B vssd1 vssd1 vccd1 vccd1 _09326_/B
+ sky130_fd_sc_hd__a22o_1
X_06537_ _06537_/A _08361_/A _06537_/C vssd1 vssd1 vccd1 vccd1 _06539_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09256_ _09988_/A _09987_/A input20/X input21/X vssd1 vssd1 vccd1 vccd1 _09256_/X
+ sky130_fd_sc_hd__and4_1
X_06468_ _06468_/A _06468_/B vssd1 vssd1 vccd1 vccd1 _06469_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__nand2_1
X_05419_ _05419_/A vssd1 vssd1 vccd1 vccd1 _05420_/B sky130_fd_sc_hd__inv_2
X_09187_ _10437_/A _09187_/B vssd1 vssd1 vccd1 vccd1 _09196_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06399_ _06399_/A _06399_/B vssd1 vssd1 vccd1 vccd1 _06399_/Y sky130_fd_sc_hd__nor2_1
X_08138_ _08138_/A _08138_/B vssd1 vssd1 vccd1 vccd1 _08180_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08069_ _08069_/A _08072_/B _08069_/C vssd1 vssd1 vccd1 vccd1 _08083_/B sky130_fd_sc_hd__nand3_1
X_10100_ _10100_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__nand2_1
X_10031_ _10032_/B _10032_/A vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__or2_1
XFILLER_0_11_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08230__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10229_ _10229_/A hold36/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__nand2_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_05770_ _05770_/A _05770_/B vssd1 vssd1 vccd1 vccd1 _05809_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07440_ _07440_/A _07440_/B vssd1 vssd1 vccd1 vccd1 _07441_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07371_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07374_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09110_ _09111_/B _09111_/A vssd1 vssd1 vccd1 vccd1 _09110_/Y sky130_fd_sc_hd__nand2_1
X_06322_ _06646_/B _06646_/C vssd1 vssd1 vccd1 vccd1 _06651_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09041_ _09041_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06253_ _06699_/C _06699_/B _06252_/Y vssd1 vssd1 vccd1 vccd1 _06264_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05204_ _09962_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _05251_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06184_ _06197_/B _06198_/B _06198_/C vssd1 vssd1 vccd1 vccd1 _06196_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_13_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09943_ _09943_/A _10176_/C vssd1 vssd1 vccd1 vccd1 _09944_/A sky130_fd_sc_hd__nand2_1
X_09874_ _09874_/A _09612_/A vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__or2b_1
XANTENNA__08140__B _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05764__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ input46/X _08825_/B vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__nand2_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _08757_/B _08757_/A vssd1 vssd1 vccd1 vccd1 _08756_/Y sky130_fd_sc_hd__nand2_1
X_05968_ _05969_/B _05969_/A vssd1 vssd1 vccd1 vccd1 _06211_/C sky130_fd_sc_hd__nand2_1
X_08687_ _08927_/B _08698_/C vssd1 vssd1 vccd1 vccd1 _08697_/A sky130_fd_sc_hd__nand2_1
X_07707_ _07707_/A _07707_/B vssd1 vssd1 vccd1 vccd1 _07708_/A sky130_fd_sc_hd__nand2_1
X_05899_ _05899_/A _05899_/B vssd1 vssd1 vccd1 vccd1 _05900_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07638_ _07640_/C vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__inv_2
XFILLER_0_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07569_ _07569_/A _07569_/B vssd1 vssd1 vccd1 vccd1 _07809_/B sky130_fd_sc_hd__nand2_2
X_09308_ _09307_/B _09308_/B _09479_/A vssd1 vssd1 vccd1 vccd1 _09520_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09239_ _09242_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _09240_/C sky130_fd_sc_hd__nand2_1
XANTENNA__05939__B _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06116__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09954__B2 _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__A1 _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05674__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _10016_/B _10016_/C vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10509__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06940_ _06940_/A _06940_/B vssd1 vssd1 vccd1 vccd1 _07093_/A sky130_fd_sc_hd__nand2_1
X_06871_ _07031_/C vssd1 vssd1 vccd1 vccd1 _07033_/B sky130_fd_sc_hd__inv_2
X_08610_ _08875_/B _08610_/B vssd1 vssd1 vccd1 vccd1 _08614_/B sky130_fd_sc_hd__nand2_1
X_05822_ _06216_/B _06213_/B vssd1 vssd1 vccd1 vccd1 _05823_/C sky130_fd_sc_hd__nand2_1
X_09590_ _09348_/A _09349_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_82_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09072__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ _08547_/A _08547_/C vssd1 vssd1 vccd1 vccd1 _08546_/A sky130_fd_sc_hd__nand2_1
X_05753_ _05773_/C _05773_/B vssd1 vssd1 vccd1 vccd1 _05762_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08472_ _08476_/B _08673_/A vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__nand2_1
X_05684_ _05684_/A _06133_/B _05687_/A vssd1 vssd1 vccd1 vccd1 _06133_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_9_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _07270_/Y _07423_/B _07423_/C vssd1 vssd1 vccd1 vccd1 _07508_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07354_ _07386_/B _07354_/B vssd1 vssd1 vccd1 vccd1 _07374_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07285_ _07285_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07471_/C sky130_fd_sc_hd__nand2_1
X_06305_ _06305_/A _06305_/B vssd1 vssd1 vccd1 vccd1 _06656_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ _09024_/A _09023_/X vssd1 vssd1 vccd1 vccd1 _09026_/A sky130_fd_sc_hd__nor2b_1
X_06236_ _10051_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _06661_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06167_ _06586_/A _06173_/C vssd1 vssd1 vccd1 vccd1 _06172_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06098_ _06404_/B _06098_/B _06098_/C vssd1 vssd1 vccd1 vccd1 _06404_/A sky130_fd_sc_hd__nand3_1
X_09926_ _09926_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09857_ input49/X _09560_/B input50/X _10083_/B vssd1 vssd1 vccd1 vccd1 _09858_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09788_ _09788_/A _09971_/A vssd1 vssd1 vccd1 vccd1 _09792_/C sky130_fd_sc_hd__nand2_1
X_08808_ _08557_/C _08557_/B _08551_/Y vssd1 vssd1 vccd1 vccd1 _08809_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_95_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08739_ _08739_/A vssd1 vssd1 vccd1 vccd1 _08740_/A sky130_fd_sc_hd__inv_2
XANTENNA__07214__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05669__B _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _10494_/CLK _10494_/D fanout99/X vssd1 vssd1 vccd1 vccd1 _10494_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08996__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10481__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07070_ _08810_/B _08248_/B vssd1 vssd1 vccd1 vccd1 _07205_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06021_ _06408_/A _06021_/B vssd1 vssd1 vccd1 vccd1 _06406_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05595__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09711_ _09199_/A _09533_/B _09548_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _09712_/B
+ sky130_fd_sc_hd__a22o_1
X_07972_ _07974_/B _07974_/A vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__nor2_1
X_06923_ _07109_/C _07109_/B _06922_/Y vssd1 vssd1 vccd1 vccd1 _06934_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09642_ _09640_/Y _09251_/B _09641_/Y vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__a21oi_2
X_06854_ _06854_/A _06854_/B _06854_/C vssd1 vssd1 vccd1 vccd1 _06857_/B sky130_fd_sc_hd__nand3_1
X_09573_ _09741_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__nand2_1
X_06785_ _06784_/B _06785_/B _06785_/C vssd1 vssd1 vccd1 vccd1 _06786_/B sky130_fd_sc_hd__nand3b_1
X_05805_ _05805_/A _05805_/B vssd1 vssd1 vccd1 vccd1 _06279_/B sky130_fd_sc_hd__nand2_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ input40/X _09022_/C vssd1 vssd1 vccd1 vccd1 _08527_/A sky130_fd_sc_hd__nand2_1
X_05736_ _06186_/A _06176_/A _05736_/C vssd1 vssd1 vccd1 vccd1 _05781_/B sky130_fd_sc_hd__nand3_1
X_08455_ _09960_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _08456_/A sky130_fd_sc_hd__nand2_1
X_05667_ input40/X _08825_/B vssd1 vssd1 vccd1 vccd1 _05672_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08386_ _08386_/A _08386_/B _08386_/C vssd1 vssd1 vccd1 vccd1 _08391_/C sky130_fd_sc_hd__nand3_1
X_05598_ _06121_/B vssd1 vssd1 vccd1 vccd1 _05599_/B sky130_fd_sc_hd__inv_2
X_07406_ _07406_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07411_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07337_ _07339_/C vssd1 vssd1 vccd1 vccd1 _07338_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ _09601_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _07269_/A sky130_fd_sc_hd__nand2_1
X_09007_ _09007_/A vssd1 vssd1 vccd1 vccd1 _09008_/C sky130_fd_sc_hd__inv_2
XFILLER_0_60_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07199_ _07346_/A _07199_/B vssd1 vssd1 vccd1 vccd1 _07228_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06219_ _06219_/A _06219_/B _06219_/C vssd1 vssd1 vccd1 vccd1 _06377_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_41_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09909_ _10141_/A _09914_/C vssd1 vssd1 vccd1 vccd1 _10156_/B sky130_fd_sc_hd__nand2_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10477_ _10509_/CLK _10477_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05862__B _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06570_ _06570_/A _06571_/A vssd1 vssd1 vccd1 vccd1 _06572_/A sky130_fd_sc_hd__or2b_1
XANTENNA__06974__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05521_ _05983_/B _05983_/A vssd1 vssd1 vccd1 vccd1 _05537_/B sky130_fd_sc_hd__nand2_1
X_08240_ _08240_/A _08240_/B _08449_/B vssd1 vssd1 vccd1 vccd1 _08449_/C sky130_fd_sc_hd__nand3_2
X_05452_ _05452_/A _05452_/B vssd1 vssd1 vccd1 vccd1 _05454_/A sky130_fd_sc_hd__nand2_1
X_08171_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08172_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07122_ _07393_/C vssd1 vssd1 vccd1 vccd1 _07390_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05383_ _05379_/Y _05369_/B _05380_/Y vssd1 vssd1 vccd1 vccd1 _05396_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07053_ _07060_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07054_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06004_ _06008_/A vssd1 vssd1 vccd1 vccd1 _06007_/A sky130_fd_sc_hd__inv_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07955_ _08337_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _07959_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06868__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ _06906_/A _06906_/B vssd1 vssd1 vccd1 vccd1 _07063_/A sky130_fd_sc_hd__nand2_1
X_09625_ _09916_/B _09625_/B vssd1 vssd1 vccd1 vccd1 _09638_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07045__A _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ _07886_/A _07886_/B vssd1 vssd1 vccd1 vccd1 _07890_/B sky130_fd_sc_hd__nand2_1
X_06837_ _06839_/A _06839_/B vssd1 vssd1 vccd1 vccd1 _06838_/A sky130_fd_sc_hd__nand2_1
X_09556_ _09851_/B _09557_/A vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__nand2_1
X_06768_ _06853_/A _06854_/A vssd1 vssd1 vccd1 vccd1 _06768_/Y sky130_fd_sc_hd__nand2_1
X_09487_ _09951_/B _09485_/C _09963_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _09488_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08507_ _08839_/B _08507_/B vssd1 vssd1 vccd1 vccd1 _08513_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05719_ _05719_/A _05719_/B vssd1 vssd1 vccd1 vccd1 _05720_/A sky130_fd_sc_hd__nand2_1
X_06699_ _06699_/A _06699_/B _06699_/C vssd1 vssd1 vccd1 vccd1 _06703_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08438_ _09951_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _08439_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08369_ _08370_/A _08371_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08378_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _10400_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _10319_/A _10319_/B _10326_/A hold109/X vssd1 vssd1 vccd1 vccd1 hold110/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08323__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ _10266_/B hold25/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__xor2_1
X_10193_ hold86/X _10193_/B vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09530__A2 _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__B1 _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05203__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 a_i[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
Xinput46 b_i[21] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_4
Xinput35 b_i[11] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 a_i[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput57 b_i[31] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05857__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07740_ _07740_/A vssd1 vssd1 vccd1 vccd1 _07826_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09999__B input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ _07695_/B _07674_/C vssd1 vssd1 vccd1 vccd1 _07697_/B sky130_fd_sc_hd__nand2_1
X_09410_ _09410_/A _09411_/A vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__nand2_1
X_06622_ _08655_/B _06622_/B vssd1 vssd1 vccd1 vccd1 _06635_/B sky130_fd_sc_hd__nand2_1
X_09341_ _09341_/A _09342_/A vssd1 vssd1 vccd1 vccd1 _09347_/B sky130_fd_sc_hd__nand2_1
X_06553_ _06553_/A _06553_/B vssd1 vssd1 vccd1 vccd1 _06555_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05504_ _05262_/C _05262_/B _05503_/Y vssd1 vssd1 vccd1 vccd1 _05983_/A sky130_fd_sc_hd__a21oi_2
X_09272_ _09270_/Y _09272_/B vssd1 vssd1 vccd1 vccd1 _09273_/B sky130_fd_sc_hd__and2b_1
X_06484_ _06484_/A _06484_/B vssd1 vssd1 vccd1 vccd1 _06484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08223_ _08223_/A _08223_/B vssd1 vssd1 vccd1 vccd1 _08228_/C sky130_fd_sc_hd__nand2_1
X_05435_ _05452_/B _05453_/C _05453_/A vssd1 vssd1 vccd1 vccd1 _05617_/B sky130_fd_sc_hd__nand3_1
X_08154_ _08184_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__and2_1
X_05366_ input5/X vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__buf_8
XFILLER_0_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07105_ _07292_/C _07292_/B _07104_/Y vssd1 vssd1 vccd1 vccd1 _07113_/A sky130_fd_sc_hd__a21o_1
X_08085_ _10394_/B _10398_/A vssd1 vssd1 vccd1 vccd1 _08086_/A sky130_fd_sc_hd__nand2_1
X_07036_ _09533_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _07177_/A sky130_fd_sc_hd__nand2_1
X_05297_ input5/X _08247_/B vssd1 vssd1 vccd1 vccd1 _05303_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09255__A _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _08990_/B _08990_/C vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__nand2_1
X_07938_ _07938_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07940_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_2__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10511_/CLK sky130_fd_sc_hd__clkbuf_16
X_07869_ _07925_/A _07925_/B vssd1 vssd1 vccd1 vccd1 _07924_/A sky130_fd_sc_hd__nand2_1
X_09608_ _09608_/A _09608_/B vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__nand2_1
X_09539_ _09703_/A _09702_/A vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08318__B _08319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08334__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10314_ _10498_/Q hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__nand2_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ _10250_/A hold41/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__xor2_1
X_10176_ _10176_/A _10176_/B _10176_/C vssd1 vssd1 vccd1 vccd1 _10177_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05220_ _05338_/B _05338_/C vssd1 vssd1 vccd1 vccd1 _05337_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06971__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09890_ _10113_/A _10113_/C _10113_/D _09890_/D vssd1 vssd1 vccd1 vccd1 _10117_/B
+ sky130_fd_sc_hd__or4_1
X_08910_ _08914_/A _09262_/A vssd1 vssd1 vccd1 vccd1 _08913_/A sky130_fd_sc_hd__nand2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08841_ _09111_/A vssd1 vssd1 vccd1 vccd1 _08842_/B sky130_fd_sc_hd__inv_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08900_/B _08772_/B vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__nand2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05984_ _05537_/B _05537_/C _05983_/Y vssd1 vssd1 vccd1 vccd1 _06406_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07307__B _09392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ _07887_/B _07887_/C vssd1 vssd1 vccd1 vccd1 _07886_/B sky130_fd_sc_hd__nand2_1
X_07654_ _07655_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07654_/Y sky130_fd_sc_hd__nand2_1
X_06605_ _08404_/B _06605_/B vssd1 vssd1 vccd1 vccd1 _06609_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08419__A _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07585_ _07586_/A _07586_/B vssd1 vssd1 vccd1 vccd1 _07589_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ _09963_/A _09962_/A _09816_/B _09496_/B vssd1 vssd1 vccd1 vccd1 _09324_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_75_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06536_ _06536_/A _06536_/B vssd1 vssd1 vccd1 vccd1 _06539_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09255_ _09986_/A input19/X vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06467_ _06467_/A _06467_/B _06467_/C vssd1 vssd1 vccd1 vccd1 _06469_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08481__A2 _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ _08206_/A _08206_/B vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__nand2_1
X_05418_ _05418_/A _05419_/A vssd1 vssd1 vccd1 vccd1 _05453_/A sky130_fd_sc_hd__nand2_1
X_09186_ _10442_/A _09186_/B vssd1 vssd1 vccd1 vccd1 _09187_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06398_ _06820_/C vssd1 vssd1 vccd1 vccd1 _06633_/A sky130_fd_sc_hd__inv_2
X_08137_ _08109_/Y _08137_/B vssd1 vssd1 vccd1 vccd1 _08138_/B sky130_fd_sc_hd__nand2b_1
X_05349_ _08420_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__buf_8
XFILLER_0_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07993__A _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08068_ _08171_/B _08068_/B vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07019_ _07021_/A _07021_/B vssd1 vssd1 vccd1 vccd1 _07020_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10030_ _10030_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10032_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08999__A _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10228_ _10226_/Y hold90/A vssd1 vssd1 vccd1 vccd1 _10230_/A sky130_fd_sc_hd__and2b_1
X_10159_ _10161_/C vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__inv_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07370_ _07370_/A _07370_/B _07370_/C vssd1 vssd1 vccd1 vccd1 _07371_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06321_ _06321_/A _06321_/B _06321_/C vssd1 vssd1 vccd1 vccd1 _06646_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09040_ _09042_/C vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06252_ _06695_/A _06696_/B vssd1 vssd1 vccd1 vccd1 _06252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05203_ input44/X vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__buf_12
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06183_ _06183_/A _06183_/B _06183_/C vssd1 vssd1 vccd1 vccd1 _06198_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09942_ _09941_/B _10171_/B _09942_/C vssd1 vssd1 vccd1 vccd1 _10176_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09873_ _09873_/A _09873_/B _09873_/C vssd1 vssd1 vccd1 vccd1 _09874_/A sky130_fd_sc_hd__and3_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _10051_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _09083_/C sky130_fd_sc_hd__nand2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09533__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08755_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__nand2_1
X_05967_ _05957_/Y _06320_/B _05966_/Y vssd1 vssd1 vccd1 vccd1 _05969_/A sky130_fd_sc_hd__a21oi_1
X_07706_ _07710_/B _07706_/B vssd1 vssd1 vccd1 vccd1 _07707_/A sky130_fd_sc_hd__nand2_1
X_08686_ _08686_/A _08686_/B vssd1 vssd1 vccd1 vccd1 _08698_/C sky130_fd_sc_hd__nand2_1
X_05898_ _05898_/A _05898_/B vssd1 vssd1 vccd1 vccd1 _05899_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07637_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07640_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07568_ _07744_/C _07733_/A vssd1 vssd1 vccd1 vccd1 _07569_/B sky130_fd_sc_hd__nand2_1
X_09307_ _09307_/A _09307_/B vssd1 vssd1 vccd1 vccd1 _09343_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06519_ _06519_/A _06519_/B _06519_/C vssd1 vssd1 vccd1 vccd1 _06598_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07499_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__nand2_1
X_09238_ _09239_/B _09242_/A vssd1 vssd1 vccd1 vccd1 _09581_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ _09169_/A _09169_/B vssd1 vssd1 vccd1 vccd1 _09182_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09954__A2 _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06116__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10013_ _10013_/A _10013_/B _10013_/C vssd1 vssd1 vccd1 vccd1 _10016_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_86_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06307__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06870_ _10043_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _07031_/C sky130_fd_sc_hd__nand2_1
X_05821_ _05821_/A _05821_/B vssd1 vssd1 vccd1 vccd1 _05823_/B sky130_fd_sc_hd__and2_1
XANTENNA__09072__B _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08540_ _08540_/A _08540_/B _08540_/C vssd1 vssd1 vccd1 vccd1 _08547_/C sky130_fd_sc_hd__nand3_1
X_05752_ _05752_/A _05752_/B vssd1 vssd1 vccd1 vccd1 _05773_/C sky130_fd_sc_hd__nand2_1
X_08471_ _08673_/B _08471_/B _08471_/C vssd1 vssd1 vccd1 vccd1 _08673_/A sky130_fd_sc_hd__nand3_2
X_05683_ _05694_/B _05683_/B vssd1 vssd1 vccd1 vccd1 _05687_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07422_ _07270_/Y _07421_/Y _07269_/A vssd1 vssd1 vccd1 vccd1 _07508_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07353_ _07202_/A _07225_/B _07203_/A vssd1 vssd1 vccd1 vccd1 _07354_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07284_ _07284_/A _07284_/B _07284_/C vssd1 vssd1 vccd1 vccd1 _07285_/B sky130_fd_sc_hd__nand3_1
X_06304_ _06962_/B _06304_/B vssd1 vssd1 vccd1 vccd1 _06305_/B sky130_fd_sc_hd__nand2_1
X_09023_ _09199_/A _10051_/B _09548_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _09023_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06235_ _06660_/B vssd1 vssd1 vccd1 vccd1 _06661_/A sky130_fd_sc_hd__inv_2
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09528__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06166_ _06166_/A _06166_/B _06166_/C vssd1 vssd1 vccd1 vccd1 _06173_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06097_ _06101_/C vssd1 vssd1 vccd1 vccd1 _06098_/C sky130_fd_sc_hd__inv_2
X_09925_ _09925_/A _09925_/B _09925_/C vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__nand3_1
X_09856_ _10084_/A _10084_/C _10084_/D _09856_/D vssd1 vssd1 vccd1 vccd1 _10091_/B
+ sky130_fd_sc_hd__or4_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08836_/A _08836_/C vssd1 vssd1 vccd1 vccd1 _08835_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05791__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09971_/A _09788_/A vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__or2_1
X_06999_ _07000_/A _06999_/B _06999_/C vssd1 vssd1 vccd1 vccd1 _07004_/A sky130_fd_sc_hd__nand3_1
X_08738_ _08738_/A _08739_/A vssd1 vssd1 vccd1 vccd1 _08754_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08669_ _08669_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08607__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09438__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ _10495_/CLK hold34/X fanout99/X vssd1 vssd1 vccd1 vccd1 _10493_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__08996__B _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10112__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06020_ _06406_/A _06408_/A _06021_/B vssd1 vssd1 vccd1 vccd1 _06049_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05595__B _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07971_ _07971_/A _07971_/B vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__and2_1
X_09710_ _10044_/A _10044_/C _10044_/D _09710_/D vssd1 vssd1 vccd1 vccd1 _10048_/B
+ sky130_fd_sc_hd__or4_1
X_06922_ _07111_/B _07110_/B vssd1 vssd1 vccd1 vccd1 _06922_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09641_ _09641_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__nor2_1
X_06853_ _06853_/A _06853_/B vssd1 vssd1 vccd1 vccd1 _06857_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09572_ _09572_/A _09572_/B _09572_/C vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__nand3_1
X_06784_ _06784_/A _06784_/B vssd1 vssd1 vccd1 vccd1 _06786_/A sky130_fd_sc_hd__nand2_1
X_05804_ _05804_/A _05804_/B vssd1 vssd1 vccd1 vccd1 _06299_/B sky130_fd_sc_hd__nand2_1
X_08523_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08593_/A sky130_fd_sc_hd__nand2_1
X_05735_ _06186_/B _05735_/B vssd1 vssd1 vccd1 vccd1 _05781_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08454_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08458_/C sky130_fd_sc_hd__nand2_1
X_05666_ _05749_/A _05749_/C _05665_/Y vssd1 vssd1 vccd1 vccd1 _06175_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _08391_/A sky130_fd_sc_hd__nand2_1
X_05597_ input36/X _09022_/C vssd1 vssd1 vccd1 vccd1 _06121_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07405_ _07407_/B _07407_/C vssd1 vssd1 vccd1 vccd1 _07643_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07336_ _07332_/Y _07450_/B _07335_/Y vssd1 vssd1 vccd1 vccd1 _07339_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ _09006_/A _09007_/A vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07267_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07423_/C sky130_fd_sc_hd__nand2_1
X_07198_ _07198_/A _07198_/B _07198_/C vssd1 vssd1 vccd1 vccd1 _07199_/B sky130_fd_sc_hd__nand3_1
X_06218_ _06277_/A _06277_/B vssd1 vssd1 vccd1 vccd1 _06276_/A sky130_fd_sc_hd__nand2_1
X_06149_ _06151_/B vssd1 vssd1 vccd1 vccd1 _06150_/B sky130_fd_sc_hd__inv_2
XFILLER_0_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09908_ _09908_/A _09908_/B _09908_/C vssd1 vssd1 vccd1 vccd1 _09914_/C sky130_fd_sc_hd__nand3_1
X_09839_ _09839_/A _09839_/B vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08337__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10476_ _10511_/CLK _10476_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06974__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08247__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05520_ _05539_/B _05539_/C vssd1 vssd1 vccd1 vccd1 _05983_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05451_ _05451_/A _05617_/B _05451_/C vssd1 vssd1 vccd1 vccd1 _05617_/A sky130_fd_sc_hd__nand3_2
X_08170_ _08170_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10387_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07121_ _07121_/A _07121_/B vssd1 vssd1 vccd1 vccd1 _07393_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05382_ _05405_/B _05405_/A vssd1 vssd1 vccd1 vccd1 _05395_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07052_ _07052_/A vssd1 vssd1 vccd1 vccd1 _07054_/B sky130_fd_sc_hd__inv_2
X_06003_ _09962_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _06008_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08710__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ _07954_/A _07954_/B vssd1 vssd1 vccd1 vccd1 _07989_/A sky130_fd_sc_hd__nand2_1
X_06905_ _06907_/B vssd1 vssd1 vccd1 vccd1 _06906_/B sky130_fd_sc_hd__inv_2
XANTENNA__07326__A _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ _07887_/A vssd1 vssd1 vccd1 vccd1 _07886_/A sky130_fd_sc_hd__inv_2
X_09624_ _09916_/A vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__inv_2
X_06836_ _06836_/A _06836_/B vssd1 vssd1 vccd1 vccd1 _06839_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07045__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07550__A2 _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ _09555_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06767_ _06865_/C _06865_/B _06766_/Y vssd1 vssd1 vccd1 vccd1 _06854_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _09486_/A vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__inv_2
X_08506_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08507_/B sky130_fd_sc_hd__inv_2
X_05718_ _05720_/B _05719_/A _05719_/B vssd1 vssd1 vccd1 vccd1 _06185_/B sky130_fd_sc_hd__nand3b_1
X_06698_ _06698_/A _06698_/B vssd1 vssd1 vccd1 vccd1 _06699_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08437_ _08437_/A _08437_/B vssd1 vssd1 vccd1 vccd1 _08441_/C sky130_fd_sc_hd__nand2_1
X_05649_ _05649_/A vssd1 vssd1 vccd1 vccd1 _05650_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ _08368_/A _08368_/B _08368_/C vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08299_ _08300_/B _08300_/A vssd1 vssd1 vccd1 vccd1 _08299_/Y sky130_fd_sc_hd__nand2_1
X_07319_ _07377_/A _07319_/B _07319_/C vssd1 vssd1 vccd1 vccd1 _07339_/B sky130_fd_sc_hd__nand3_1
X_10330_ hold14/X _10322_/Y hold108/X vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10471__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ hold100/A hold24/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__nand2_1
X_10192_ _10193_/B hold86/A vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__or2_1
XANTENNA__06140__A _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__B2 _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__A1 _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput36 b_i[12] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 a_i[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
Xinput14 a_i[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput47 b_i[22] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_1
Xinput58 b_i[3] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10491__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10459_ _10495_/CLK _10459_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07670_ _07691_/B _07691_/A vssd1 vssd1 vccd1 vccd1 _07674_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09361__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ _06196_/C _06196_/B _06399_/Y vssd1 vssd1 vccd1 vccd1 _06622_/B sky130_fd_sc_hd__a21o_1
X_09340_ _09340_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__nand2_1
X_06552_ _10043_/A _09601_/B vssd1 vssd1 vccd1 vccd1 _06553_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09271_ _09762_/A _09270_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09272_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05503_ _05503_/A _05503_/B vssd1 vssd1 vccd1 vccd1 _05503_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _08223_/B _08223_/A vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__or2_1
X_06483_ _06501_/A _08281_/A vssd1 vssd1 vccd1 vccd1 _06500_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10494__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08705__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05434_ _05461_/C _05461_/B _05431_/Y vssd1 vssd1 vccd1 vccd1 _05452_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10508__RESET_B fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08184_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05365_ _05370_/A _05370_/B vssd1 vssd1 vccd1 vccd1 _05369_/A sky130_fd_sc_hd__nand2_1
X_07104_ _07104_/A _07104_/B vssd1 vssd1 vccd1 vccd1 _07104_/Y sky130_fd_sc_hd__nor2_1
X_08084_ _08084_/A vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__inv_2
X_05296_ input62/X vssd1 vssd1 vccd1 vccd1 _08247_/B sky130_fd_sc_hd__clkbuf_8
X_07035_ _10043_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _07178_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06225__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08986_ _08986_/A _08986_/B vssd1 vssd1 vccd1 vccd1 _08990_/C sky130_fd_sc_hd__nand2_1
X_07937_ _08035_/C _08035_/B vssd1 vssd1 vccd1 vccd1 _07980_/B sky130_fd_sc_hd__nand2_1
X_07868_ _07935_/B _07922_/C _07867_/Y vssd1 vssd1 vccd1 vccd1 _07880_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09607_ _09607_/A _09873_/A vssd1 vssd1 vccd1 vccd1 _09611_/C sky130_fd_sc_hd__nand2_1
X_06819_ _07709_/B vssd1 vssd1 vccd1 vccd1 _06820_/B sky130_fd_sc_hd__inv_2
X_07799_ _07799_/A _07799_/B _07799_/C vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__nand3_1
X_09538_ _09702_/A _09703_/A vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__or2_1
XFILLER_0_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09469_ _09469_/A _09469_/B vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08334__B _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ _10498_/Q hold13/X vssd1 vssd1 vccd1 vccd1 _10313_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10244_ _10244_/A hold40/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__nand2_1
X_10175_ _10175_/A vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__inv_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05214__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08838_/Y _08512_/B _08839_/Y vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__a21oi_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08900_/B _08771_/B _08772_/B vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__nand3_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05983_ _05983_/A _05983_/B vssd1 vssd1 vccd1 vccd1 _05983_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09803__B _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _07721_/B _07722_/B _07722_/C vssd1 vssd1 vccd1 vccd1 _07887_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07653_ _08205_/B vssd1 vssd1 vccd1 vccd1 _07677_/B sky130_fd_sc_hd__inv_2
XANTENNA__08419__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06604_ _06604_/A _06604_/B vssd1 vssd1 vccd1 vccd1 _06605_/B sky130_fd_sc_hd__nand2_1
X_09323_ _09960_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07584_ _09601_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _07586_/B sky130_fd_sc_hd__nand2_1
X_06535_ _06535_/A _08365_/B _06538_/A vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_47_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09254_ _09350_/B vssd1 vssd1 vccd1 vccd1 _09348_/A sky130_fd_sc_hd__inv_2
XFILLER_0_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08435__A _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06466_ _08268_/B _06466_/B _06466_/C vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09185_ _10449_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _09186_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08205_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08206_/A sky130_fd_sc_hd__nand2_1
X_05417_ input35/X _09022_/C vssd1 vssd1 vccd1 vccd1 _05419_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08136_ _08136_/A _08161_/A vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06397_ _06641_/A _06641_/B _06397_/C vssd1 vssd1 vccd1 vccd1 _06820_/C sky130_fd_sc_hd__nand3_4
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05348_ _05928_/B _05928_/C vssd1 vssd1 vccd1 vccd1 _05927_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07993__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05279_ _05279_/A _05280_/A vssd1 vssd1 vccd1 vccd1 _05282_/A sky130_fd_sc_hd__nand2_1
X_08067_ _08067_/A _08079_/B vssd1 vssd1 vccd1 vccd1 _08083_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07018_ _07018_/A _07018_/B vssd1 vssd1 vccd1 vccd1 _07021_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05794__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08969_ _09951_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10227_ _10487_/Q hold89/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__nand2_1
X_10158_ _10158_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10161_/C sky130_fd_sc_hd__nor2_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10089_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10093_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06320_ _06320_/A _06320_/B vssd1 vssd1 vccd1 vccd1 _06646_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06251_ _06697_/C vssd1 vssd1 vccd1 vccd1 _06699_/B sky130_fd_sc_hd__inv_2
XFILLER_0_25_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05202_ input10/X vssd1 vssd1 vccd1 vccd1 _09962_/B sky130_fd_sc_hd__clkbuf_8
X_06182_ _06182_/A _06182_/B vssd1 vssd1 vccd1 vccd1 _06198_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09872_ _09872_/A vssd1 vssd1 vccd1 vccd1 _09876_/A sky130_fd_sc_hd__inv_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08828_/B sky130_fd_sc_hd__inv_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09533__B _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08754_ _08754_/A _08754_/B _08754_/C vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__nand3_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05966_ _06316_/A _06318_/A vssd1 vssd1 vccd1 vccd1 _05966_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07705_ _07678_/Y _08209_/B _07704_/Y vssd1 vssd1 vccd1 vccd1 _07714_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08685_ _08428_/B _08428_/A _08674_/B vssd1 vssd1 vccd1 vccd1 _08686_/B sky130_fd_sc_hd__o21a_1
X_05897_ _05897_/A _05897_/B vssd1 vssd1 vccd1 vccd1 _05898_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07636_ _07640_/A _07640_/B vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07567_ _07733_/A _07733_/B _07567_/C vssd1 vssd1 vccd1 vccd1 _07744_/C sky130_fd_sc_hd__nand3_1
X_09306_ _09306_/A _09306_/B vssd1 vssd1 vccd1 vccd1 _09307_/B sky130_fd_sc_hd__and2_1
XANTENNA__05789__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06518_ _06518_/A _08268_/A _06518_/C vssd1 vssd1 vccd1 vccd1 _06519_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _09237_/A _09542_/A vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07498_ _07498_/A vssd1 vssd1 vccd1 vccd1 _07499_/B sky130_fd_sc_hd__inv_2
XFILLER_0_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06449_ _06448_/B _08260_/B _06449_/C vssd1 vssd1 vccd1 vccd1 _08260_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09168_ _09178_/B vssd1 vssd1 vccd1 vccd1 _09169_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _09385_/B _09099_/B _09099_/C vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__nand3_1
X_08119_ _08134_/A _08134_/B _08119_/C vssd1 vssd1 vccd1 vccd1 _08164_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_101_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10012_ _10013_/A _10013_/C _10013_/B vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07244__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05699__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06307__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05820_ _09199_/A _10111_/B _09548_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _05821_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05751_ _05751_/A _05751_/B vssd1 vssd1 vccd1 vccd1 _05752_/A sky130_fd_sc_hd__nand2_1
X_08470_ _08470_/A vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__inv_2
X_05682_ _05685_/B _06126_/A _05686_/A vssd1 vssd1 vccd1 vccd1 _06133_/B sky130_fd_sc_hd__nand3_1
X_07421_ _07423_/C vssd1 vssd1 vccd1 vccd1 _07421_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07352_ _07352_/A _07352_/B vssd1 vssd1 vccd1 vccd1 _07386_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06303_ _06303_/A _06304_/B _06720_/A vssd1 vssd1 vccd1 vccd1 _06962_/B sky130_fd_sc_hd__nand3_1
X_07283_ _07283_/A _07283_/B _07283_/C vssd1 vssd1 vccd1 vccd1 _07284_/B sky130_fd_sc_hd__nand3_1
X_09022_ _09199_/A _09548_/A _09022_/C _09022_/D vssd1 vssd1 vccd1 vccd1 _09024_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06234_ _10052_/A _10000_/A vssd1 vssd1 vccd1 vccd1 _06660_/B sky130_fd_sc_hd__nand2_1
X_06165_ _06165_/A _06165_/B vssd1 vssd1 vccd1 vccd1 _06586_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09528__B _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06096_ _06096_/A _06096_/B vssd1 vssd1 vccd1 vccd1 _06101_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06233__A _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09924_ _09924_/A vssd1 vssd1 vccd1 vccd1 _09925_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09855_ input50/X vssd1 vssd1 vccd1 vccd1 _10084_/C sky130_fd_sc_hd__inv_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08806_/A _08806_/B _09055_/A vssd1 vssd1 vccd1 vccd1 _08836_/C sky130_fd_sc_hd__nand3_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _09971_/B vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__inv_2
X_06998_ _07690_/B _07690_/C vssd1 vssd1 vccd1 vccd1 _07689_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08737_ _08737_/A _08737_/B vssd1 vssd1 vccd1 vccd1 _08739_/A sky130_fd_sc_hd__nand2_1
X_05949_ _05949_/A _05949_/B _05949_/C vssd1 vssd1 vccd1 vccd1 _05950_/A sky130_fd_sc_hd__nand3_1
X_08668_ _09188_/A _08668_/B _08668_/C vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07619_ _07906_/A vssd1 vssd1 vccd1 vccd1 _07620_/C sky130_fd_sc_hd__inv_2
XFILLER_0_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08607__B input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _09147_/A vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__inv_2
XFILLER_0_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ _10494_/CLK _10492_/D fanout99/X vssd1 vssd1 vccd1 vccd1 _10492_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09438__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06143__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__A _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05222__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09629__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07970_ _07970_/A _07970_/B vssd1 vssd1 vccd1 vccd1 _07974_/B sky130_fd_sc_hd__nand2_1
X_06921_ _07112_/C vssd1 vssd1 vccd1 vccd1 _07109_/B sky130_fd_sc_hd__inv_2
X_09640_ _09641_/B _09641_/A vssd1 vssd1 vccd1 vccd1 _09640_/Y sky130_fd_sc_hd__nand2_1
X_06852_ _06854_/A vssd1 vssd1 vccd1 vccd1 _06853_/B sky130_fd_sc_hd__inv_2
X_09571_ _09571_/A _09571_/B vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__nand2_1
X_06783_ _06785_/B _06785_/C vssd1 vssd1 vccd1 vccd1 _06784_/A sky130_fd_sc_hd__nand2_1
X_05803_ _05805_/B vssd1 vssd1 vccd1 vccd1 _05804_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08522_ _08854_/B _08522_/B vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__nand2_1
X_05734_ _06186_/A vssd1 vssd1 vccd1 vccd1 _05735_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08453_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08719_/B sky130_fd_sc_hd__or2_1
X_05665_ _05665_/A _05665_/B vssd1 vssd1 vccd1 vccd1 _05665_/Y sky130_fd_sc_hd__nor2_1
X_07404_ _07403_/B _07404_/B _07404_/C vssd1 vssd1 vccd1 vccd1 _07407_/C sky130_fd_sc_hd__nand3b_1
X_08384_ _08386_/C vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__inv_2
X_05596_ _06121_/A vssd1 vssd1 vccd1 vccd1 _05599_/A sky130_fd_sc_hd__inv_2
XANTENNA__06228__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07335_ _07448_/B _07447_/A vssd1 vssd1 vccd1 vccd1 _07335_/Y sky130_fd_sc_hd__nor2_1
X_07266_ _10083_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _07270_/B sky130_fd_sc_hd__nand2_1
X_09005_ _08747_/Y _08750_/B _08748_/A vssd1 vssd1 vccd1 vccd1 _09007_/A sky130_fd_sc_hd__a21oi_1
X_06217_ _05823_/B _06217_/B _06217_/C vssd1 vssd1 vccd1 vccd1 _06277_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07197_ _07197_/A _07197_/B _07197_/C vssd1 vssd1 vccd1 vccd1 _07198_/B sky130_fd_sc_hd__nand3_1
X_06148_ _05717_/B _05717_/C _05711_/A vssd1 vssd1 vccd1 vccd1 _06151_/B sky130_fd_sc_hd__a21oi_2
X_06079_ _06083_/B _06084_/C _06084_/A vssd1 vssd1 vccd1 vccd1 _06511_/B sky130_fd_sc_hd__nand3_1
X_09907_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _10141_/A sky130_fd_sc_hd__nand2_1
X_09838_ _09840_/C vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__inv_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _09769_/A _09993_/A vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05307__A _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08337__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10475_ _10509_/CLK _10475_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08528__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08247__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05450_ _05454_/C vssd1 vssd1 vccd1 vccd1 _05451_/C sky130_fd_sc_hd__inv_2
XFILLER_0_55_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05381_ _05379_/Y _05369_/B _05380_/Y vssd1 vssd1 vccd1 vccd1 _05405_/A sky130_fd_sc_hd__a21oi_1
X_07120_ _07119_/B _07120_/B _07120_/C vssd1 vssd1 vccd1 vccd1 _07121_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07051_ _07051_/A _07051_/B vssd1 vssd1 vccd1 vccd1 _07054_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09221__B1 _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06002_ _06017_/B _06018_/C _06018_/A vssd1 vssd1 vccd1 vccd1 _06463_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08710__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _07966_/B vssd1 vssd1 vccd1 vccd1 _07954_/B sky130_fd_sc_hd__inv_2
X_07884_ _07882_/Y _07932_/B _07883_/Y vssd1 vssd1 vccd1 vccd1 _08049_/B sky130_fd_sc_hd__a21oi_1
X_06904_ _10050_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _06907_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07326__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _09621_/Y _09382_/B _09622_/Y vssd1 vssd1 vccd1 vccd1 _09916_/A sky130_fd_sc_hd__a21oi_2
X_06835_ _06999_/B _06835_/B vssd1 vssd1 vccd1 vccd1 _06836_/A sky130_fd_sc_hd__nand2_1
X_09554_ _09716_/A _09558_/C vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08438__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06766_ _06862_/B _06861_/A vssd1 vssd1 vccd1 vccd1 _06766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09485_ _09951_/B _09963_/B _09485_/C _09804_/A vssd1 vssd1 vccd1 vccd1 _09486_/A
+ sky130_fd_sc_hd__and4_1
X_08505_ _08503_/Y _08261_/B _08504_/Y vssd1 vssd1 vccd1 vccd1 _08839_/A sky130_fd_sc_hd__a21oi_2
X_05717_ _05717_/A _05717_/B _05717_/C vssd1 vssd1 vccd1 vccd1 _05719_/B sky130_fd_sc_hd__nand3_1
X_06697_ _06697_/A _06697_/B _06697_/C vssd1 vssd1 vccd1 vccd1 _06703_/B sky130_fd_sc_hd__nand3_1
X_08436_ _08437_/A _08437_/B vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__or2_1
X_05648_ _05648_/A _05649_/A vssd1 vssd1 vccd1 vccd1 _05694_/C sky130_fd_sc_hd__nand2_1
X_08367_ _08367_/A vssd1 vssd1 vccd1 vccd1 _08368_/A sky130_fd_sc_hd__inv_2
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07318_ _07377_/B _07318_/B vssd1 vssd1 vccd1 vccd1 _07339_/A sky130_fd_sc_hd__nand2_1
X_05579_ _06065_/A vssd1 vssd1 vccd1 vccd1 _05582_/A sky130_fd_sc_hd__inv_2
XANTENNA__09269__A _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08298_ _08511_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08582_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07249_ _07489_/C _07489_/B _07486_/A vssd1 vssd1 vccd1 vccd1 _07475_/C sky130_fd_sc_hd__a21oi_2
X_10260_ _10260_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09763__A1 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10191_/A _10191_/B vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__nand2_1
XANTENNA__09818__A2 _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07252__A _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput37 b_i[13] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput26 a_i[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 a_i[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
Xinput48 b_i[23] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_1
Xinput59 b_i[4] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10458_ _10494_/CLK _10458_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfrtp_1
X_10389_ _10389_/A vssd1 vssd1 vccd1 vccd1 _10458_/D sky130_fd_sc_hd__clkbuf_1
X_06620_ _08413_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _08655_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09361__B input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ _09361_/D vssd1 vssd1 vccd1 vccd1 _09601_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ _09762_/A _09270_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09270_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06482_ _08281_/B _06482_/B _06482_/C vssd1 vssd1 vccd1 vccd1 _08281_/A sky130_fd_sc_hd__nand3_2
X_05502_ _05502_/A _05502_/B vssd1 vssd1 vccd1 vccd1 _05573_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08221_ _08221_/A _08221_/B vssd1 vssd1 vccd1 vccd1 _08223_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05433_ _05452_/A _05453_/B vssd1 vssd1 vccd1 vccd1 _05451_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08154_/B _08152_/B vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05364_ _05364_/A _05380_/A vssd1 vssd1 vccd1 vccd1 _05370_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07103_ _07103_/A vssd1 vssd1 vccd1 vccd1 _07292_/B sky130_fd_sc_hd__inv_2
X_05295_ _05335_/A _05335_/B vssd1 vssd1 vccd1 vccd1 _05334_/A sky130_fd_sc_hd__nand2_1
X_08083_ _08083_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08084_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09817__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ _07197_/B _07197_/C vssd1 vssd1 vccd1 vccd1 _07196_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06225__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _08985_/A _09337_/A vssd1 vssd1 vccd1 vccd1 _08986_/B sky130_fd_sc_hd__nand2_1
X_07936_ _07936_/A _07936_/B _07936_/C vssd1 vssd1 vccd1 vccd1 _08035_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07867_ _07935_/A vssd1 vssd1 vccd1 vccd1 _07867_/Y sky130_fd_sc_hd__inv_2
X_09606_ _09873_/A _09607_/A vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__or2_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06818_ _06818_/A _07709_/B vssd1 vssd1 vccd1 vccd1 _06821_/A sky130_fd_sc_hd__nand2_1
X_07798_ _07796_/Y _07889_/B _07797_/Y vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__a21o_1
X_09537_ _09698_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__nand2_1
X_06749_ _06749_/A _06749_/B vssd1 vssd1 vccd1 vccd1 _06751_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _09468_/A _09468_/B vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09399_ _09399_/A _09399_/B vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _09986_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _08428_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ _10312_/A hold11/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__xor2_1
XFILLER_0_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10243_ _10241_/Y _10243_/B vssd1 vssd1 vccd1 vccd1 _10250_/A sky130_fd_sc_hd__and2b_1
X_10174_ _10174_/A _10175_/A vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05214__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08525__B _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08770_ _08770_/A _08770_/B vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__nand2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05982_ _05571_/C _05571_/B _05981_/Y vssd1 vssd1 vccd1 vccd1 _06099_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07721_ _07721_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07887_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10461__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _07652_/A _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__nand3_1
X_06603_ _06604_/B _06604_/A vssd1 vssd1 vccd1 vccd1 _08404_/B sky130_fd_sc_hd__or2_1
X_07583_ _08337_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _07586_/A sky130_fd_sc_hd__nand2_1
X_09322_ _09330_/C vssd1 vssd1 vccd1 vccd1 _09322_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_87_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06534_ _06534_/A _06534_/B vssd1 vssd1 vccd1 vccd1 _06538_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09253_ _09253_/A _09253_/B vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06465_ _06468_/A _06467_/A vssd1 vssd1 vccd1 vccd1 _06466_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08435__B _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09184_ _09191_/A vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05416_ input32/X vssd1 vssd1 vccd1 vccd1 _09022_/C sky130_fd_sc_hd__clkbuf_8
X_08204_ _08204_/A vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__inv_2
X_06396_ _06816_/B _06816_/A vssd1 vssd1 vccd1 vccd1 _06397_/C sky130_fd_sc_hd__nor2_1
X_08135_ _08160_/B _08135_/B _08135_/C vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05347_ _05347_/A _05347_/B _05347_/C vssd1 vssd1 vccd1 vccd1 _05928_/C sky130_fd_sc_hd__nand3_1
XANTENNA__06236__A _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09547__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05278_ _09496_/B _09980_/A vssd1 vssd1 vccd1 vccd1 _05280_/A sky130_fd_sc_hd__nand2_1
X_08066_ _08072_/B _08069_/C vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__nand2_1
X_07017_ _07345_/B _07017_/B vssd1 vssd1 vccd1 vccd1 _07018_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05794__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _08968_/A _09230_/A vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09282__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ _09141_/C _08899_/B vssd1 vssd1 vccd1 vccd1 _09069_/A sky130_fd_sc_hd__nand2_1
X_07919_ _08075_/C _08075_/B vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05985__A _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10226_ _10487_/Q hold89/X vssd1 vssd1 vccd1 vccd1 _10226_/Y sky130_fd_sc_hd__nor2_1
X_10157_ _10157_/A vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__inv_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10484__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ _10089_/B _10089_/A vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__or2_1
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06250_ input35/X _08825_/B vssd1 vssd1 vccd1 vccd1 _06697_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06181_ _06183_/C vssd1 vssd1 vccd1 vccd1 _06182_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08271__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09940_ _10171_/B _09942_/C vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__nand2_1
X_09871_ _09878_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__nor2_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _10050_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__nand2_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__nand2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05965_ _06321_/C vssd1 vssd1 vccd1 vccd1 _06320_/B sky130_fd_sc_hd__inv_2
X_07704_ _10416_/B _07703_/Y _07694_/A vssd1 vssd1 vccd1 vccd1 _07704_/Y sky130_fd_sc_hd__o21ai_1
X_08684_ _08684_/A _08911_/A vssd1 vssd1 vccd1 vccd1 _08686_/A sky130_fd_sc_hd__nand2_1
X_05896_ _05898_/B _05897_/B _05897_/A vssd1 vssd1 vccd1 vccd1 _05899_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07635_ _07655_/A _07635_/B _07635_/C vssd1 vssd1 vccd1 vccd1 _07640_/B sky130_fd_sc_hd__nand3_1
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07569_/A sky130_fd_sc_hd__nand2_1
X_09305_ _09308_/B _09479_/A vssd1 vssd1 vccd1 vccd1 _09307_/A sky130_fd_sc_hd__nand2_1
X_06517_ _06517_/A _06517_/B vssd1 vssd1 vccd1 vccd1 _06519_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09236_ _09235_/B _09236_/B _09542_/B vssd1 vssd1 vccd1 vccd1 _09542_/A sky130_fd_sc_hd__nand3b_1
X_07497_ _07497_/A vssd1 vssd1 vccd1 vccd1 _07499_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06448_ _06448_/A _06448_/B vssd1 vssd1 vccd1 vccd1 _06455_/B sky130_fd_sc_hd__nand2_1
X_09167_ _09165_/Y _08644_/B _09166_/Y vssd1 vssd1 vccd1 vccd1 _09178_/B sky130_fd_sc_hd__a21oi_2
X_06379_ _06379_/A _06379_/B vssd1 vssd1 vccd1 vccd1 _06380_/A sky130_fd_sc_hd__nand2_1
X_09098_ _09098_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09104_/B sky130_fd_sc_hd__nand2_1
X_08118_ _08160_/B _08160_/A vssd1 vssd1 vccd1 vccd1 _08119_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08049_ _08049_/A _08049_/B vssd1 vssd1 vccd1 vccd1 _08053_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10011_ _09796_/C _09796_/B _09772_/A vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07244__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05699__B input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09187__A _10437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10126__A input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10209_ hold98/X vssd1 vssd1 vccd1 vccd1 _10484_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07435__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07154__B _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05750_ _05886_/C _05886_/B vssd1 vssd1 vccd1 vccd1 _05888_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05681_ _05448_/C _05448_/B _05678_/Y vssd1 vssd1 vccd1 vccd1 _05685_/B sky130_fd_sc_hd__a21o_1
X_07420_ _07610_/B vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__inv_2
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07351_ _07386_/A _07352_/A _07352_/B vssd1 vssd1 vccd1 vccd1 _07374_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06302_ _06302_/A _06302_/B _06302_/C vssd1 vssd1 vccd1 vccd1 _06656_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ _07315_/B _07315_/A vssd1 vssd1 vccd1 vccd1 _07284_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09021_ _09021_/A vssd1 vssd1 vccd1 vccd1 _09026_/B sky130_fd_sc_hd__inv_2
X_06233_ _08248_/B vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__buf_6
XFILLER_0_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06164_ _06166_/C vssd1 vssd1 vccd1 vccd1 _06165_/B sky130_fd_sc_hd__inv_2
XFILLER_0_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09528__C _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06095_ _06094_/B _06095_/B _06095_/C vssd1 vssd1 vccd1 vccd1 _06096_/B sky130_fd_sc_hd__nand3b_1
X_09923_ _09923_/A _09924_/A vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__nand2_1
X_09854_ input51/X _09854_/B vssd1 vssd1 vccd1 vccd1 _09860_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _09055_/B _08805_/B vssd1 vssd1 vccd1 vccd1 _08836_/A sky130_fd_sc_hd__nand2_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09468_/A _09784_/Y _09467_/A vssd1 vssd1 vccd1 vccd1 _09971_/B sky130_fd_sc_hd__o21a_1
X_06997_ _06997_/A _07146_/B _07146_/C vssd1 vssd1 vccd1 vccd1 _07690_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09857__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ _08740_/B _08740_/C vssd1 vssd1 vccd1 vccd1 _08738_/A sky130_fd_sc_hd__nand2_1
X_05948_ _05948_/A _05948_/B vssd1 vssd1 vccd1 vccd1 _05949_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09560__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08667_ _09188_/B _09188_/A vssd1 vssd1 vccd1 vccd1 _08669_/A sky130_fd_sc_hd__nand2_1
X_05879_ _05760_/Y _05879_/B _05879_/C vssd1 vssd1 vccd1 vccd1 _05880_/B sky130_fd_sc_hd__nand3b_1
X_07618_ _07914_/B vssd1 vssd1 vccd1 vccd1 _07621_/B sky130_fd_sc_hd__inv_2
XANTENNA__08607__C _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ _08596_/Y _08385_/B _08597_/Y vssd1 vssd1 vccd1 vccd1 _09147_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07549_ _08810_/B input44/X vssd1 vssd1 vccd1 vccd1 _07553_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08904__A _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _10026_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _09224_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10491_ _10494_/CLK hold26/X fanout99/X vssd1 vssd1 vccd1 vccd1 _10491_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__09438__C _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06143__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__B _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08814__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05222__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__B input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07149__B _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09000__A1 _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06920_ _09951_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _07112_/C sky130_fd_sc_hd__nand2_1
X_06851_ _07008_/B _07008_/C vssd1 vssd1 vccd1 vccd1 _07007_/A sky130_fd_sc_hd__nand2_1
X_09570_ _09572_/B vssd1 vssd1 vccd1 vccd1 _09571_/B sky130_fd_sc_hd__inv_2
X_06782_ _06782_/A _06782_/B _06782_/C vssd1 vssd1 vccd1 vccd1 _06785_/C sky130_fd_sc_hd__nand3_1
X_05802_ _09528_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _05805_/B sky130_fd_sc_hd__nand2_1
X_08521_ _08521_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _08522_/B sky130_fd_sc_hd__nand2_1
X_05733_ _05731_/Y _05492_/A _05732_/Y vssd1 vssd1 vccd1 vccd1 _06186_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08452_ _09963_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _08454_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05664_ _05773_/B _05751_/A vssd1 vssd1 vccd1 vccd1 _05749_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07403_ _07403_/A _07403_/B vssd1 vssd1 vccd1 vccd1 _07407_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08383_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08386_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05595_ input37/X _09022_/D vssd1 vssd1 vccd1 vccd1 _06121_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06228__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07334_ _07451_/B vssd1 vssd1 vccd1 vccd1 _07450_/B sky130_fd_sc_hd__inv_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07265_ _09854_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__nand2_1
X_09004_ _09008_/A _09233_/A vssd1 vssd1 vccd1 vccd1 _09006_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06216_ _06216_/A _06216_/B vssd1 vssd1 vccd1 vccd1 _06217_/C sky130_fd_sc_hd__nand2_1
X_07196_ _07196_/A _07196_/B vssd1 vssd1 vccd1 vccd1 _07198_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06147_ _06151_/A _06151_/C vssd1 vssd1 vccd1 vccd1 _06150_/A sky130_fd_sc_hd__nand2_1
X_06078_ _06078_/A _06078_/B vssd1 vssd1 vccd1 vccd1 _06084_/A sky130_fd_sc_hd__nand2_1
X_09906_ _09908_/B vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__inv_2
X_09837_ _09837_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09840_/C sky130_fd_sc_hd__nand2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _09993_/B _09768_/B _09768_/C vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__nand3_1
XANTENNA__05307__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _08719_/A _08719_/B vssd1 vssd1 vccd1 vccd1 _08720_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09699_ _10023_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _09701_/A sky130_fd_sc_hd__nand2_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06138__B _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06154__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ _10511_/CLK _10474_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05993__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08528__B _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05233__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05380_ _05380_/A _05380_/B vssd1 vssd1 vccd1 vccd1 _05380_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07050_ _07050_/A _07050_/B _07052_/A vssd1 vssd1 vccd1 vccd1 _07055_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_42_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06001_ _05515_/C _05515_/B _05998_/Y vssd1 vssd1 vccd1 vccd1 _06017_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09221__B2 _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A1 _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07952_ _08003_/A _08003_/B _07951_/A vssd1 vssd1 vccd1 vccd1 _07966_/B sky130_fd_sc_hd__o21ai_1
X_07883_ _07921_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _07883_/Y sky130_fd_sc_hd__nor2_1
X_06903_ _06907_/A vssd1 vssd1 vccd1 vccd1 _06906_/A sky130_fd_sc_hd__inv_2
XANTENNA__05408__A _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ _09622_/A _09622_/B vssd1 vssd1 vccd1 vccd1 _09622_/Y sky130_fd_sc_hd__nor2_1
X_06834_ _06835_/B _06834_/B _06834_/C vssd1 vssd1 vccd1 vccd1 _06999_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_37_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09553_ _09553_/A _09553_/B vssd1 vssd1 vccd1 vccd1 _09558_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08438__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08504_/Y sky130_fd_sc_hd__nor2_1
X_06765_ _06863_/C vssd1 vssd1 vccd1 vccd1 _06865_/B sky130_fd_sc_hd__inv_2
X_09484_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09495_/B sky130_fd_sc_hd__nand2_1
X_05716_ _05716_/A vssd1 vssd1 vccd1 vccd1 _05717_/C sky130_fd_sc_hd__inv_2
XANTENNA__06239__A _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ _06698_/A _06696_/B vssd1 vssd1 vccd1 vccd1 _06697_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _09981_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _08437_/B sky130_fd_sc_hd__nand2_1
X_05647_ _10026_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _05649_/A sky130_fd_sc_hd__nand2_1
X_08366_ _08366_/A _08367_/A vssd1 vssd1 vccd1 vccd1 _08371_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07317_ _07377_/A vssd1 vssd1 vccd1 vccd1 _07318_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05578_ input3/X _09313_/D vssd1 vssd1 vccd1 vccd1 _06065_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09269__B input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ _08297_/A _08297_/B _08297_/C vssd1 vssd1 vccd1 vccd1 _08304_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07248_ _07248_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _07486_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07179_ _07179_/A _07179_/B _07179_/C vssd1 vssd1 vccd1 vccd1 _07182_/A sky130_fd_sc_hd__nand3_1
X_10190_ _10190_/A hold18/X vssd1 vssd1 vccd1 vccd1 _10193_/B sky130_fd_sc_hd__and2_1
XFILLER_0_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05318__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08348__B _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07252__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05988__A _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 a_i[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 a_i[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
Xinput49 b_i[24] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_4
Xinput38 b_i[14] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_2
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10457_ _10457_/A _10457_/B vssd1 vssd1 vccd1 vccd1 _10478_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10388_ _10390_/A _10388_/B vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__and2_1
XANTENNA__09361__C _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06550_ _08322_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06553_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06481_ _06481_/A vssd1 vssd1 vccd1 vccd1 _06482_/C sky130_fd_sc_hd__inv_2
XFILLER_0_47_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05501_ _05335_/C _05499_/Y _05500_/Y vssd1 vssd1 vccd1 vccd1 _05627_/B sky130_fd_sc_hd__o21bai_1
X_08220_ _08220_/A vssd1 vssd1 vccd1 vccd1 _08221_/B sky130_fd_sc_hd__inv_2
XFILLER_0_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05432_ _05461_/C _05461_/B _05431_/Y vssd1 vssd1 vccd1 vccd1 _05453_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08151_ _08151_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _08152_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05363_ _05380_/B vssd1 vssd1 vccd1 vccd1 _05364_/A sky130_fd_sc_hd__inv_2
XFILLER_0_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05294_ _05294_/A _05500_/B vssd1 vssd1 vccd1 vccd1 _05335_/B sky130_fd_sc_hd__nand2_1
X_07102_ _09951_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _07103_/A sky130_fd_sc_hd__nand2_1
X_08082_ _08082_/A vssd1 vssd1 vccd1 vccd1 _10394_/B sky130_fd_sc_hd__inv_2
XFILLER_0_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07033_ _07033_/A _07033_/B _07033_/C vssd1 vssd1 vccd1 vccd1 _07197_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09817__B _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06522__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08984_ _08958_/Y _08720_/B _08959_/Y vssd1 vssd1 vccd1 vccd1 _08986_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07935_ _07935_/A _07935_/B vssd1 vssd1 vccd1 vccd1 _07936_/A sky130_fd_sc_hd__nand2_1
X_09605_ _09873_/C _09873_/B vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__nand2_1
X_07866_ _07866_/A _07866_/B vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__nand2_2
X_06817_ _07153_/A _06817_/B _07153_/B vssd1 vssd1 vccd1 vccd1 _07709_/B sky130_fd_sc_hd__nand3_4
X_07797_ _07887_/A _07886_/B vssd1 vssd1 vccd1 vccd1 _07797_/Y sky130_fd_sc_hd__nor2_1
X_09536_ _09536_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__nand2_1
X_06748_ _06842_/B _06842_/C vssd1 vssd1 vccd1 vccd1 _06841_/A sky130_fd_sc_hd__nand2_1
X_09467_ _09467_/A _09784_/A vssd1 vssd1 vccd1 vccd1 _09468_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08418_ _08312_/A _08312_/B _08521_/B vssd1 vssd1 vccd1 vccd1 _08854_/A sky130_fd_sc_hd__a21boi_1
X_06679_ _06892_/B _06891_/B vssd1 vssd1 vccd1 vccd1 _06680_/C sky130_fd_sc_hd__nand2_1
X_09398_ _09648_/A _09404_/B vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08349_ _09528_/A _09022_/C vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10311_ _10311_/A hold10/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__nand2_1
X_10242_ _10489_/Q _10467_/Q vssd1 vssd1 vccd1 vccd1 _10243_/B sky130_fd_sc_hd__nand2_1
X_10173_ _10173_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _10509_/CLK hold2/X fanout99/A vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__08822__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07438__A _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07157__B _07709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _07722_/B _07722_/C vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__nand2_1
X_05981_ _05981_/A _05981_/B vssd1 vssd1 vccd1 vccd1 _05981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07651_ _07651_/A _07697_/A _07651_/C vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__nand3_2
X_06602_ _06151_/B _06150_/A _06163_/A vssd1 vssd1 vccd1 vccd1 _06604_/A sky130_fd_sc_hd__o21a_1
X_07582_ _10111_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _07765_/B sky130_fd_sc_hd__nand2_1
X_09321_ _09321_/A _09321_/B vssd1 vssd1 vccd1 vccd1 _09330_/C sky130_fd_sc_hd__nand2_1
X_06533_ _06537_/A _08361_/A _06536_/B vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _09251_/B _09252_/B _09252_/C vssd1 vssd1 vccd1 vccd1 _09253_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_62_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06464_ _06016_/A _06016_/C _06463_/Y vssd1 vssd1 vccd1 vccd1 _06467_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ _09183_/A _10448_/B vssd1 vssd1 vccd1 vccd1 _09191_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08203_ _08205_/B _08203_/B vssd1 vssd1 vccd1 vccd1 _08204_/A sky130_fd_sc_hd__xor2_1
X_06395_ _06643_/C _06643_/B vssd1 vssd1 vccd1 vccd1 _06816_/A sky130_fd_sc_hd__nand2_1
X_05415_ _05420_/A _05420_/C vssd1 vssd1 vccd1 vccd1 _05418_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08134_ _08134_/A _08134_/B vssd1 vssd1 vccd1 vccd1 _08136_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05346_ _05346_/A _05346_/B vssd1 vssd1 vccd1 vccd1 _05347_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06236__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09547__B _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05277_ _07960_/B vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__buf_8
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ _08065_/A _08065_/B vssd1 vssd1 vccd1 vccd1 _08069_/C sky130_fd_sc_hd__nand2_1
X_07016_ _07017_/B _07016_/B _07016_/C vssd1 vssd1 vccd1 vccd1 _07345_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08967_ _08967_/A _08967_/B vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09282__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ _08856_/Y _09143_/B _08897_/Y vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__a21o_1
X_07918_ _07918_/A _07918_/B _08206_/B vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__nand3_1
X_07849_ _07849_/A _07849_/B vssd1 vssd1 vccd1 vccd1 _07855_/B sky130_fd_sc_hd__nand2_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ _09523_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08907__A _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05985__B _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10225_ hold74/X vssd1 vssd1 vccd1 vccd1 _10486_/D sky130_fd_sc_hd__clkbuf_1
X_10156_ _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__nor2_1
X_10087_ _10087_/A _10087_/B vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__xnor2_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05241__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06180_ _06180_/A _06180_/B vssd1 vssd1 vccd1 vccd1 _06183_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_13_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08271__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09870_ _09877_/C _10100_/A vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__nand2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08832_/A _08832_/C vssd1 vssd1 vccd1 vccd1 _08830_/A sky130_fd_sc_hd__nand2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08754_/C vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__inv_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05964_ _05964_/A _05964_/B vssd1 vssd1 vccd1 vccd1 _06321_/C sky130_fd_sc_hd__nand2_1
X_08683_ _08683_/A _08684_/A _08911_/A vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__nand3_1
X_07703_ _07703_/A vssd1 vssd1 vccd1 vccd1 _07703_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07634_ _07655_/B _07634_/B vssd1 vssd1 vccd1 vccd1 _07640_/A sky130_fd_sc_hd__nand2_1
X_05895_ _05895_/A _05895_/B vssd1 vssd1 vccd1 vccd1 _05897_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07565_ _07577_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07808_/B sky130_fd_sc_hd__xor2_1
X_09304_ _09479_/B _09304_/B _09304_/C vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__nand3_1
X_06516_ _08317_/B _06516_/B _06516_/C vssd1 vssd1 vccd1 vccd1 _08317_/A sky130_fd_sc_hd__nand3_2
X_07496_ _07556_/B vssd1 vssd1 vccd1 vccd1 _07496_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06247__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09235_ _09235_/A _09235_/B vssd1 vssd1 vccd1 vccd1 _09237_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06447_ _09496_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _06448_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09166_ _09166_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09166_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06378_ _06380_/B _06379_/A _06379_/B vssd1 vssd1 vccd1 vccd1 _06381_/A sky130_fd_sc_hd__nand3b_1
X_09097_ _09099_/C vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__inv_2
X_08117_ _08135_/B _08135_/C vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05329_ _05329_/A _05559_/A _05576_/A vssd1 vssd1 vccd1 vccd1 _05331_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08048_ _08048_/A _08048_/B _08048_/C vssd1 vssd1 vccd1 vccd1 _08056_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10010_ _10010_/A _10010_/B _10010_/C vssd1 vssd1 vccd1 vccd1 _10013_/C sky130_fd_sc_hd__nand3_1
X_09999_ _09999_/A input17/X vssd1 vssd1 vccd1 vccd1 _10001_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10126__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__B1 _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ hold97/X _10213_/A vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__and2_1
X_10139_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07435__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__B1 _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05680_ _06107_/B _06107_/A vssd1 vssd1 vccd1 vccd1 _05684_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ _07350_/A _07350_/B _07350_/C vssd1 vssd1 vccd1 vccd1 _07352_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06301_ _06302_/C _06302_/B vssd1 vssd1 vccd1 vccd1 _06305_/A sky130_fd_sc_hd__nand2_1
X_09020_ _10043_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07281_ _07284_/C _07281_/B _07281_/C vssd1 vssd1 vccd1 vccd1 _07285_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06232_ _06365_/A _06366_/A vssd1 vssd1 vccd1 vccd1 _06232_/Y sky130_fd_sc_hd__nand2_1
X_06163_ _06163_/A _06163_/B vssd1 vssd1 vccd1 vccd1 _06166_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09528__D _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06094_ _06094_/A _06094_/B vssd1 vssd1 vccd1 vccd1 _06096_/A sky130_fd_sc_hd__nand2_1
X_09922_ _10157_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09924_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ _09873_/C _09853_/B vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__nand2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _09784_/A vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__inv_2
X_08804_ _09055_/A vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__inv_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _08735_/A _08735_/B _08735_/C vssd1 vssd1 vccd1 vccd1 _08740_/C sky130_fd_sc_hd__nand3_1
X_06996_ _06996_/A _07146_/A vssd1 vssd1 vccd1 vccd1 _07690_/B sky130_fd_sc_hd__nand2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09857__B2 _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05947_ _05947_/A _05947_/B vssd1 vssd1 vccd1 vccd1 _05949_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09560__B _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _08668_/B _08668_/C vssd1 vssd1 vccd1 vccd1 _09188_/B sky130_fd_sc_hd__nand2_1
X_05878_ _05760_/Y _05877_/Y _05759_/A vssd1 vssd1 vccd1 vccd1 _05880_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08597_ _08597_/A _08597_/B vssd1 vssd1 vccd1 vccd1 _08597_/Y sky130_fd_sc_hd__nor2_1
X_07617_ _07906_/A _07617_/B _07906_/B vssd1 vssd1 vccd1 vccd1 _07914_/B sky130_fd_sc_hd__nand3_2
XANTENNA__08607__D _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07548_ _08422_/A vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10474__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ _07539_/B _07539_/C vssd1 vssd1 vccd1 vccd1 _07542_/A sky130_fd_sc_hd__nand2_1
X_09218_ _09242_/B vssd1 vssd1 vccd1 vccd1 _09239_/B sky130_fd_sc_hd__inv_2
XANTENNA__09288__A input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10490_ _10494_/CLK _10490_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfrtp_1
X_09149_ _09161_/A _09162_/A vssd1 vssd1 vccd1 vccd1 _09171_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09438__D _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09751__A _09751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09198__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08814__B _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09629__C _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07149__C _07150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06850_ _06850_/A _06850_/B _06850_/C vssd1 vssd1 vccd1 vccd1 _07008_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05801_ _05805_/A vssd1 vssd1 vccd1 vccd1 _05804_/A sky130_fd_sc_hd__inv_2
X_06781_ _06781_/A _06781_/B vssd1 vssd1 vccd1 vccd1 _06785_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08520_ _08520_/A _08672_/A vssd1 vssd1 vccd1 vccd1 _08854_/B sky130_fd_sc_hd__nand2_1
X_05732_ _05732_/A _05732_/B vssd1 vssd1 vccd1 vccd1 _05732_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08451_ _09962_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__nand2_1
X_05663_ _05752_/B _05751_/A _05751_/B vssd1 vssd1 vccd1 vccd1 _05773_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10497__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07403_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_85_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08382_ _08381_/B _08382_/B _08382_/C vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__nand3b_1
X_05594_ _05609_/B _05610_/C _05610_/A vssd1 vssd1 vccd1 vccd1 _06093_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07333_ _09963_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _07451_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07264_ _07468_/B _07467_/A vssd1 vssd1 vccd1 vccd1 _07264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09003_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__nand2_1
X_06215_ _06302_/B _06298_/B vssd1 vssd1 vccd1 vccd1 _06216_/A sky130_fd_sc_hd__nand2_1
X_07195_ _07346_/B _07195_/B _07195_/C vssd1 vssd1 vccd1 vccd1 _07346_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_13_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06146_ _06146_/A _06146_/B _06146_/C vssd1 vssd1 vccd1 vccd1 _06151_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06077_ _06077_/A _06077_/B vssd1 vssd1 vccd1 vccd1 _06078_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _09905_/A _10168_/B vssd1 vssd1 vccd1 vccd1 _09908_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ _09840_/A _10019_/A vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__nand2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _09993_/B _09768_/C _09768_/B vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__a21o_1
X_06979_ _07098_/B _07096_/A vssd1 vssd1 vccd1 vccd1 _07399_/A sky130_fd_sc_hd__and2_1
XFILLER_0_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ _09698_/A _09698_/B vssd1 vssd1 vccd1 vccd1 _10023_/B sky130_fd_sc_hd__nand2_1
X_08718_ _08721_/B _08721_/C vssd1 vssd1 vccd1 vccd1 _08720_/A sky130_fd_sc_hd__nand2_1
X_08649_ _09181_/B _09181_/A vssd1 vssd1 vccd1 vccd1 _08660_/C sky130_fd_sc_hd__nand2_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06138__C _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06154__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10473_ _10509_/CLK _10473_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05993__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07266__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__A _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08825__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06345__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06000_ _06017_/A _06018_/B vssd1 vssd1 vccd1 vccd1 _06016_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09221__A2 _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07951_ _07951_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _08003_/B sky130_fd_sc_hd__nand2_1
X_06902_ _09720_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _06907_/A sky130_fd_sc_hd__nand2_1
X_07882_ _07930_/B _07921_/A vssd1 vssd1 vccd1 vccd1 _07882_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05408__B _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ _09622_/B _09622_/A vssd1 vssd1 vccd1 vccd1 _09621_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09391__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ _06841_/B _06842_/B _06842_/C vssd1 vssd1 vccd1 vccd1 _06835_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09552_ _09553_/B _09553_/A vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__or2_1
X_06764_ _09533_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _06863_/C sky130_fd_sc_hd__nand2_1
X_08503_ _08504_/B _08504_/A vssd1 vssd1 vccd1 vccd1 _08503_/Y sky130_fd_sc_hd__nand2_1
X_05715_ _05715_/A _05716_/A vssd1 vssd1 vccd1 vccd1 _05719_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05424__A _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _09518_/B _09837_/B vssd1 vssd1 vccd1 vccd1 _09517_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06239__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06695_ _06695_/A vssd1 vssd1 vccd1 vccd1 _06698_/A sky130_fd_sc_hd__inv_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ _09981_/B _09437_/B vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05646_ input26/X vssd1 vssd1 vccd1 vccd1 _09361_/D sky130_fd_sc_hd__buf_6
X_08365_ _08365_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__nand2_1
X_05577_ _05327_/A _05330_/A _05576_/Y vssd1 vssd1 vccd1 vccd1 _06169_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07316_ _07284_/A _07284_/C _07315_/Y vssd1 vssd1 vccd1 vccd1 _07377_/A sky130_fd_sc_hd__a21oi_2
X_08296_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07247_ _07488_/B vssd1 vssd1 vccd1 vccd1 _07489_/B sky130_fd_sc_hd__inv_2
X_07178_ _07180_/B _07178_/B vssd1 vssd1 vccd1 vccd1 _07179_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06129_ _06129_/A _06129_/B _06534_/A vssd1 vssd1 vccd1 vccd1 _06131_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05318__B _08247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _09817_/X _09819_/B vssd1 vssd1 vccd1 vccd1 _09820_/B sky130_fd_sc_hd__and2b_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05988__B _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 a_i[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
Xinput17 a_i[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_4
Xinput39 b_i[15] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
X_10456_ _10456_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10477_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10387_ _10387_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10388_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05509__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09361__D _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06480_ _06480_/A _06481_/A vssd1 vssd1 vccd1 vccd1 _06501_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05500_ _05500_/A _05500_/B vssd1 vssd1 vccd1 vccd1 _05500_/Y sky130_fd_sc_hd__nor2_1
X_05431_ _05462_/B _05463_/B vssd1 vssd1 vccd1 vccd1 _05431_/Y sky130_fd_sc_hd__nor2_1
X_08150_ _08150_/A vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05362_ _05362_/A _05380_/B vssd1 vssd1 vccd1 vccd1 _05370_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07101_ _07104_/A _07104_/B vssd1 vssd1 vccd1 vccd1 _07292_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05293_ _05502_/A _05293_/B vssd1 vssd1 vccd1 vccd1 _05500_/B sky130_fd_sc_hd__nand2_1
X_08081_ _10397_/B _08081_/B vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07032_ _07032_/A _07032_/B vssd1 vssd1 vccd1 vccd1 _07033_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09817__C _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06522__B _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08983_ _08983_/A _09337_/A _08985_/A vssd1 vssd1 vccd1 vccd1 _08990_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07934_ _07986_/A _07986_/C vssd1 vssd1 vccd1 vccd1 _07984_/A sky130_fd_sc_hd__nand2_1
X_07865_ _07865_/A vssd1 vssd1 vccd1 vccd1 _07866_/B sky130_fd_sc_hd__inv_2
X_09604_ _09604_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06816_ _06816_/A _06816_/B vssd1 vssd1 vccd1 vccd1 _07153_/B sky130_fd_sc_hd__nand2_2
X_07796_ _07886_/B _07887_/A vssd1 vssd1 vccd1 vccd1 _07796_/Y sky130_fd_sc_hd__nand2_1
X_09535_ _09535_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _09698_/A sky130_fd_sc_hd__nand2_1
X_06747_ _06747_/A _06747_/B _06747_/C vssd1 vssd1 vccd1 vccd1 _06842_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ _09981_/A input19/X _09981_/B input18/X vssd1 vssd1 vccd1 vccd1 _09784_/A
+ sky130_fd_sc_hd__a22o_1
X_06678_ _06893_/C vssd1 vssd1 vccd1 vccd1 _06680_/B sky130_fd_sc_hd__inv_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08417_ _08415_/Y _08654_/B _08416_/Y vssd1 vssd1 vccd1 vccd1 _08646_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_19_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05629_ _05629_/A _05629_/B _05629_/C vssd1 vssd1 vccd1 vccd1 _05631_/B sky130_fd_sc_hd__nand3_1
X_09397_ _09397_/A _09397_/B _09397_/C vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10028__B1 _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ input40/X _09022_/D vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__nand2_1
X_08279_ _08279_/A _08279_/B vssd1 vssd1 vccd1 vccd1 _08284_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09296__A _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10310_ _10308_/Y hold118/A vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__and2b_1
X_10241_ _10489_/Q _10467_/Q vssd1 vssd1 vccd1 vccd1 _10241_/Y sky130_fd_sc_hd__nor2_1
X_10172_ _10171_/B _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _10173_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10508_ _10509_/CLK _10508_/D fanout99/A vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__08822__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ _10439_/A vssd1 vssd1 vccd1 vccd1 _10472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07438__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05239__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07157__C _07709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05980_ _05626_/C _05626_/B _05979_/Y vssd1 vssd1 vccd1 vccd1 _06402_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07650_ _07913_/B vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__inv_2
X_06601_ _06616_/B _08388_/A _06617_/C vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__nand3_1
X_07581_ _07592_/B _07600_/B vssd1 vssd1 vccd1 vccd1 _07591_/A sky130_fd_sc_hd__nand2_1
X_09320_ _09321_/B _09321_/A vssd1 vssd1 vccd1 vccd1 _09320_/Y sky130_fd_sc_hd__nor2_1
X_06532_ _06537_/C vssd1 vssd1 vccd1 vccd1 _06536_/B sky130_fd_sc_hd__inv_2
X_09251_ _09251_/A _09251_/B vssd1 vssd1 vccd1 vccd1 _09253_/A sky130_fd_sc_hd__nand2_1
X_06463_ _06463_/A vssd1 vssd1 vccd1 vccd1 _06463_/Y sky130_fd_sc_hd__inv_2
X_08202_ _08202_/A _08202_/B vssd1 vssd1 vccd1 vccd1 _10407_/B sky130_fd_sc_hd__nand2_2
X_09182_ _09182_/A _09182_/B _09182_/C vssd1 vssd1 vccd1 vccd1 _10448_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06394_ _05974_/Y _06394_/B _06394_/C vssd1 vssd1 vccd1 vccd1 _06643_/B sky130_fd_sc_hd__nand3b_1
X_05414_ _05590_/A _05590_/B vssd1 vssd1 vccd1 vccd1 _05420_/C sky130_fd_sc_hd__nand2_1
X_08133_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__nand2_1
X_05345_ _05345_/A _05345_/B _05345_/C vssd1 vssd1 vccd1 vccd1 _05928_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08732__B _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _08064_/A _08064_/B _08064_/C vssd1 vssd1 vccd1 vccd1 _08072_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _07023_/B _07024_/C _07024_/B vssd1 vssd1 vccd1 vccd1 _07017_/B sky130_fd_sc_hd__nand3_1
X_05276_ _05281_/A _05281_/C vssd1 vssd1 vccd1 vccd1 _05279_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08966_ _08967_/B _08967_/A vssd1 vssd1 vccd1 vccd1 _08968_/A sky130_fd_sc_hd__or2_1
XANTENNA__09282__C _09437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ _09141_/A _09140_/A vssd1 vssd1 vccd1 vccd1 _08897_/Y sky130_fd_sc_hd__nor2_1
X_07917_ _08071_/B vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__inv_2
XFILLER_0_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07848_ _07865_/A _07941_/B _07938_/A vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__nand3_1
X_09518_ _09517_/B _09518_/B _09837_/B vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _07855_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _07789_/C sky130_fd_sc_hd__nand2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09451_/A _09451_/C _09451_/B vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06443__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ hold73/X _10229_/A vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__and2_1
X_10155_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10087_/B sky130_fd_sc_hd__nand2_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05522__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05241__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08820_ _08820_/A _08820_/B vssd1 vssd1 vccd1 vccd1 _08832_/C sky130_fd_sc_hd__nand2_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07184__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08751_ _08751_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08754_/C sky130_fd_sc_hd__nand2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05963_ _05962_/B _05963_/B _05963_/C vssd1 vssd1 vccd1 vccd1 _05964_/B sky130_fd_sc_hd__nand3b_1
X_08682_ _08911_/B _08682_/B _08682_/C vssd1 vssd1 vccd1 vccd1 _08911_/A sky130_fd_sc_hd__nand3_1
X_07702_ _10417_/A _10410_/A vssd1 vssd1 vccd1 vccd1 _08209_/B sky130_fd_sc_hd__nor2_1
X_05894_ _05894_/A vssd1 vssd1 vccd1 vccd1 _05895_/B sky130_fd_sc_hd__inv_2
X_07633_ _07655_/A vssd1 vssd1 vccd1 vccd1 _07634_/B sky130_fd_sc_hd__inv_2
XFILLER_0_88_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07564_ _07562_/Y _07564_/B vssd1 vssd1 vccd1 vccd1 _07761_/B sky130_fd_sc_hd__nand2b_1
X_09303_ _09303_/A vssd1 vssd1 vccd1 vccd1 _09304_/C sky130_fd_sc_hd__inv_2
X_06515_ _06519_/C vssd1 vssd1 vccd1 vccd1 _06516_/C sky130_fd_sc_hd__inv_2
XFILLER_0_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07495_ _07497_/A _07498_/A vssd1 vssd1 vccd1 vccd1 _07556_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09234_ _09234_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09235_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06446_ _08260_/B _06449_/C vssd1 vssd1 vccd1 vccd1 _06448_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06247__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09165_ _09166_/B _09166_/A vssd1 vssd1 vccd1 vccd1 _09165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08116_ _08116_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _08135_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06377_ _06377_/A _06377_/B _06377_/C vssd1 vssd1 vccd1 vccd1 _06379_/B sky130_fd_sc_hd__nand3_1
X_09096_ _09096_/A _09096_/B vssd1 vssd1 vccd1 vccd1 _09099_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05328_ _05576_/B _05328_/B vssd1 vssd1 vccd1 vccd1 _05331_/A sky130_fd_sc_hd__nand2_1
X_08047_ _07882_/Y _07932_/B _07883_/Y vssd1 vssd1 vccd1 vccd1 _08048_/A sky130_fd_sc_hd__a21o_1
X_05259_ _09962_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _05265_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09998_ _09998_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _10002_/A sky130_fd_sc_hd__nand2_1
X_08949_ _09332_/A _08949_/B vssd1 vssd1 vccd1 vccd1 _08951_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08918__A _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06173__A _06173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09563__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06901__A _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__B2 _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__nand2_1
X_10138_ _10138_/A _10138_/B _10138_/C vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__nand3_1
X_10069_ _09706_/B _09701_/Y _09738_/A vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09315__B2 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__A1 _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06348__A _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07280_ _07283_/A _07283_/C _07315_/A vssd1 vssd1 vccd1 vccd1 _07281_/C sky130_fd_sc_hd__nand3_1
X_06300_ _06300_/A _06300_/B vssd1 vssd1 vccd1 vccd1 _06302_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06231_ _06358_/C _06358_/B _06230_/Y vssd1 vssd1 vccd1 vccd1 _06366_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06162_ _06162_/A _06162_/B _06162_/C vssd1 vssd1 vccd1 vccd1 _06163_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06093_ _06093_/A _06093_/B vssd1 vssd1 vccd1 vccd1 _06094_/B sky130_fd_sc_hd__nand2_1
X_09921_ _09921_/A _09921_/B _09921_/C vssd1 vssd1 vccd1 vccd1 _09922_/B sky130_fd_sc_hd__nand3_1
X_09852_ _09850_/Y _09567_/B _09851_/Y vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__a21oi_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09996_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__nand2_1
X_08803_ _08801_/Y _08539_/A _08802_/Y vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__a21oi_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05427__A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__B input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _08735_/A _08735_/C _08735_/B vssd1 vssd1 vccd1 vccd1 _08740_/B sky130_fd_sc_hd__a21o_1
X_06995_ _06997_/A vssd1 vssd1 vccd1 vccd1 _07146_/A sky130_fd_sc_hd__inv_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09857__A2 _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05946_ _06333_/A _06334_/A vssd1 vssd1 vccd1 vccd1 _06325_/B sky130_fd_sc_hd__nand2_1
X_08665_ _08665_/A _08665_/B vssd1 vssd1 vccd1 vccd1 _08668_/B sky130_fd_sc_hd__nand2_1
X_05877_ _05879_/C vssd1 vssd1 vccd1 vccd1 _05877_/Y sky130_fd_sc_hd__inv_2
X_08596_ _08597_/B _08597_/A vssd1 vssd1 vccd1 vccd1 _08596_/Y sky130_fd_sc_hd__nand2_1
X_07616_ _07616_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _07906_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07547_ _09022_/D vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07478_ _07478_/A _07478_/B _07478_/C vssd1 vssd1 vccd1 vccd1 _07539_/C sky130_fd_sc_hd__nand3_1
X_09217_ _09217_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06429_ _06429_/A _06429_/B vssd1 vssd1 vccd1 vccd1 _06436_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_91_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09148_ _09146_/Y _08634_/B _09147_/Y vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09079_ _09079_/A _09079_/B vssd1 vssd1 vccd1 vccd1 _09087_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06721__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09198__B _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05800__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__D _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10494__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05800_ _09685_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _05805_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06780_ _06782_/A vssd1 vssd1 vccd1 vccd1 _06781_/B sky130_fd_sc_hd__inv_2
X_05731_ _05732_/B _05732_/A vssd1 vssd1 vccd1 vccd1 _05731_/Y sky130_fd_sc_hd__nand2_1
X_08450_ _08673_/B _08471_/C vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__nand2_1
X_05662_ _05662_/A _05662_/B vssd1 vssd1 vccd1 vccd1 _05751_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08381_ _08381_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07401_ _07362_/A _07363_/A _07371_/A vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__o21a_1
X_07332_ _07447_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07332_/Y sky130_fd_sc_hd__nand2_1
X_05593_ _05420_/C _05420_/B _05590_/Y vssd1 vssd1 vccd1 vccd1 _05609_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ _07250_/Y _07477_/B _07262_/Y vssd1 vssd1 vccd1 vccd1 _07467_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09002_ _09003_/B _09003_/A vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__or2_1
XFILLER_0_73_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07194_ _07196_/B _07197_/C _07197_/B vssd1 vssd1 vccd1 vccd1 _07346_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06214_ _06298_/A _06298_/B _06214_/C vssd1 vssd1 vccd1 vccd1 _06302_/B sky130_fd_sc_hd__nand3_1
X_06145_ _06145_/A vssd1 vssd1 vccd1 vccd1 _06146_/C sky130_fd_sc_hd__inv_2
XFILLER_0_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06076_ _06077_/A _06076_/B _06077_/B vssd1 vssd1 vccd1 vccd1 _06084_/C sky130_fd_sc_hd__nand3_1
X_09904_ _09903_/B _09904_/B _09904_/C vssd1 vssd1 vccd1 vccd1 _10168_/B sky130_fd_sc_hd__nand3b_2
X_09835_ _09835_/A _09835_/B _10019_/B vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__nand3_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _09766_/A vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__inv_2
X_06978_ _07097_/B _07096_/A _07096_/B vssd1 vssd1 vccd1 vccd1 _07098_/B sky130_fd_sc_hd__nand3b_1
X_09697_ _09700_/B _09700_/C vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__nand2_1
X_08717_ _08717_/A _08932_/A _08959_/A vssd1 vssd1 vccd1 vccd1 _08721_/C sky130_fd_sc_hd__nand3_1
X_05929_ _05929_/A _05929_/B _05929_/C vssd1 vssd1 vccd1 vccd1 _06328_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08648_ _08415_/Y _08654_/B _08416_/Y vssd1 vssd1 vccd1 vccd1 _09181_/A sky130_fd_sc_hd__a21oi_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08579_ _08579_/A _08579_/B _08579_/C vssd1 vssd1 vccd1 vccd1 _08586_/C sky130_fd_sc_hd__nand3_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10472_ _10494_/CLK _10472_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07547__A _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07266__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__B _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06345__B _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07950_ _07950_/A _07950_/B vssd1 vssd1 vccd1 vccd1 _07951_/B sky130_fd_sc_hd__nand2_1
X_06901_ _09560_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _07064_/B sky130_fd_sc_hd__nand2_1
X_07881_ _07928_/B _07928_/C _07880_/Y vssd1 vssd1 vccd1 vccd1 _07921_/A sky130_fd_sc_hd__a21oi_1
X_09620_ _09626_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09916_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08288__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ _06779_/Y _06849_/B _06788_/Y vssd1 vssd1 vccd1 vccd1 _06841_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10464__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _09716_/B _09551_/B vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__nand2_1
X_06763_ _06862_/B _06861_/A vssd1 vssd1 vccd1 vccd1 _06865_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08502_ _08508_/A _08763_/A vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__nand2_1
X_05714_ _10043_/A input12/X vssd1 vssd1 vccd1 vccd1 _05716_/A sky130_fd_sc_hd__nand2_1
X_09482_ _09482_/A _09799_/A _09482_/C vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06694_ _06698_/B _06695_/A vssd1 vssd1 vccd1 vccd1 _06697_/A sky130_fd_sc_hd__nand2_1
X_05645_ input41/X vssd1 vssd1 vccd1 vccd1 _10026_/A sky130_fd_sc_hd__clkbuf_8
X_08433_ _08445_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__nand2_1
X_08364_ _08368_/B _08368_/C vssd1 vssd1 vccd1 vccd1 _08366_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05576_ _05576_/A _05576_/B vssd1 vssd1 vccd1 vccd1 _05576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07315_ _07315_/A _07315_/B vssd1 vssd1 vccd1 vccd1 _07315_/Y sky130_fd_sc_hd__nor2_1
X_08295_ _08295_/A _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08511_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07246_ _10050_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _07488_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07177_ _07177_/A vssd1 vssd1 vccd1 vccd1 _07180_/B sky130_fd_sc_hd__inv_2
XFILLER_0_5_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06128_ _06128_/A _06128_/B vssd1 vssd1 vccd1 vccd1 _06131_/A sky130_fd_sc_hd__nand2_1
X_06059_ _06063_/A _06063_/C vssd1 vssd1 vccd1 vccd1 _06061_/A sky130_fd_sc_hd__nand2_1
X_09818_ _09963_/A _09962_/B _09962_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09819_/B
+ sky130_fd_sc_hd__a22o_1
X_09749_ input24/X vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__inv_2
XFILLER_0_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05350__A _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 a_i[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput29 a_i[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
X_10455_ _10455_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__nand2_1
X_10386_ _10387_/B _10387_/A vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__or2_1
XANTENNA__05509__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10487__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05525__A _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05430_ _05464_/C vssd1 vssd1 vccd1 vccd1 _05461_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05361_ input7/X _08689_/A vssd1 vssd1 vccd1 vccd1 _05380_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07100_ _09854_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _07104_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05292_ _05908_/B _05292_/B vssd1 vssd1 vccd1 vccd1 _05294_/A sky130_fd_sc_hd__nand2_1
X_08080_ _08080_/A _08176_/C vssd1 vssd1 vccd1 vccd1 _08081_/B sky130_fd_sc_hd__nand2_1
X_07031_ _07031_/A _07031_/B _07031_/C vssd1 vssd1 vccd1 vccd1 _07197_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__D _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08982_ _08982_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07933_ _07932_/B _07933_/B _07933_/C vssd1 vssd1 vccd1 vccd1 _07986_/C sky130_fd_sc_hd__nand3b_1
X_07864_ _07941_/B _07938_/A vssd1 vssd1 vccd1 vccd1 _07866_/A sky130_fd_sc_hd__nand2_1
X_09603_ _09604_/A _09602_/Y vssd1 vssd1 vccd1 vccd1 _09873_/C sky130_fd_sc_hd__or2b_1
X_06815_ _07148_/B _07148_/A vssd1 vssd1 vccd1 vccd1 _06817_/B sky130_fd_sc_hd__nor2_1
X_07795_ _07815_/C _07815_/B _07794_/Y vssd1 vssd1 vccd1 vccd1 _07887_/A sky130_fd_sc_hd__a21oi_2
X_09534_ _09536_/B vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__inv_2
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08746__A _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06746_ _06746_/A _06746_/B vssd1 vssd1 vccd1 vccd1 _06842_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _09465_/A vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__inv_2
XFILLER_0_66_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06677_ _09720_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _06893_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08416_ _08652_/C _08651_/A vssd1 vssd1 vccd1 vccd1 _08416_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05628_ _05979_/A _05628_/B _05628_/C vssd1 vssd1 vccd1 vccd1 _05629_/B sky130_fd_sc_hd__nand3_1
X_09396_ _09396_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _09648_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10028__A1 _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10028__B2 _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08347_ _10026_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _08354_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05559_ _05559_/A _05559_/B vssd1 vssd1 vccd1 vccd1 _05563_/A sky130_fd_sc_hd__nand2_2
X_08278_ _08279_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07229_ _07229_/A _07229_/B _07229_/C vssd1 vssd1 vccd1 vccd1 _07417_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10240_ hold93/X vssd1 vssd1 vccd1 vccd1 _10488_/D sky130_fd_sc_hd__clkbuf_1
X_10171_ _10171_/A _10171_/B vssd1 vssd1 vccd1 vccd1 _10173_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07560__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06904__A _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10507_ _10509_/CLK _10507_/D fanout99/A vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10438_ _10438_/A _10440_/A vssd1 vssd1 vccd1 vccd1 _10439_/A sky130_fd_sc_hd__and2_1
X_10369_ hold63/X hold49/X hold60/X hold57/X vssd1 vssd1 vccd1 vccd1 _10376_/C sky130_fd_sc_hd__and4_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08566__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06600_ _06600_/A _06600_/B _06600_/C vssd1 vssd1 vccd1 vccd1 _06617_/C sky130_fd_sc_hd__nand3_1
X_07580_ _07579_/B _07580_/B _07580_/C vssd1 vssd1 vccd1 vccd1 _07600_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10502__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06531_ _06536_/A _06537_/C vssd1 vssd1 vccd1 vccd1 _06535_/A sky130_fd_sc_hd__nand2_1
X_09250_ _09018_/A _09017_/A _09053_/A vssd1 vssd1 vccd1 vccd1 _09251_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06462_ _06467_/B _06467_/C vssd1 vssd1 vccd1 vccd1 _06468_/A sky130_fd_sc_hd__nand2_1
X_08201_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08202_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09181_ _09181_/A _09181_/B vssd1 vssd1 vccd1 vccd1 _09182_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06393_ _05974_/Y _06392_/Y _06394_/B vssd1 vssd1 vccd1 vccd1 _06643_/C sky130_fd_sc_hd__o21bai_1
X_05413_ _05413_/A _05413_/B vssd1 vssd1 vccd1 vccd1 _05420_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08132_ _08132_/A _08194_/A vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05344_ _05346_/B _05344_/B vssd1 vssd1 vccd1 vccd1 _05345_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05275_ _05554_/A _05554_/B vssd1 vssd1 vccd1 vccd1 _05281_/C sky130_fd_sc_hd__nand2_1
X_08063_ _08065_/B vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07014_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07023_/B sky130_fd_sc_hd__inv_2
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08965_ _09227_/C _08965_/B vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__xor2_1
X_07916_ _07916_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08075_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09282__D _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08896_ _09144_/C vssd1 vssd1 vccd1 vccd1 _09143_/B sky130_fd_sc_hd__inv_2
X_07847_ _07938_/A _07939_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07941_/B sky130_fd_sc_hd__nand3_1
X_07778_ _07849_/B _07849_/A vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__or2_1
X_09517_ _09517_/A _09517_/B vssd1 vssd1 vccd1 vccd1 _09523_/B sky130_fd_sc_hd__nand2_1
X_06729_ _06962_/A _06962_/B _06963_/A vssd1 vssd1 vccd1 vccd1 _06965_/B sky130_fd_sc_hd__nand3_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09448_ _09448_/A _09448_/B vssd1 vssd1 vccd1 vccd1 _09451_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_54_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09379_ _09622_/A _09379_/B _09379_/C vssd1 vssd1 vccd1 vccd1 _09383_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_46_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06443__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ hold72/X _10223_/B vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__nand2_1
X_10154_ _10154_/A _10154_/B _10154_/C vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__nand3_1
X_10085_ input49/X _09720_/B input50/X _09560_/B vssd1 vssd1 vccd1 vccd1 _10086_/B
+ sky130_fd_sc_hd__a22o_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08750_ _08750_/A _08750_/B vssd1 vssd1 vccd1 vccd1 _08751_/B sky130_fd_sc_hd__nand2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05962_ _05962_/A _05962_/B vssd1 vssd1 vccd1 vccd1 _05964_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07184__B _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08681_ _08911_/B _08682_/C _08682_/B vssd1 vssd1 vccd1 vccd1 _08684_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07701_ _07701_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__nand2_1
X_05893_ _05893_/A _05893_/B vssd1 vssd1 vccd1 vccd1 _05895_/A sky130_fd_sc_hd__nand2_1
X_07632_ _07630_/Y _07403_/B _07631_/Y vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ _09302_/A _09303_/A vssd1 vssd1 vccd1 vccd1 _09308_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07563_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07564_/B sky130_fd_sc_hd__nand2_1
X_06514_ _08375_/A _06514_/B vssd1 vssd1 vccd1 vccd1 _06519_/C sky130_fd_sc_hd__nand2_1
X_07494_ _10051_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _07498_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ _09233_/A vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06445_ _06445_/A _06445_/B vssd1 vssd1 vccd1 vccd1 _06449_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _09164_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09169_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08115_ _08116_/B _08116_/A vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__or2_1
X_06376_ _06376_/A _06376_/B vssd1 vssd1 vccd1 vccd1 _06379_/A sky130_fd_sc_hd__nand2_1
X_09095_ _09385_/B _09099_/B vssd1 vssd1 vccd1 vccd1 _09098_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05327_ _05327_/A _05614_/B _05330_/A vssd1 vssd1 vccd1 vccd1 _05614_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09855__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _08172_/B vssd1 vssd1 vccd1 vccd1 _08054_/A sky130_fd_sc_hd__inv_2
X_05258_ _05263_/A _05264_/A vssd1 vssd1 vccd1 vccd1 _05262_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09997_ _09997_/A vssd1 vssd1 vccd1 vccd1 _10008_/A sky130_fd_sc_hd__inv_2
X_08948_ _08946_/Y _08948_/B _08948_/C vssd1 vssd1 vccd1 vccd1 _08949_/B sky130_fd_sc_hd__nand3b_1
X_08879_ _08879_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _08882_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08918__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _10207_/B _10207_/A vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__or2_1
XANTENNA__06901__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__A2 _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ _10137_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__nand2_1
X_10068_ _10071_/B _10071_/C vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09315__A2 _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06348__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06230_ _06353_/A _06354_/A vssd1 vssd1 vccd1 vccd1 _06230_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06161_ _06161_/A _06161_/B vssd1 vssd1 vccd1 vccd1 _06163_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06092_ _06095_/B _06095_/C vssd1 vssd1 vccd1 vccd1 _06094_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09920_ _09920_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09851_ _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09851_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__05708__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A _09782_/B vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__nand2_1
X_08802_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _08802_/Y sky130_fd_sc_hd__nor2_1
X_06994_ _06991_/Y _07680_/C _06993_/Y vssd1 vssd1 vccd1 vccd1 _06997_/A sky130_fd_sc_hd__a21oi_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08733_/A vssd1 vssd1 vccd1 vccd1 _08735_/B sky130_fd_sc_hd__inv_2
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05945_ _06343_/C _06343_/B _05944_/Y vssd1 vssd1 vccd1 vccd1 _06334_/A sky130_fd_sc_hd__a21oi_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08664_/A vssd1 vssd1 vccd1 vccd1 _08665_/B sky130_fd_sc_hd__inv_2
X_05876_ _06219_/A _06219_/B vssd1 vssd1 vccd1 vccd1 _05882_/A sky130_fd_sc_hd__nand2_1
X_08595_ _08601_/B _08601_/C vssd1 vssd1 vccd1 vccd1 _09147_/B sky130_fd_sc_hd__nand2_1
X_07615_ _07523_/B _07523_/C _07524_/B vssd1 vssd1 vccd1 vccd1 _07616_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_76_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07546_ _07717_/B _07717_/C vssd1 vssd1 vccd1 vccd1 _07719_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09216_ _09216_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09243_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07477_ _07477_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07539_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06428_ _08214_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _06429_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09147_ _09147_/A _09147_/B vssd1 vssd1 vccd1 vccd1 _09147_/Y sky130_fd_sc_hd__nor2_1
X_06359_ _06359_/A _06359_/B vssd1 vssd1 vccd1 vccd1 _06751_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_16_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09078_ _09079_/B _09079_/A vssd1 vssd1 vccd1 vccd1 _09087_/A sky130_fd_sc_hd__or2_1
X_08029_ _08029_/A _08030_/B _08030_/A vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_31_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08668__A_N _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05800__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09942__B _10171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05730_ _06176_/A _05736_/C vssd1 vssd1 vccd1 vccd1 _06186_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05661_ _05661_/A _05661_/B vssd1 vssd1 vccd1 vccd1 _05751_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08380_ _06544_/A _06543_/A _06583_/A vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07400_ _07400_/A _07400_/B vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07331_ _07327_/Y _07329_/Y _07458_/A vssd1 vssd1 vccd1 vccd1 _07448_/B sky130_fd_sc_hd__a21oi_2
X_05592_ _05609_/A _05610_/B vssd1 vssd1 vccd1 vccd1 _05608_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07262_ _07475_/C _07474_/A vssd1 vssd1 vccd1 vccd1 _07262_/Y sky130_fd_sc_hd__nor2_1
X_09001_ _09234_/A _09000_/Y vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__nor2b_1
X_07193_ _07181_/C _07181_/B _07040_/Y vssd1 vssd1 vccd1 vccd1 _07196_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06213_ _06216_/B _06213_/B vssd1 vssd1 vccd1 vccd1 _06217_/B sky130_fd_sc_hd__nand2b_1
X_06144_ _06144_/A _06145_/A vssd1 vssd1 vccd1 vccd1 _06151_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06075_ _06484_/A _06484_/B vssd1 vssd1 vccd1 vccd1 _06077_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _09903_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09905_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09527__A2 _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ _09834_/A vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__inv_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09765_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__xor2_1
X_06977_ _06977_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _07096_/B sky130_fd_sc_hd__nand2_1
X_09696_ _10034_/A _10039_/B _09696_/C vssd1 vssd1 vccd1 vccd1 _09700_/C sky130_fd_sc_hd__nand3_1
X_08716_ _08716_/A vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__inv_2
X_05928_ _05928_/A _05928_/B _05928_/C vssd1 vssd1 vccd1 vccd1 _05929_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08647_ _08647_/A _08647_/B vssd1 vssd1 vccd1 vccd1 _09181_/B sky130_fd_sc_hd__nand2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05859_ _08272_/B vssd1 vssd1 vccd1 vccd1 _09485_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _08578_/A _08578_/B vssd1 vssd1 vccd1 vccd1 _08586_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07529_ _07529_/A _07529_/B vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10471_ _10495_/CLK _10471_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__07828__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09953__A _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06900_ _06911_/B _06911_/C vssd1 vssd1 vccd1 vccd1 _06910_/A sky130_fd_sc_hd__nand2_1
X_07880_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07880_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08288__B _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ _06831_/A _06831_/B _06831_/C vssd1 vssd1 vccd1 vccd1 _06839_/A sky130_fd_sc_hd__nand3_1
X_09550_ _09199_/A _10043_/B _09548_/A _10052_/A vssd1 vssd1 vccd1 vccd1 _09551_/B
+ sky130_fd_sc_hd__a22o_1
X_06762_ _10026_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _06861_/A sky130_fd_sc_hd__nand2_1
X_09481_ _09481_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09518_/B sky130_fd_sc_hd__nand2_1
X_08501_ _08500_/B _08501_/B _08763_/B vssd1 vssd1 vccd1 vccd1 _08763_/A sky130_fd_sc_hd__nand3b_1
X_05713_ _05717_/A _05717_/B vssd1 vssd1 vccd1 vccd1 _05715_/A sky130_fd_sc_hd__nand2_1
X_08432_ _08431_/B _08674_/A _08432_/C vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_53_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06693_ _06696_/B vssd1 vssd1 vccd1 vccd1 _06698_/B sky130_fd_sc_hd__inv_2
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05644_ _05683_/B _05650_/C vssd1 vssd1 vccd1 vccd1 _05648_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ _08362_/B _08363_/B _08363_/C vssd1 vssd1 vccd1 vccd1 _08368_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_58_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05575_ _05627_/B _05628_/B _05628_/C vssd1 vssd1 vccd1 vccd1 _05626_/A sky130_fd_sc_hd__nand3_1
X_08294_ _08294_/A _08532_/A vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07314_ _07319_/B _07319_/C vssd1 vssd1 vccd1 vccd1 _07377_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07245_ _07248_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _07489_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06552__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _07180_/A _07177_/A vssd1 vssd1 vccd1 vccd1 _07179_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06127_ _06127_/A _06127_/B _06130_/A vssd1 vssd1 vccd1 vccd1 _06134_/A sky130_fd_sc_hd__nand3_1
X_06058_ _06058_/A _06058_/B vssd1 vssd1 vccd1 vccd1 _06063_/C sky130_fd_sc_hd__nand2_1
X_09817_ _09963_/A _09962_/A _09962_/B _09960_/B vssd1 vssd1 vccd1 vccd1 _09817_/X
+ sky130_fd_sc_hd__and4_1
X_09748_ _09986_/A input21/X vssd1 vssd1 vccd1 vccd1 _09754_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _10455_/B vssd1 vssd1 vccd1 vccd1 _09679_/Y sky130_fd_sc_hd__inv_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05350__B _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 a_i[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_2
X_10454_ _10454_/A vssd1 vssd1 vccd1 vccd1 _10476_/D sky130_fd_sc_hd__buf_1
X_10385_ _10385_/A _10385_/B _10385_/C vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__or3_1
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05360_ _05380_/A vssd1 vssd1 vccd1 vccd1 _05362_/A sky130_fd_sc_hd__inv_2
XFILLER_0_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05291_ _05292_/B _05291_/B _05291_/C vssd1 vssd1 vccd1 vccd1 _05908_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07030_ _07032_/B _07030_/B vssd1 vssd1 vccd1 vccd1 _07031_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08981_ _08981_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07932_ _07932_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _07986_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09363__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ _07936_/C _07936_/B vssd1 vssd1 vccd1 vccd1 _07922_/C sky130_fd_sc_hd__nand2_1
X_09602_ _09604_/B vssd1 vssd1 vccd1 vccd1 _09602_/Y sky130_fd_sc_hd__inv_2
X_06814_ _07147_/B _07147_/C vssd1 vssd1 vccd1 vccd1 _07148_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09533_ _10026_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _09536_/B sky130_fd_sc_hd__nand2_1
X_07794_ _07816_/A _07817_/A vssd1 vssd1 vccd1 vccd1 _07794_/Y sky130_fd_sc_hd__nor2_1
X_06745_ _06747_/A _06747_/B vssd1 vssd1 vccd1 vccd1 _06746_/A sky130_fd_sc_hd__nand2_1
X_09464_ _09981_/A _09981_/B input18/X input19/X vssd1 vssd1 vccd1 vccd1 _09465_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__06547__A _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06676_ _06891_/A _06892_/A vssd1 vssd1 vccd1 vccd1 _06681_/B sky130_fd_sc_hd__nand2_1
X_09395_ _09397_/C vssd1 vssd1 vccd1 vccd1 _09396_/B sky130_fd_sc_hd__inv_2
X_08415_ _08651_/A _08652_/C vssd1 vssd1 vccd1 vccd1 _08415_/Y sky130_fd_sc_hd__nand2_1
X_05627_ _05979_/B _05627_/B vssd1 vssd1 vccd1 vccd1 _05629_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10028__A2 _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08346_ _08346_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05558_ _05561_/B _06043_/A _05562_/A vssd1 vssd1 vccd1 vccd1 _05560_/B sky130_fd_sc_hd__nand3_1
X_08277_ _08279_/B vssd1 vssd1 vccd1 vccd1 _08278_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05489_ _05489_/A _05490_/B _05489_/C vssd1 vssd1 vccd1 vccd1 _05960_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_6_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07228_ _07228_/A _07228_/B vssd1 vssd1 vccd1 vccd1 _07229_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06282__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ _07713_/A _07159_/B vssd1 vssd1 vccd1 vccd1 _07162_/A sky130_fd_sc_hd__nand2_1
X_10170_ _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _10171_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08937__A _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07560__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10506_ _10509_/CLK _10506_/D fanout99/A vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06904__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10437_ _10437_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _10440_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10368_ hold69/X _10368_/B vssd1 vssd1 vccd1 vccd1 _10368_/Y sky130_fd_sc_hd__nor2_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06920__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10298_/Y _10299_/B _10299_/C vssd1 vssd1 vccd1 vccd1 _10299_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07751__A _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08566__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06530_ _06063_/C _06063_/B _06057_/A vssd1 vssd1 vccd1 vccd1 _06537_/C sky130_fd_sc_hd__a21oi_2
X_06461_ _06469_/C vssd1 vssd1 vccd1 vccd1 _06466_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05412_ _05590_/B vssd1 vssd1 vccd1 vccd1 _05413_/B sky130_fd_sc_hd__inv_2
X_08200_ _08200_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08201_/B sky130_fd_sc_hd__nand2_1
X_09180_ _09180_/A _09180_/B vssd1 vssd1 vccd1 vccd1 _09183_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06392_ _06394_/C vssd1 vssd1 vccd1 vccd1 _06392_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ _08169_/B _08175_/A vssd1 vssd1 vccd1 vccd1 _08168_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05343_ _05343_/A vssd1 vssd1 vccd1 vccd1 _05346_/B sky130_fd_sc_hd__inv_2
X_05274_ _05274_/A _05274_/B vssd1 vssd1 vccd1 vccd1 _05281_/A sky130_fd_sc_hd__nand2_1
X_08062_ _08176_/C _08080_/A vssd1 vssd1 vccd1 vccd1 _08062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07013_ _07013_/A _07013_/B _07013_/C vssd1 vssd1 vccd1 vccd1 _07021_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08964_ _09963_/A _09496_/B vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__nand2_1
X_07915_ _07918_/A _08206_/B vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__nand2_1
X_08895_ _08895_/A _09132_/A vssd1 vssd1 vccd1 vccd1 _09144_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07846_ _07846_/A _07846_/B _07846_/C vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__nand3_1
X_07777_ _07779_/B _07777_/B vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__nand2_1
X_09516_ _09516_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09517_/B sky130_fd_sc_hd__nand2_1
X_06728_ _06982_/B _06982_/A vssd1 vssd1 vccd1 vccd1 _06963_/A sky130_fd_sc_hd__nor2_1
X_09447_ _09447_/A vssd1 vssd1 vccd1 vccd1 _09448_/B sky130_fd_sc_hd__inv_2
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10477__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06659_ _06791_/B _06791_/C vssd1 vssd1 vccd1 vccd1 _06793_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ _09378_/A _09378_/B vssd1 vssd1 vccd1 vccd1 _09622_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08492__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08330_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10222_ _10223_/B hold72/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__or2_1
X_10153_ _10153_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10084_ _10084_/A _10084_/B _10084_/C _10084_/D vssd1 vssd1 vccd1 vccd1 _10086_/A
+ sky130_fd_sc_hd__or4_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06618__C _06618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10488__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10437__A _10437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07746__A _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _07700_/A _07700_/B _07700_/C vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__nand3_1
X_05961_ _05963_/B _05963_/C vssd1 vssd1 vccd1 vccd1 _05962_/A sky130_fd_sc_hd__nand2_1
X_08680_ _08680_/A vssd1 vssd1 vccd1 vccd1 _08682_/B sky130_fd_sc_hd__inv_2
X_05892_ _05894_/A _05893_/A _05893_/B vssd1 vssd1 vccd1 vccd1 _05897_/B sky130_fd_sc_hd__nand3_1
X_07631_ _07631_/A _07631_/B vssd1 vssd1 vccd1 vccd1 _07631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07562_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07562_/Y sky130_fd_sc_hd__nor2_1
X_09301_ _09301_/A _09301_/B vssd1 vssd1 vccd1 vccd1 _09303_/A sky130_fd_sc_hd__nand2_1
X_06513_ _06512_/B _06513_/B _06513_/C vssd1 vssd1 vccd1 vccd1 _06514_/B sky130_fd_sc_hd__nand3b_1
X_07493_ _10050_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _07497_/A sky130_fd_sc_hd__nand2_1
X_09232_ _09236_/B _09542_/B vssd1 vssd1 vccd1 vccd1 _09235_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06444_ _06445_/A _06445_/B vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09163_ _09172_/A _09172_/B _09171_/C vssd1 vssd1 vccd1 vccd1 _09164_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06375_ _06377_/A vssd1 vssd1 vccd1 vccd1 _06376_/B sky130_fd_sc_hd__inv_2
XFILLER_0_28_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08114_ _08020_/Y _08114_/B vssd1 vssd1 vccd1 vccd1 _08116_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05326_ _05397_/C _05376_/A vssd1 vssd1 vccd1 vccd1 _05330_/A sky130_fd_sc_hd__nand2_1
X_09094_ _09094_/A _09094_/B vssd1 vssd1 vccd1 vccd1 _09099_/B sky130_fd_sc_hd__nand2_1
X_08045_ _08087_/A _08087_/B _08045_/C vssd1 vssd1 vccd1 vccd1 _08172_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05257_ _05503_/B vssd1 vssd1 vccd1 vccd1 _05264_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09996_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__nand2_1
X_08947_ _08947_/A _08947_/B vssd1 vssd1 vccd1 vccd1 _08948_/C sky130_fd_sc_hd__nand2_1
X_08878_ _08879_/B _08879_/A vssd1 vssd1 vccd1 vccd1 _08878_/Y sky130_fd_sc_hd__nor2_1
X_07829_ _09560_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _07833_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10510__RESET_B fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10205_ hold86/A _10193_/B _10200_/A hold96/X vssd1 vssd1 vccd1 vccd1 _10207_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10136_ _10138_/C vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__inv_2
X_10067_ _10067_/A _10067_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10071_/C sky130_fd_sc_hd__nand3_1
Xclkbuf_2_3__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10509_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06645__A _06820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06160_ _06162_/C vssd1 vssd1 vccd1 vccd1 _06161_/B sky130_fd_sc_hd__inv_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06091_ _06579_/A _06511_/A _06091_/C vssd1 vssd1 vccd1 vccd1 _06095_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_40_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09850_ _09851_/B _09851_/A vssd1 vssd1 vccd1 vccd1 _09850_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05708__B _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09782_/B _09782_/A vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__or2_1
X_08801_ _08802_/B _08802_/A vssd1 vssd1 vccd1 vccd1 _08801_/Y sky130_fd_sc_hd__nand2_1
X_06993_ _07138_/A _07137_/A vssd1 vssd1 vccd1 vccd1 _06993_/Y sky130_fd_sc_hd__nor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _09951_/A _09496_/B vssd1 vssd1 vccd1 vccd1 _08733_/A sky130_fd_sc_hd__nand2_1
X_05944_ _06340_/B _06339_/A vssd1 vssd1 vccd1 vccd1 _05944_/Y sky130_fd_sc_hd__nor2_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__B1 _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _08663_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08665_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05875_ _05875_/A _05875_/B _05875_/C vssd1 vssd1 vccd1 vccd1 _06219_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08594_ _08594_/A _08594_/B _08594_/C vssd1 vssd1 vccd1 vccd1 _08601_/C sky130_fd_sc_hd__nand3_2
X_07614_ _07614_/A _07614_/B vssd1 vssd1 vccd1 vccd1 _07616_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07545_ _07545_/A _07545_/B _07545_/C vssd1 vssd1 vccd1 vccd1 _07717_/C sky130_fd_sc_hd__nand3_1
XANTENNA__10085__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07476_ _07478_/A _07478_/B vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__nand2_1
X_09215_ _09215_/A _09215_/B _09215_/C vssd1 vssd1 vccd1 vccd1 _09216_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06427_ _08225_/B _06430_/C vssd1 vssd1 vccd1 vccd1 _06429_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09146_ _09147_/B _09147_/A vssd1 vssd1 vccd1 vccd1 _09146_/Y sky130_fd_sc_hd__nand2_1
X_06358_ _06358_/A _06358_/B _06358_/C vssd1 vssd1 vccd1 vccd1 _06359_/B sky130_fd_sc_hd__nand3_1
X_09077_ _09077_/A _09076_/Y vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__nor2b_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05309_ _05308_/B _05559_/B _05309_/C vssd1 vssd1 vccd1 vccd1 _05559_/A sky130_fd_sc_hd__nand3b_2
X_06289_ _06707_/C _06707_/B _06288_/Y vssd1 vssd1 vccd1 vccd1 _06296_/A sky130_fd_sc_hd__a21o_1
X_08028_ _08028_/A _08028_/B vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _10016_/A vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__inv_2
XANTENNA__09106__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09776__A _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10119_ _10120_/B _10120_/A vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05660_ _05662_/B vssd1 vssd1 vccd1 vccd1 _05661_/B sky130_fd_sc_hd__inv_2
X_05591_ _05420_/C _05420_/B _05590_/Y vssd1 vssd1 vccd1 vccd1 _05610_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ _07330_/A _07330_/B vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_73_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ _10027_/A _10044_/D _08999_/C vssd1 vssd1 vccd1 vccd1 _09000_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07261_ _07478_/C vssd1 vssd1 vccd1 vccd1 _07477_/B sky130_fd_sc_hd__inv_2
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09686__A _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ _07234_/B _07234_/C _07191_/Y vssd1 vssd1 vccd1 vccd1 _07227_/A sky130_fd_sc_hd__a21oi_2
X_06212_ _06810_/B _06810_/C vssd1 vssd1 vccd1 vccd1 _06809_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06143_ _10043_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _06145_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06074_ _06078_/B vssd1 vssd1 vccd1 vccd1 _06076_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _09904_/B _09904_/C vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09527__A3 _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09833_ _09833_/A _09834_/A vssd1 vssd1 vccd1 vccd1 _09840_/A sky130_fd_sc_hd__nand2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09762_/Y _09764_/B vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__and2b_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06976_ _06976_/A _06976_/B vssd1 vssd1 vccd1 vccd1 _07096_/A sky130_fd_sc_hd__nand2_1
X_09695_ _10039_/A _09695_/B vssd1 vssd1 vccd1 vccd1 _09700_/B sky130_fd_sc_hd__nand2_1
X_08715_ _08959_/B _08716_/A vssd1 vssd1 vccd1 vccd1 _08721_/B sky130_fd_sc_hd__nand2_1
X_05927_ _05927_/A _05927_/B vssd1 vssd1 vccd1 vccd1 _05929_/A sky130_fd_sc_hd__nand2_1
X_08646_ _08646_/A _08647_/A _08647_/B vssd1 vssd1 vccd1 vccd1 _09180_/B sky130_fd_sc_hd__nand3_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05858_ _09022_/D vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08577_ _08579_/C vssd1 vssd1 vccd1 vccd1 _08578_/B sky130_fd_sc_hd__inv_2
X_05789_ input37/X vssd1 vssd1 vccd1 vccd1 _09962_/A sky130_fd_sc_hd__clkbuf_8
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ _07528_/A _07528_/B vssd1 vssd1 vccd1 vccd1 _07529_/B sky130_fd_sc_hd__nand2_1
X_07459_ _07459_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07598_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470_ _10494_/CLK _10470_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfrtp_1
X_09129_ _09136_/B _09414_/A vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07828__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08005__A _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08675__A _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06830_ _07146_/B _07146_/C vssd1 vssd1 vccd1 vccd1 _06996_/A sky130_fd_sc_hd__nand2_1
X_06761_ _09684_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _06862_/B sky130_fd_sc_hd__nand2_1
X_09480_ _09482_/A vssd1 vssd1 vccd1 vccd1 _09481_/B sky130_fd_sc_hd__inv_2
X_08500_ _08500_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08508_/A sky130_fd_sc_hd__nand2_1
X_05712_ _05712_/A _05712_/B vssd1 vssd1 vccd1 vccd1 _05717_/B sky130_fd_sc_hd__nand2_1
X_06692_ _06930_/C _06930_/B _06691_/Y vssd1 vssd1 vccd1 vccd1 _06703_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08431_ _08431_/A _08431_/B vssd1 vssd1 vccd1 vccd1 _08445_/A sky130_fd_sc_hd__nand2_1
X_05643_ _05643_/A _05643_/B vssd1 vssd1 vccd1 vccd1 _05650_/C sky130_fd_sc_hd__nand2_1
X_08362_ _08362_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08368_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05574_ _05574_/A _05574_/B _05574_/C vssd1 vssd1 vccd1 vccd1 _05628_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08293_ _08532_/A _08294_/A vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__or2_1
X_07313_ _07313_/A _07313_/B _07313_/C vssd1 vssd1 vccd1 vccd1 _07319_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07244_ _10052_/A _08422_/A vssd1 vssd1 vccd1 vccd1 _07248_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06552__B _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ _07178_/B vssd1 vssd1 vccd1 vccd1 _07180_/A sky130_fd_sc_hd__inv_2
X_06126_ _06126_/A _06126_/B vssd1 vssd1 vccd1 vccd1 _06130_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06057_ _06057_/A vssd1 vssd1 vccd1 vccd1 _06063_/A sky130_fd_sc_hd__inv_2
XANTENNA__08479__B _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _09960_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__nand2_1
X_09747_ _09843_/B vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__inv_2
X_06959_ _06959_/A _06959_/B vssd1 vssd1 vccd1 vccd1 _06959_/Y sky130_fd_sc_hd__nor2_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _10452_/A _09678_/B vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08495__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08629_ _09150_/B _08631_/C vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07839__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10453_ _10453_/A _10455_/A vssd1 vssd1 vccd1 vccd1 _10454_/A sky130_fd_sc_hd__and2_1
XFILLER_0_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10384_ _08179_/A _10384_/B _10384_/C vssd1 vssd1 vccd1 vccd1 _10385_/C sky130_fd_sc_hd__nand3b_1
XANTENNA__05359__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08389__B _08390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06918__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05290_ _05337_/B _05338_/C _05338_/B vssd1 vssd1 vccd1 vccd1 _05292_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10175__A _10175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _08982_/B _08981_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09337_/A sky130_fd_sc_hd__nand3b_1
X_07931_ _07933_/B _07933_/C vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09363__B2 _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _07862_/A _07970_/A _07862_/C vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__nand3_1
X_09601_ input51/X _09601_/B vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__nand2_1
X_06813_ _06812_/B _06813_/B _06813_/C vssd1 vssd1 vccd1 vccd1 _07147_/C sky130_fd_sc_hd__nand3b_2
X_09532_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__inv_2
X_07793_ _07889_/B _07818_/B vssd1 vssd1 vccd1 vccd1 _07815_/B sky130_fd_sc_hd__nor2b_1
X_06744_ _06744_/A _06744_/B vssd1 vssd1 vccd1 vccd1 _06747_/B sky130_fd_sc_hd__nand2_1
X_09463_ _09980_/A input17/X vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06547__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ _06891_/B vssd1 vssd1 vccd1 vccd1 _06892_/A sky130_fd_sc_hd__inv_2
X_09394_ _09634_/B _09394_/B vssd1 vssd1 vccd1 vccd1 _09397_/C sky130_fd_sc_hd__nand2_1
X_08414_ _08651_/B vssd1 vssd1 vccd1 vccd1 _08652_/C sky130_fd_sc_hd__inv_2
X_05626_ _05626_/A _05626_/B _05626_/C vssd1 vssd1 vccd1 vccd1 _05631_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08345_ _08331_/Y _08345_/B _08345_/C vssd1 vssd1 vccd1 vccd1 _08346_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05557_ _05281_/C _05281_/B _05554_/Y vssd1 vssd1 vccd1 vccd1 _05561_/B sky130_fd_sc_hd__a21o_1
X_08276_ _09951_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _08279_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05488_ _05827_/B vssd1 vssd1 vccd1 vccd1 _05489_/C sky130_fd_sc_hd__inv_2
XFILLER_0_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07227_ _07227_/A vssd1 vssd1 vccd1 vccd1 _07228_/A sky130_fd_sc_hd__inv_2
XANTENNA__06282__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07158_ _10428_/A _07156_/Y _10429_/B vssd1 vssd1 vccd1 vccd1 _07159_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06109_ _09685_/A _08814_/B vssd1 vssd1 vccd1 vccd1 _06114_/A sky130_fd_sc_hd__nand2_1
X_07089_ _07078_/B _07081_/A _07088_/Y vssd1 vssd1 vccd1 vccd1 _07091_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08937__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05361__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10505_ _10511_/CLK hold51/X fanout99/A vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10436_ _10437_/B _10437_/A vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10367_ hold59/X vssd1 vssd1 vccd1 vccd1 _10507_/D sky130_fd_sc_hd__clkbuf_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06920__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10298_/A _10298_/B vssd1 vssd1 vccd1 vccd1 _10298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07751__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06460_ _06460_/A _06460_/B vssd1 vssd1 vccd1 vccd1 _06469_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05411_ input3/X _08272_/B vssd1 vssd1 vccd1 vccd1 _05590_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ _08130_/A _08172_/B _08130_/C vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06391_ _06388_/Y _06812_/B _06390_/Y vssd1 vssd1 vccd1 vccd1 _06816_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05342_ _05346_/A _05343_/A vssd1 vssd1 vccd1 vccd1 _05345_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05273_ _05554_/B vssd1 vssd1 vccd1 vccd1 _05274_/B sky130_fd_sc_hd__inv_2
X_08061_ _08079_/C _08079_/B vssd1 vssd1 vccd1 vccd1 _08080_/A sky130_fd_sc_hd__nand2_1
X_07012_ _07623_/B _07623_/C vssd1 vssd1 vccd1 vccd1 _07625_/A sky130_fd_sc_hd__nand2_1
X_08963_ _09962_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _09227_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07914_ _07914_/A _07914_/B vssd1 vssd1 vccd1 vccd1 _07918_/A sky130_fd_sc_hd__nand2_1
X_08894_ _09132_/B _08894_/B _08894_/C vssd1 vssd1 vccd1 vccd1 _09132_/A sky130_fd_sc_hd__nand3_1
X_07845_ _07845_/A _07845_/B vssd1 vssd1 vccd1 vccd1 _07939_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06558__A input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ _07776_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07777_/B sky130_fd_sc_hd__nand2_1
X_09515_ _09514_/B _09515_/B _09515_/C vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__nand3b_1
X_06727_ _06938_/B _06936_/A vssd1 vssd1 vccd1 vccd1 _06982_/A sky130_fd_sc_hd__and2_1
X_09446_ _09802_/B _09446_/B vssd1 vssd1 vccd1 vccd1 _09451_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06658_ _06658_/A _06658_/B _06658_/C vssd1 vssd1 vccd1 vccd1 _06791_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ _09378_/A _09378_/B _09622_/B vssd1 vssd1 vccd1 vccd1 _09383_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08492__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06589_ _06589_/A _06589_/B vssd1 vssd1 vccd1 vccd1 _06591_/A sky130_fd_sc_hd__nand2_1
X_05609_ _05609_/A _05609_/B vssd1 vssd1 vccd1 vccd1 _05611_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06293__A _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ _08328_/A vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__inv_2
XFILLER_0_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ _08262_/B _08262_/C vssd1 vssd1 vccd1 vccd1 _08261_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10221_ _10221_/A hold71/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10152_ _10154_/A vssd1 vssd1 vccd1 vccd1 _10153_/B sky130_fd_sc_hd__inv_2
XANTENNA__08013__A _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05637__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10083_ input51/X _10083_/B vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__nand2_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08667__B _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07746__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _10407_/B _08210_/C _07714_/A vssd1 vssd1 vccd1 vccd1 _10427_/A sky130_fd_sc_hd__a21bo_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05960_ _05960_/A _05960_/B _05960_/C vssd1 vssd1 vccd1 vccd1 _05963_/C sky130_fd_sc_hd__nand3_1
X_05891_ _05891_/A _05891_/B _05891_/C vssd1 vssd1 vccd1 vccd1 _05893_/B sky130_fd_sc_hd__nand3_1
X_07630_ _07631_/B _07631_/A vssd1 vssd1 vccd1 vccd1 _07630_/Y sky130_fd_sc_hd__nand2_1
X_07561_ _09560_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _07563_/B sky130_fd_sc_hd__nand2_1
X_09300_ _09300_/A _09506_/A _09300_/C vssd1 vssd1 vccd1 vccd1 _09301_/B sky130_fd_sc_hd__nand3_1
X_06512_ _06512_/A _06512_/B vssd1 vssd1 vccd1 vccd1 _08375_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07492_ _09720_/B _09986_/A vssd1 vssd1 vccd1 vccd1 _07556_/C sky130_fd_sc_hd__nand2_1
X_09231_ _09525_/A _09231_/B _09231_/C vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06443_ _09960_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _06445_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09162_ _09162_/A _09162_/B _09162_/C vssd1 vssd1 vccd1 vccd1 _09172_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_61_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06374_ _06735_/A _06736_/A vssd1 vssd1 vccd1 vccd1 _06649_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08113_ _08158_/C _08158_/B _08112_/Y vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05325_ _05376_/A _05325_/B _05376_/B vssd1 vssd1 vccd1 vccd1 _05397_/C sky130_fd_sc_hd__nand3_2
X_09093_ _08832_/C _08832_/B _08819_/A vssd1 vssd1 vccd1 vccd1 _09094_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08044_ _08127_/B _08123_/A vssd1 vssd1 vccd1 vccd1 _08045_/C sky130_fd_sc_hd__nor2_1
X_05256_ _09951_/B _08422_/A vssd1 vssd1 vccd1 vccd1 _05503_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09995_ _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _10010_/C sky130_fd_sc_hd__nand2_1
X_08946_ _08947_/B _08947_/A vssd1 vssd1 vccd1 vccd1 _08946_/Y sky130_fd_sc_hd__nor2_1
X_08877_ _08877_/A _09096_/A vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07828_ _10083_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _07833_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07759_ _07812_/B vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09429_ _09429_/A _09430_/A vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05367__A _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ hold18/X _10196_/Y hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10135_ _10133_/Y _09744_/B _10134_/Y vssd1 vssd1 vccd1 vccd1 _10138_/C sky130_fd_sc_hd__a21oi_2
X_10066_ _10066_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10071_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07582__A _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06645__B _06820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06090_ _06579_/B _06090_/B vssd1 vssd1 vccd1 vccd1 _06095_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05277__A _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08800_/A _08800_/B vssd1 vssd1 vccd1 vccd1 _08802_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09996_/B _09780_/B vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__nand2_1
X_06992_ _06992_/A _06992_/B vssd1 vssd1 vccd1 vccd1 _07680_/C sky130_fd_sc_hd__nand2_2
XANTENNA__10467__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08729_/A _09953_/A _08729_/C vssd1 vssd1 vccd1 vccd1 _08735_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__07492__A _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05943_ _06341_/C vssd1 vssd1 vccd1 vccd1 _06343_/B sky130_fd_sc_hd__inv_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__A1 _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__B2 _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ _08662_/A vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__inv_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05874_ _05874_/A _05874_/B vssd1 vssd1 vccd1 vccd1 _06219_/A sky130_fd_sc_hd__nand2_1
X_07613_ _07899_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _07617_/B sky130_fd_sc_hd__nor2_1
X_08593_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08601_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07544_ _07544_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07717_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10085__B2 _09560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07475_ _07475_/A _07475_/B _07475_/C vssd1 vssd1 vccd1 vccd1 _07478_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_91_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09214_ _09215_/A _09215_/C _09215_/B vssd1 vssd1 vccd1 vccd1 _09216_/A sky130_fd_sc_hd__a21o_1
X_06426_ _06426_/A _06426_/B vssd1 vssd1 vccd1 vccd1 _06430_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09145_ _09162_/B _09162_/C vssd1 vssd1 vccd1 vccd1 _09161_/A sky130_fd_sc_hd__nand2_1
X_06357_ _06357_/A _06357_/B vssd1 vssd1 vccd1 vccd1 _06359_/A sky130_fd_sc_hd__nand2_1
X_09076_ _10084_/A _10113_/D _09075_/C vssd1 vssd1 vccd1 vccd1 _09076_/Y sky130_fd_sc_hd__o21ai_1
X_05308_ _05308_/A _05308_/B vssd1 vssd1 vccd1 vccd1 _05329_/A sky130_fd_sc_hd__nand2_1
X_06288_ _06288_/A _06288_/B vssd1 vssd1 vccd1 vccd1 _06288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08028_/A sky130_fd_sc_hd__nand2_1
X_05239_ input6/X vssd1 vssd1 vccd1 vccd1 _10026_/B sky130_fd_sc_hd__buf_8
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ _09978_/A _09978_/B vssd1 vssd1 vccd1 vccd1 _10016_/A sky130_fd_sc_hd__nand2_1
X_08929_ _08929_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09106__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09466__B1 _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08961__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10118_ _10118_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05544__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10049_ _10049_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05590_ _05590_/A _05590_/B vssd1 vssd1 vccd1 vccd1 _05590_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10472__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07260_ _07260_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _07478_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07191_ _07235_/B _07236_/A vssd1 vssd1 vccd1 vccd1 _07191_/Y sky130_fd_sc_hd__nor2_1
X_06211_ _05969_/Y _06211_/B _06211_/C vssd1 vssd1 vccd1 vccd1 _06810_/C sky130_fd_sc_hd__nand3b_1
X_06142_ _06146_/A _06146_/B vssd1 vssd1 vccd1 vccd1 _06144_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06073_ _09951_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _06078_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _10110_/B _10110_/A vssd1 vssd1 vccd1 vccd1 _09904_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09832_ _09832_/A _09832_/B vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__nand2_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09763_ _09762_/A _09762_/B _09762_/C vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__o21ai_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08716_/A sky130_fd_sc_hd__nand2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06975_ _06977_/B vssd1 vssd1 vccd1 vccd1 _06976_/B sky130_fd_sc_hd__inv_2
X_09694_ _10039_/B vssd1 vssd1 vccd1 vccd1 _09695_/B sky130_fd_sc_hd__inv_2
X_05926_ _06331_/C vssd1 vssd1 vccd1 vccd1 _06330_/B sky130_fd_sc_hd__inv_2
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08645_ _08644_/B _08645_/B _08645_/C vssd1 vssd1 vccd1 vccd1 _08647_/B sky130_fd_sc_hd__nand3b_1
X_05857_ _09720_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _06257_/B sky130_fd_sc_hd__nand2_2
X_08576_ _08576_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _08579_/C sky130_fd_sc_hd__nand2_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07527_ _07527_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07529_/A sky130_fd_sc_hd__nand2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05788_ _05809_/B _05809_/C vssd1 vssd1 vccd1 vccd1 _05798_/A sky130_fd_sc_hd__nand2_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08781__A _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07458_ _07458_/A _07327_/Y vssd1 vssd1 vccd1 vccd1 _07459_/B sky130_fd_sc_hd__nor2b_1
X_06409_ _09963_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _06413_/A sky130_fd_sc_hd__nand2_1
X_07389_ _07391_/B _07392_/B _07392_/C vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__nand3_1
X_09128_ _09135_/B _09414_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_44_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09059_ _09059_/A _09059_/B vssd1 vssd1 vccd1 vccd1 _09400_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08005__B _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09687__B1 _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07100__A _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput90 hold3/A vssd1 vssd1 vccd1 vccd1 y_o[31] sky130_fd_sc_hd__buf_12
XFILLER_0_37_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08866__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ _06854_/B _06854_/C vssd1 vssd1 vccd1 vccd1 _06853_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10505__CLK _10511_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05711_ _05711_/A vssd1 vssd1 vccd1 vccd1 _05717_/A sky130_fd_sc_hd__inv_2
X_06691_ _06926_/A _06927_/B vssd1 vssd1 vccd1 vccd1 _06691_/Y sky130_fd_sc_hd__nor2_1
X_08430_ _08220_/A _08223_/B _08221_/A vssd1 vssd1 vccd1 vccd1 _08431_/B sky130_fd_sc_hd__a21oi_1
X_05642_ _05642_/A _05642_/B vssd1 vssd1 vccd1 vccd1 _05683_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08361_ _08361_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _08362_/B sky130_fd_sc_hd__nand2_1
X_05573_ _05981_/B _05573_/B vssd1 vssd1 vccd1 vccd1 _05574_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08292_ _08292_/A _08292_/B vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07312_ _07312_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07319_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07243_ _10051_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07174_ _07237_/B vssd1 vssd1 vccd1 vccd1 _07234_/B sky130_fd_sc_hd__inv_2
X_06125_ _06128_/B _06534_/A _06129_/A vssd1 vssd1 vccd1 vccd1 _06127_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06056_ _06058_/A _06058_/B vssd1 vssd1 vccd1 vccd1 _06057_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08708__A2 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _09822_/B _09975_/B vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08479__C _08479_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__A1 _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__nand2_1
X_06958_ _06959_/B _06959_/A vssd1 vssd1 vccd1 vccd1 _06958_/Y sky130_fd_sc_hd__nand2_1
X_09677_ _10450_/A _10456_/A vssd1 vssd1 vccd1 vccd1 _09678_/B sky130_fd_sc_hd__nor2_1
X_05909_ _05928_/A vssd1 vssd1 vccd1 vccd1 _05927_/B sky130_fd_sc_hd__inv_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08495__B _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ _08628_/A _08628_/B vssd1 vssd1 vccd1 vccd1 _08631_/C sky130_fd_sc_hd__nand2_1
X_06889_ _07016_/B _07016_/C _06888_/Y vssd1 vssd1 vccd1 vccd1 _07013_/A sky130_fd_sc_hd__a21oi_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ _08559_/A vssd1 vssd1 vccd1 vccd1 _08559_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07839__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10452_ _10452_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10383_ _10383_/A _10383_/B _10383_/C vssd1 vssd1 vccd1 vccd1 _10384_/C sky130_fd_sc_hd__and3_1
XANTENNA__05359__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06918__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ _07930_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _07933_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09363__A2 _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _07861_/A vssd1 vssd1 vccd1 vccd1 _07970_/A sky130_fd_sc_hd__inv_2
XANTENNA__09980__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ _09853_/B _09600_/B vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06812_ _06812_/A _06812_/B vssd1 vssd1 vccd1 vccd1 _07147_/B sky130_fd_sc_hd__nand2_1
X_07792_ _07792_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07818_/B sky130_fd_sc_hd__nand2_1
X_09531_ _09698_/B _09531_/B vssd1 vssd1 vccd1 vccd1 _09536_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06743_ _06845_/B _06743_/B vssd1 vssd1 vccd1 vccd1 _06744_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _09470_/B _09770_/B vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__nand2_1
X_06674_ _10051_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _06891_/B sky130_fd_sc_hd__nand2_1
X_09393_ input52/X _10111_/B input53/X _10126_/B vssd1 vssd1 vccd1 vccd1 _09394_/B
+ sky130_fd_sc_hd__a22o_1
X_08413_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08651_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05625_ _05979_/B _05979_/A vssd1 vssd1 vccd1 vccd1 _05626_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ _08344_/A vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__inv_2
XFILLER_0_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05556_ _06087_/B _06087_/A vssd1 vssd1 vccd1 vccd1 _05560_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09220__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08275_ _08489_/B _08275_/B vssd1 vssd1 vccd1 vccd1 _08279_/A sky130_fd_sc_hd__nand2_1
X_05487_ _05487_/A _05487_/B vssd1 vssd1 vccd1 vccd1 _05827_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07226_ _07228_/B _07227_/A vssd1 vssd1 vccd1 vccd1 _07229_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07157_ _07157_/A _07709_/B _07709_/A vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__nand3_1
X_06108_ _05684_/A _05687_/A _06107_/Y vssd1 vssd1 vccd1 vccd1 _06585_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07088_ _07088_/A _07088_/B vssd1 vssd1 vccd1 vccd1 _07088_/Y sky130_fd_sc_hd__nor2_1
X_06039_ _06505_/A vssd1 vssd1 vccd1 vccd1 _06040_/B sky130_fd_sc_hd__inv_2
X_09729_ _09718_/Y _09729_/B _09729_/C vssd1 vssd1 vccd1 vccd1 _09730_/B sky130_fd_sc_hd__nand3b_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504_ _10511_/CLK _10504_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ _10435_/A _10435_/B vssd1 vssd1 vccd1 vccd1 _10471_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10366_ _10368_/B hold58/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__and2b_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10295_/Y hold10/X vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_87_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05410_ input64/X vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__buf_4
XFILLER_0_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06664__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06390_ _06810_/A _06809_/A vssd1 vssd1 vccd1 vccd1 _06390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05341_ _05344_/B vssd1 vssd1 vccd1 vccd1 _05346_/A sky130_fd_sc_hd__inv_2
XFILLER_0_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05272_ _09960_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _05554_/B sky130_fd_sc_hd__nand2_1
X_08060_ _08060_/A _08060_/B _08065_/B vssd1 vssd1 vccd1 vccd1 _08079_/B sky130_fd_sc_hd__nand3_1
X_07011_ _07011_/A _07011_/B _07011_/C vssd1 vssd1 vccd1 vccd1 _07623_/C sky130_fd_sc_hd__nand3_1
X_08962_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08967_/B sky130_fd_sc_hd__inv_2
X_08893_ _08893_/A vssd1 vssd1 vccd1 vccd1 _08894_/C sky130_fd_sc_hd__inv_2
X_07913_ _07913_/A _07913_/B vssd1 vssd1 vccd1 vccd1 _07914_/A sky130_fd_sc_hd__nand2_1
X_07844_ _07844_/A _07851_/A vssd1 vssd1 vccd1 vccd1 _07845_/B sky130_fd_sc_hd__nand2_1
X_07775_ _07776_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07779_/B sky130_fd_sc_hd__or2_1
X_09514_ _09514_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06726_ _06937_/B _06936_/A _06936_/B vssd1 vssd1 vccd1 vccd1 _06938_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _09446_/B _09802_/B vssd1 vssd1 vccd1 vccd1 _09451_/A sky130_fd_sc_hd__or2_1
XFILLER_0_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06657_ _06716_/B _06716_/C vssd1 vssd1 vccd1 vccd1 _06715_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05608_ _05608_/A _06093_/B _05608_/C vssd1 vssd1 vccd1 vccd1 _06093_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09376_ _09379_/B _09379_/C vssd1 vssd1 vccd1 vccd1 _09622_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06588_ _06590_/C vssd1 vssd1 vccd1 vccd1 _06589_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08327_ _10044_/A _10084_/D _08326_/C vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__o21ai_1
X_05539_ _05983_/A _05539_/B _05539_/C vssd1 vssd1 vccd1 vccd1 _05540_/B sky130_fd_sc_hd__nand3_1
X_08258_ _08464_/A _08504_/A _08258_/C vssd1 vssd1 vccd1 vccd1 _08262_/C sky130_fd_sc_hd__nand3_1
X_07209_ _07209_/A _07209_/B vssd1 vssd1 vccd1 vccd1 _07359_/B sky130_fd_sc_hd__nand2_1
X_08189_ _08189_/A _08189_/B _08189_/C vssd1 vssd1 vccd1 vccd1 _08191_/A sky130_fd_sc_hd__nor3_1
X_10220_ _10220_/A hold36/X vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__and2_1
XFILLER_0_42_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _09925_/A _09925_/B _09925_/C vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__05637__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ _10082_/A vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__inv_2
XANTENNA__08013__B _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08964__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10418_ _10418_/A vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__inv_2
X_10349_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__and2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05890_ _05890_/A _05890_/B vssd1 vssd1 vccd1 vccd1 _05893_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07560_ _10083_/B _09981_/B vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__nand2_1
X_06511_ _06511_/A _06511_/B vssd1 vssd1 vccd1 vccd1 _06512_/B sky130_fd_sc_hd__nand2_1
X_09230_ _09230_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09231_/C sky130_fd_sc_hd__nand2_1
X_07491_ _08214_/A vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__clkbuf_8
X_06442_ _09816_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _06445_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _09161_/A _09161_/B vssd1 vssd1 vccd1 vccd1 _09172_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06373_ _06363_/Y _06746_/B _06372_/Y vssd1 vssd1 vccd1 vccd1 _06736_/A sky130_fd_sc_hd__a21oi_1
X_09092_ _09381_/A _09092_/B vssd1 vssd1 vccd1 vccd1 _09094_/A sky130_fd_sc_hd__nand2_1
X_08112_ _08112_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _08112_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05324_ _05324_/A _05324_/B vssd1 vssd1 vccd1 vccd1 _05376_/B sky130_fd_sc_hd__nand2_1
X_08043_ _08091_/B _08091_/C vssd1 vssd1 vccd1 vccd1 _08123_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05255_ input13/X vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__buf_4
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05738__A input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09994_ _09995_/B _09995_/A vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__or2_1
X_08945_ _08948_/B _09332_/B _08945_/C vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__nand3b_1
X_08876_ _08876_/A _09096_/B _08876_/C vssd1 vssd1 vccd1 vccd1 _09096_/A sky130_fd_sc_hd__nand3_1
X_07827_ _07846_/A _07846_/C vssd1 vssd1 vccd1 vccd1 _07836_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07758_ _07823_/B _07821_/B vssd1 vssd1 vccd1 vccd1 _07812_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08784__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06709_ _06946_/C vssd1 vssd1 vccd1 vccd1 _06710_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07689_ _07689_/A _07692_/B vssd1 vssd1 vccd1 vccd1 _07693_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09428_ _09431_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09429_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ _09039_/A _09038_/B _09358_/Y vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_81_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05367__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ _10203_/A hold76/X vssd1 vssd1 vccd1 vccd1 _10207_/B sky130_fd_sc_hd__and2_1
XFILLER_0_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _10134_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10134_/Y sky130_fd_sc_hd__nor2_1
X_10065_ _10067_/C vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__inv_2
XANTENNA__06479__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07773__A _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _07137_/A _07138_/A vssd1 vssd1 vccd1 vccd1 _06991_/Y sky130_fd_sc_hd__nand2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08730_/A vssd1 vssd1 vccd1 vccd1 _08735_/A sky130_fd_sc_hd__inv_2
XANTENNA__07492__B _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05942_ _10026_/B _08214_/A vssd1 vssd1 vccd1 vccd1 _06341_/C sky130_fd_sc_hd__nand2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__A2 _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ _09189_/A _09190_/B vssd1 vssd1 vccd1 vccd1 _08662_/A sky130_fd_sc_hd__nand2_1
X_05873_ _05875_/B vssd1 vssd1 vccd1 vccd1 _05874_/B sky130_fd_sc_hd__inv_2
X_07612_ _07898_/C _07898_/B vssd1 vssd1 vccd1 vccd1 _07899_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08592_ _08594_/C vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07543_ _07545_/A _07545_/B vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10085__A2 _09720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _07474_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09213_ _09213_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _09215_/B sky130_fd_sc_hd__xor2_1
X_06425_ _06425_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09144_ _09144_/A _09144_/B _09144_/C vssd1 vssd1 vccd1 vccd1 _09162_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07948__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06356_ _06358_/A _06358_/C vssd1 vssd1 vccd1 vccd1 _06357_/A sky130_fd_sc_hd__nand2_1
X_09075_ _10084_/A _10113_/D _09075_/C vssd1 vssd1 vccd1 vccd1 _09077_/A sky130_fd_sc_hd__nor3_1
X_05307_ _09533_/B _07216_/B vssd1 vssd1 vccd1 vccd1 _05308_/B sky130_fd_sc_hd__nand2_1
X_06287_ _06287_/A vssd1 vssd1 vccd1 vccd1 _06707_/B sky130_fd_sc_hd__inv_2
X_08026_ _08027_/A _08027_/B _08026_/C vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__nand3_1
X_05238_ _05243_/B _05311_/A vssd1 vssd1 vccd1 vccd1 _05242_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _09976_/B _09977_/B _09977_/C vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__nand3b_1
X_08928_ _08930_/A vssd1 vssd1 vccd1 vccd1 _08929_/B sky130_fd_sc_hd__inv_2
X_08859_ _08857_/Y _08589_/B _08858_/Y vssd1 vssd1 vccd1 vccd1 _08887_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09466__A1 _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08961__B _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07858__A _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06762__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08689__A _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__nand2_1
X_10048_ _10048_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__nand2_1
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09313__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06210_ _05969_/Y _06209_/Y _05900_/A vssd1 vssd1 vccd1 vccd1 _06810_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07190_ _07236_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07234_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06672__A _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06141_ _10044_/A _10113_/B _06137_/Y vssd1 vssd1 vccd1 vccd1 _06146_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06072_ _06072_/A _06072_/B vssd1 vssd1 vccd1 vccd1 _06077_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _09904_/B sky130_fd_sc_hd__or2_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09831_ _09830_/B _09831_/B _09831_/C vssd1 vssd1 vccd1 vccd1 _09832_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__09393__B1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09762_ _09762_/A _09762_/B _09762_/C vssd1 vssd1 vccd1 vccd1 _09762_/Y sky130_fd_sc_hd__nor3_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _09963_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _06977_/B sky130_fd_sc_hd__nand2_1
X_08713_ _08717_/A _08932_/A vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__nand2_1
X_05925_ _05925_/A _05925_/B vssd1 vssd1 vccd1 vccd1 _06331_/C sky130_fd_sc_hd__nand2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _09501_/A _09692_/Y _09500_/A vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_96_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08644_ _08644_/A _08644_/B vssd1 vssd1 vccd1 vccd1 _08647_/A sky130_fd_sc_hd__nand2_1
X_05856_ _09313_/D vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__buf_6
X_08575_ _08575_/A _08575_/B _08575_/C vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_49_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05787_ _05787_/A _05787_/B _05787_/C vssd1 vssd1 vccd1 vccd1 _05809_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_49_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07526_ _07527_/A _07526_/B _07527_/B vssd1 vssd1 vccd1 vccd1 _07614_/B sky130_fd_sc_hd__nand3_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07457_ _07457_/A vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__inv_2
X_06408_ _06408_/A _06463_/A vssd1 vssd1 vccd1 vccd1 _06468_/B sky130_fd_sc_hd__nand2_1
X_07388_ _07059_/Y _07349_/B _07085_/Y vssd1 vssd1 vccd1 vccd1 _07391_/B sky130_fd_sc_hd__a21o_1
X_09127_ _09127_/A _09127_/B vssd1 vssd1 vccd1 vccd1 _09136_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06339_ _06339_/A vssd1 vssd1 vccd1 vccd1 _06342_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09058_ _09060_/C vssd1 vssd1 vccd1 vccd1 _09059_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08009_ _08010_/B _08010_/A vssd1 vssd1 vccd1 vccd1 _08095_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09687__B2 _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__A1 _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08972__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06492__A _09960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07100__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput80 hold66/A vssd1 vssd1 vccd1 vccd1 y_o[22] sky130_fd_sc_hd__buf_12
Xoutput91 _10483_/Q vssd1 vssd1 vccd1 vccd1 y_o[3] sky130_fd_sc_hd__buf_12
XFILLER_0_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08866__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05710_ _05712_/A _05712_/B vssd1 vssd1 vccd1 vccd1 _05711_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06667__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ _06928_/C vssd1 vssd1 vccd1 vccd1 _06930_/B sky130_fd_sc_hd__inv_2
X_05641_ _05643_/B vssd1 vssd1 vccd1 vccd1 _05642_/B sky130_fd_sc_hd__inv_2
X_08360_ _08363_/B _08363_/C vssd1 vssd1 vccd1 vccd1 _08362_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07311_ _07313_/C vssd1 vssd1 vccd1 vccd1 _07312_/B sky130_fd_sc_hd__inv_2
X_05572_ _05981_/A _06022_/A _05572_/C vssd1 vssd1 vccd1 vccd1 _05574_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08291_ _09227_/A _10044_/D _08289_/C vssd1 vssd1 vccd1 vccd1 _08292_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07242_ _07475_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07474_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07173_ _07173_/A _07173_/B vssd1 vssd1 vccd1 vccd1 _07237_/B sky130_fd_sc_hd__nand2_1
X_06124_ _05605_/C _05605_/B _06121_/Y vssd1 vssd1 vccd1 vccd1 _06128_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_26_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06055_ _09963_/A _10052_/A vssd1 vssd1 vccd1 vccd1 _06058_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09814_ _09957_/A _09814_/B _09814_/C vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06719__A2 _09392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ _09745_/A _09745_/B _09745_/C vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06957_ _07001_/B _07000_/A vssd1 vssd1 vccd1 vccd1 _06957_/Y sky130_fd_sc_hd__nand2_1
X_09676_ _09676_/A _09676_/B vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__nand2_1
X_06888_ _07024_/A _07023_/A vssd1 vssd1 vccd1 vccd1 _06888_/Y sky130_fd_sc_hd__nor2_1
X_05908_ _05908_/A _05908_/B _05908_/C vssd1 vssd1 vccd1 vccd1 _05916_/A sky130_fd_sc_hd__nand3_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _08627_/A _08627_/B vssd1 vssd1 vccd1 vccd1 _09150_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05481__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05839_ _05947_/A _05948_/A vssd1 vssd1 vccd1 vccd1 _05919_/B sky130_fd_sc_hd__nand2_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _08558_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08563_/A sky130_fd_sc_hd__nand2_1
X_08489_ _08489_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08490_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07509_ _07511_/B _07511_/C vssd1 vssd1 vccd1 vccd1 _07510_/A sky130_fd_sc_hd__nand2_1
X_10451_ _10452_/B _10452_/A vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__or2_1
X_10382_ hold45/X vssd1 vssd1 vccd1 vccd1 _10480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05656__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06487__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07860_ _07860_/A _07861_/A vssd1 vssd1 vccd1 vccd1 _07936_/C sky130_fd_sc_hd__nand2_1
X_06811_ _06813_/B _06813_/C vssd1 vssd1 vccd1 vccd1 _06812_/A sky130_fd_sc_hd__nand2_1
X_07791_ _07792_/B _07792_/A vssd1 vssd1 vccd1 vccd1 _07889_/B sky130_fd_sc_hd__nor2_2
X_09530_ _09528_/A _10026_/B _09685_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09531_/B
+ sky130_fd_sc_hd__a22o_1
X_06742_ _06743_/B _06742_/B _06742_/C vssd1 vssd1 vccd1 vccd1 _06845_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09461_ _09461_/A _09461_/B _09461_/C vssd1 vssd1 vccd1 vccd1 _09770_/B sky130_fd_sc_hd__nand3_2
X_06673_ _06892_/B vssd1 vssd1 vccd1 vccd1 _06891_/A sky130_fd_sc_hd__inv_2
X_09392_ _10113_/A _10113_/C _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09634_/B
+ sky130_fd_sc_hd__or4_2
X_08412_ _08652_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08651_/A sky130_fd_sc_hd__nand2_1
X_05624_ _05499_/A _05334_/B _05500_/Y vssd1 vssd1 vccd1 vccd1 _05979_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ _08331_/Y _08333_/Y _08344_/A vssd1 vssd1 vccd1 vccd1 _08346_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05555_ _05281_/C _05281_/B _05554_/Y vssd1 vssd1 vccd1 vccd1 _06087_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__09220__B _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ _08274_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05486_ _05478_/Y _05486_/B _05486_/C vssd1 vssd1 vccd1 vccd1 _05487_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ _07225_/A _07225_/B vssd1 vssd1 vccd1 vccd1 _07417_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07956__A _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07156_ _07709_/A _07709_/B _07157_/A vssd1 vssd1 vccd1 vccd1 _07156_/Y sky130_fd_sc_hd__a21oi_1
X_06107_ _06107_/A _06107_/B vssd1 vssd1 vccd1 vccd1 _06107_/Y sky130_fd_sc_hd__nor2_1
X_07087_ _07391_/A _07392_/A vssd1 vssd1 vccd1 vccd1 _07390_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05476__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06038_ _05534_/C _05534_/B _06037_/Y vssd1 vssd1 vccd1 vccd1 _06505_/A sky130_fd_sc_hd__a21oi_2
Xfanout100 fanout99/A vssd1 vssd1 vccd1 vccd1 fanout100/X sky130_fd_sc_hd__clkbuf_8
X_09728_ _09728_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09729_/C sky130_fd_sc_hd__nand2_1
X_07989_ _07989_/A _07989_/B _07989_/C vssd1 vssd1 vccd1 vccd1 _07990_/B sky130_fd_sc_hd__nand3_1
X_09659_ _09661_/A vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__inv_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ _10509_/CLK hold48/X fanout100/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfrtp_1
X_10434_ _10434_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10435_/B sky130_fd_sc_hd__nand2_1
X_10365_ _10365_/A _10365_/B vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__nand2_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05386__A _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10496_/Q hold9/X vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__nand2_1
XANTENNA__06010__A _09960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06664__B _09981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05340_ _05908_/B _05908_/C vssd1 vssd1 vccd1 vccd1 _05913_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05271_ _05554_/A vssd1 vssd1 vccd1 vccd1 _05274_/A sky130_fd_sc_hd__inv_2
XFILLER_0_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07010_ _07010_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07623_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ _09960_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08892_ _08892_/A _08893_/A vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__nand2_1
X_07912_ _07912_/A _08071_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__nand3_1
X_07843_ _07851_/A _07844_/A vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__or2_1
XFILLER_0_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07774_ _08337_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _07776_/B sky130_fd_sc_hd__nand2_1
X_09513_ _09330_/C _09330_/B _09320_/Y vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06725_ _06725_/A _06725_/B vssd1 vssd1 vccd1 vccd1 _06936_/B sky130_fd_sc_hd__nand2_1
X_09444_ _09789_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06656_ _06656_/A _06656_/B _06656_/C vssd1 vssd1 vccd1 vccd1 _06716_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05607_ _05611_/C vssd1 vssd1 vccd1 vccd1 _05608_/C sky130_fd_sc_hd__inv_2
X_09375_ _09375_/A _09375_/B _09375_/C vssd1 vssd1 vccd1 vccd1 _09379_/C sky130_fd_sc_hd__nand3_1
X_06587_ _06587_/A _06587_/B vssd1 vssd1 vccd1 vccd1 _06590_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08326_ _10044_/A _10084_/D _08326_/C vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05538_ _05983_/B _05538_/B vssd1 vssd1 vccd1 vccd1 _05540_/A sky130_fd_sc_hd__nand2_1
X_08257_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__inv_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05469_ input35/X _08810_/B vssd1 vssd1 vccd1 vccd1 _05870_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ _10383_/A _08188_/B _08188_/C vssd1 vssd1 vccd1 vccd1 _08189_/C sky130_fd_sc_hd__nand3_1
X_07208_ _07208_/A _07209_/B _07209_/A vssd1 vssd1 vccd1 vccd1 _07222_/A sky130_fd_sc_hd__nand3_1
X_07139_ _07680_/A _07680_/B vssd1 vssd1 vccd1 vccd1 _07679_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10150_ _10154_/B _10154_/C vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _09723_/X _09725_/A _09724_/A vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08964__B _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09141__A _09141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10417_ _10417_/A _10417_/B vssd1 vssd1 vccd1 vccd1 _10467_/D sky130_fd_sc_hd__xnor2_1
X_10348_ _10349_/B _10349_/A vssd1 vssd1 vccd1 vccd1 _10376_/B sky130_fd_sc_hd__nor2_2
XANTENNA__06005__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _10299_/C hold33/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__xor2_1
XANTENNA__09723__B1 _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05844__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06510_ _06513_/B _06513_/C vssd1 vssd1 vccd1 vccd1 _06512_/A sky130_fd_sc_hd__nand2_1
X_07490_ _07503_/B _07503_/C vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06441_ _08247_/B vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__buf_12
XFILLER_0_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _09171_/A _09171_/B _09172_/C vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09986__A _09986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06372_ _06739_/A _06744_/A vssd1 vssd1 vccd1 vccd1 _06372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ _09091_/A _09381_/A _09092_/B vssd1 vssd1 vccd1 vccd1 _09385_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08111_ _08112_/B _08112_/A vssd1 vssd1 vccd1 vccd1 _08158_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05323_ _05377_/B vssd1 vssd1 vccd1 vccd1 _05325_/B sky130_fd_sc_hd__inv_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08042_ _08042_/A _08042_/B vssd1 vssd1 vccd1 vccd1 _08091_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05254_ _05503_/A vssd1 vssd1 vccd1 vccd1 _05263_/A sky130_fd_sc_hd__inv_2
XFILLER_0_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _09993_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ _08947_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08945_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09226__A _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05754__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _08875_/A _08875_/B vssd1 vssd1 vccd1 vccd1 _08877_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07826_ _07826_/A _07826_/B vssd1 vssd1 vccd1 vccd1 _07846_/C sky130_fd_sc_hd__nand2_1
X_07757_ _07821_/A _07821_/B _07757_/C vssd1 vssd1 vccd1 vccd1 _07823_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_79_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08784__B _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ _06708_/A _06708_/B vssd1 vssd1 vccd1 vccd1 _06946_/C sky130_fd_sc_hd__nand2_1
X_07688_ _07688_/A _07707_/B _07688_/C vssd1 vssd1 vccd1 vccd1 _07694_/A sky130_fd_sc_hd__nand3_1
X_09427_ _09427_/A _09669_/A _09427_/C vssd1 vssd1 vccd1 vccd1 _09674_/B sky130_fd_sc_hd__nand3_1
X_06639_ _06639_/A _06639_/B _06820_/C vssd1 vssd1 vccd1 vccd1 _06640_/B sky130_fd_sc_hd__nand3_2
X_09358_ _09358_/A vssd1 vssd1 vccd1 vccd1 _09358_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08309_ _08309_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08315_/B sky130_fd_sc_hd__nand2_1
X_09289_ _09762_/A _09777_/B _09289_/C vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10490__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ _10484_/Q hold75/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__nand2_1
X_10133_ _10134_/B _10134_/A vssd1 vssd1 vccd1 vccd1 _10133_/Y sky130_fd_sc_hd__nand2_1
X_10064_ _10062_/Y _09830_/B _10063_/Y vssd1 vssd1 vccd1 vccd1 _10067_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__06479__B _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08747__A1 _09227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07773__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06990_ _06957_/Y _07003_/B _06989_/Y vssd1 vssd1 vccd1 vccd1 _07138_/A sky130_fd_sc_hd__a21oi_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05941_ _06340_/B _06339_/A vssd1 vssd1 vccd1 vccd1 _06343_/C sky130_fd_sc_hd__nand2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _08668_/C _09180_/B _08660_/C vssd1 vssd1 vccd1 vccd1 _09190_/B sky130_fd_sc_hd__nand3b_1
X_05872_ _05875_/A _05875_/C vssd1 vssd1 vccd1 vccd1 _05874_/A sky130_fd_sc_hd__nand2_1
X_07611_ _07523_/B _07611_/B _07611_/C vssd1 vssd1 vccd1 vccd1 _07898_/C sky130_fd_sc_hd__nand3b_1
X_08591_ _08591_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _08594_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07542_ _07542_/A _07542_/B vssd1 vssd1 vccd1 vccd1 _07545_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07473_ _07475_/C vssd1 vssd1 vccd1 vccd1 _07474_/B sky130_fd_sc_hd__inv_2
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09212_ _09210_/X _09212_/B vssd1 vssd1 vccd1 vccd1 _09213_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_63_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06424_ _06426_/B vssd1 vssd1 vccd1 vccd1 _06425_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09143_ _09143_/A _09143_/B vssd1 vssd1 vccd1 vccd1 _09162_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06355_ _06355_/A _06355_/B vssd1 vssd1 vccd1 vccd1 _06358_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07948__B _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05306_ input63/X vssd1 vssd1 vccd1 vccd1 _07216_/B sky130_fd_sc_hd__buf_6
X_09074_ input50/X _10112_/B vssd1 vssd1 vccd1 vccd1 _09075_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06286_ _09960_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _06287_/A sky130_fd_sc_hd__nand2_1
X_08025_ _08025_/A _08025_/B vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__nand2_1
X_05237_ _05311_/B vssd1 vssd1 vccd1 vccd1 _05243_/B sky130_fd_sc_hd__inv_2
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09976_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__nand2_1
X_08927_ _08927_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__nand2_1
X_08858_ _08858_/A _08858_/B vssd1 vssd1 vccd1 vccd1 _08858_/Y sky130_fd_sc_hd__nor2_1
X_07809_ _07809_/A _07809_/B _07809_/C vssd1 vssd1 vccd1 vccd1 _07810_/B sky130_fd_sc_hd__nand3_1
X_08789_ _09227_/A _10044_/B _08790_/C vssd1 vssd1 vccd1 vccd1 _08789_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07858__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__B _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05659__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07874__A _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__B _09998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _10116_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__xnor2_1
X_10047_ _10047_/A _10047_/B vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__xnor2_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09313__B _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06672__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06140_ _09361_/C vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__inv_2
X_06071_ _06484_/B vssd1 vssd1 vccd1 vccd1 _06072_/B sky130_fd_sc_hd__inv_2
XFILLER_0_53_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09393__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _09830_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _09832_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09393__B2 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09981_/B input19/X vssd1 vssd1 vccd1 vccd1 _09762_/C sky130_fd_sc_hd__nand2_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _06977_/A vssd1 vssd1 vccd1 vccd1 _06976_/A sky130_fd_sc_hd__inv_2
X_08712_ _08711_/B _08932_/B _08712_/C vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__nand3b_1
X_05924_ _05924_/A _05924_/B _05924_/C vssd1 vssd1 vccd1 vccd1 _05925_/B sky130_fd_sc_hd__nand3_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _09692_/A vssd1 vssd1 vccd1 vccd1 _09692_/Y sky130_fd_sc_hd__inv_2
X_08643_ _08645_/B _08645_/C vssd1 vssd1 vccd1 vccd1 _08644_/A sky130_fd_sc_hd__nand2_1
X_05855_ _08810_/B vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__buf_6
X_08574_ _08574_/A vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__inv_2
XFILLER_0_49_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05786_ _05786_/A _05786_/B vssd1 vssd1 vccd1 vccd1 _05974_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07525_ _07525_/A vssd1 vssd1 vccd1 vccd1 _07527_/A sky130_fd_sc_hd__inv_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07456_ _10111_/B _08866_/B _09485_/C _09804_/A vssd1 vssd1 vccd1 vccd1 _07457_/A
+ sky130_fd_sc_hd__and4_1
X_06407_ _06405_/Y _06048_/B _06406_/Y vssd1 vssd1 vccd1 vccd1 _06517_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07387_ _07385_/Y _07373_/B _07386_/Y vssd1 vssd1 vccd1 vccd1 _07631_/A sky130_fd_sc_hd__a21oi_1
X_09126_ _09414_/B _09126_/B vssd1 vssd1 vccd1 vccd1 _09127_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06338_ _06342_/A _06339_/A vssd1 vssd1 vccd1 vccd1 _06341_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ _09057_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _09060_/C sky130_fd_sc_hd__nor2_1
X_06269_ _06269_/A _06269_/B vssd1 vssd1 vccd1 vccd1 _06658_/C sky130_fd_sc_hd__nand2_1
X_08008_ _08004_/X _08006_/Y _08102_/A vssd1 vssd1 vccd1 vccd1 _08010_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09959_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__and2_1
XANTENNA__09687__A2 _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05942__A _10026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08972__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06492__B _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05389__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput70 _10493_/Q vssd1 vssd1 vccd1 vccd1 y_o[13] sky130_fd_sc_hd__buf_12
Xoutput81 hold46/A vssd1 vssd1 vccd1 vccd1 y_o[23] sky130_fd_sc_hd__buf_12
Xoutput92 _10484_/Q vssd1 vssd1 vccd1 vccd1 y_o[4] sky130_fd_sc_hd__buf_12
XANTENNA__09324__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05640_ _09528_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _05643_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06667__B _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05571_ _05571_/A _05571_/B _05571_/C vssd1 vssd1 vccd1 vccd1 _05628_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07310_ _07380_/B _07310_/B vssd1 vssd1 vccd1 vccd1 _07313_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08290_ _08290_/A vssd1 vssd1 vccd1 vccd1 _08292_/A sky130_fd_sc_hd__inv_2
XFILLER_0_73_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07241_ _07188_/Y _07241_/B _07241_/C vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_54_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07172_ _07172_/A _07172_/B _07172_/C vssd1 vssd1 vccd1 vccd1 _07173_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06123_ _06128_/A _06129_/B vssd1 vssd1 vccd1 vccd1 _06127_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06054_ input37/X _09022_/C vssd1 vssd1 vccd1 vccd1 _06058_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ _09813_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__nand2_1
X_09744_ _09744_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__nand2_1
X_06956_ _06916_/Y _07010_/B _06955_/Y vssd1 vssd1 vccd1 vccd1 _07000_/A sky130_fd_sc_hd__a21oi_2
X_09675_ _09674_/B _09675_/B _09941_/B vssd1 vssd1 vccd1 vccd1 _09676_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06887_ _07025_/C vssd1 vssd1 vccd1 vccd1 _07016_/C sky130_fd_sc_hd__inv_2
X_05907_ _05907_/A _05907_/B vssd1 vssd1 vccd1 vccd1 _05969_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08626_ _08628_/B vssd1 vssd1 vccd1 vccd1 _08627_/B sky130_fd_sc_hd__inv_2
X_05838_ _05947_/B vssd1 vssd1 vccd1 vccd1 _05948_/A sky130_fd_sc_hd__inv_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08557_ _08551_/Y _08557_/B _08557_/C vssd1 vssd1 vccd1 vccd1 _08558_/B sky130_fd_sc_hd__nand3b_1
X_05769_ _05787_/C vssd1 vssd1 vccd1 vccd1 _05770_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ _08488_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08501_/B sky130_fd_sc_hd__nand2_1
X_07508_ _07508_/A _07508_/B _07508_/C vssd1 vssd1 vccd1 vccd1 _07511_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07439_ _07439_/A vssd1 vssd1 vccd1 vccd1 _07441_/B sky130_fd_sc_hd__inv_2
XFILLER_0_91_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10450_ _10450_/A vssd1 vssd1 vccd1 vccd1 _10452_/B sky130_fd_sc_hd__inv_2
X_09109_ _09115_/B _09406_/A vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ hold44/X _10381_/B vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__and2_1
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05656__B _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06487__B _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05847__A _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07790_ _07807_/B _07790_/B vssd1 vssd1 vccd1 vccd1 _07792_/A sky130_fd_sc_hd__and2_1
X_06810_ _06810_/A _06810_/B _06810_/C vssd1 vssd1 vccd1 vccd1 _06813_/C sky130_fd_sc_hd__nand3_1
X_06741_ _06749_/B _06750_/C _06750_/B vssd1 vssd1 vccd1 vccd1 _06743_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09460_ _09461_/A _09461_/C _09461_/B vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__a21o_1
X_08411_ _08410_/B _08411_/B _08411_/C vssd1 vssd1 vccd1 vccd1 _08652_/B sky130_fd_sc_hd__nand3b_1
X_06672_ _10050_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _06892_/B sky130_fd_sc_hd__nand2_1
X_09391_ input53/X vssd1 vssd1 vccd1 vccd1 _10113_/C sky130_fd_sc_hd__inv_2
XFILLER_0_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05623_ _05628_/B _05628_/C vssd1 vssd1 vccd1 vccd1 _05979_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08342_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__xor2_1
X_05554_ _05554_/A _05554_/B vssd1 vssd1 vccd1 vccd1 _05554_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08273_ _08274_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _08489_/B sky130_fd_sc_hd__or2_1
X_05485_ _05485_/A vssd1 vssd1 vccd1 vccd1 _05486_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09220__C _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07224_ _07229_/C vssd1 vssd1 vccd1 vccd1 _07225_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07956__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _07710_/B vssd1 vssd1 vccd1 vccd1 _07157_/A sky130_fd_sc_hd__inv_2
X_06106_ _06183_/A _06183_/B vssd1 vssd1 vccd1 vccd1 _06182_/A sky130_fd_sc_hd__nand2_1
X_07086_ _07059_/Y _07349_/B _07085_/Y vssd1 vssd1 vccd1 vccd1 _07392_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__05476__B _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06037_ _06037_/A _06037_/B vssd1 vssd1 vccd1 vccd1 _06037_/Y sky130_fd_sc_hd__nor2_1
Xfanout101 input65/X vssd1 vssd1 vccd1 vccd1 fanout99/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07988_ _07988_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07990_/A sky130_fd_sc_hd__nand2_1
X_09727_ _09727_/A vssd1 vssd1 vccd1 vccd1 _09729_/B sky130_fd_sc_hd__inv_2
X_06939_ _07090_/B vssd1 vssd1 vccd1 vccd1 _06940_/B sky130_fd_sc_hd__inv_2
XFILLER_0_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09658_ _09658_/A _09658_/B vssd1 vssd1 vccd1 vccd1 _09661_/A sky130_fd_sc_hd__nand2_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09589_ _09589_/A _09845_/A vssd1 vssd1 vccd1 vccd1 _09591_/A sky130_fd_sc_hd__nand2_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ input49/X _10111_/B input50/X _08866_/B vssd1 vssd1 vccd1 vccd1 _08610_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10502_ _10511_/CLK _10502_/D fanout100/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10433_ _10433_/A vssd1 vssd1 vccd1 vccd1 _10470_/D sky130_fd_sc_hd__clkbuf_1
X_10364_ _10365_/B _10365_/A vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09139__A _09141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05667__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05386__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _10496_/Q hold9/X vssd1 vssd1 vccd1 vccd1 _10295_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06010__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05270_ _09816_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _05554_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08960_ _08958_/Y _08720_/B _08959_/Y vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08891_ _09132_/B _08894_/B vssd1 vssd1 vccd1 vccd1 _08892_/A sky130_fd_sc_hd__nand2_1
X_07911_ _07911_/A _07911_/B _07914_/B vssd1 vssd1 vccd1 vccd1 _08071_/B sky130_fd_sc_hd__nand3_2
X_07842_ _07842_/A _07841_/Y vssd1 vssd1 vccd1 vccd1 _07844_/A sky130_fd_sc_hd__nor2b_1
X_09512_ _09515_/B _09515_/C vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__nand2_1
X_07773_ _08862_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _07776_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06724_ _06725_/A _06725_/B vssd1 vssd1 vccd1 vccd1 _06936_/A sky130_fd_sc_hd__or2_1
XFILLER_0_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09443_ _09443_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09444_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06655_ _06823_/B _06823_/C vssd1 vssd1 vccd1 vccd1 _06825_/A sky130_fd_sc_hd__nand2_1
X_09374_ _09375_/A _09375_/C _09375_/B vssd1 vssd1 vccd1 vccd1 _09379_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09257__B1 _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05606_ _05606_/A _05606_/B vssd1 vssd1 vccd1 vccd1 _05611_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08325_ _09548_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08326_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06586_ _06586_/A vssd1 vssd1 vccd1 vccd1 _06587_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05537_ _06022_/B _05537_/B _05537_/C vssd1 vssd1 vccd1 vccd1 _06022_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08256_ _08504_/B _08257_/A vssd1 vssd1 vccd1 vccd1 _08262_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05468_ _05866_/A _05867_/A vssd1 vssd1 vccd1 vccd1 _05871_/C sky130_fd_sc_hd__nand2_1
X_08187_ _10383_/C _10383_/B _08186_/A vssd1 vssd1 vccd1 vccd1 _08188_/C sky130_fd_sc_hd__a21o_1
X_07207_ _07207_/A _07207_/B _07207_/C vssd1 vssd1 vccd1 vccd1 _07209_/A sky130_fd_sc_hd__nand3_1
X_07138_ _07138_/A _07138_/B _07138_/C vssd1 vssd1 vccd1 vccd1 _07680_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05399_ _05399_/A _05399_/B _05399_/C vssd1 vssd1 vccd1 vccd1 _05400_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ _07206_/B vssd1 vssd1 vccd1 vccd1 _07205_/A sky130_fd_sc_hd__inv_2
X_10080_ _10149_/A _10149_/C vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06111__A _09528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10416_ _10416_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10417_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10347_ hold46/X vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__inv_2
XANTENNA__06005__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10278_ _10278_/A hold32/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__nand2_1
XANTENNA__09723__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__B2 _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05844__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__B1 _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05860__A _10050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06440_ _06468_/B _06467_/B _06467_/C vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06371_ _06747_/C vssd1 vssd1 vccd1 vccd1 _06746_/B sky130_fd_sc_hd__inv_2
X_09090_ _09090_/A _09090_/B vssd1 vssd1 vccd1 vccd1 _09092_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _08137_/B _08138_/A _08109_/Y vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__a21oi_1
X_05322_ _10043_/B _07216_/B vssd1 vssd1 vccd1 vccd1 _05377_/B sky130_fd_sc_hd__nand2_1
X_08041_ _08037_/B _08036_/B _07980_/Y vssd1 vssd1 vccd1 vccd1 _08042_/B sky130_fd_sc_hd__a21oi_1
X_05253_ _09963_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _05503_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__xor2_1
X_08943_ _08944_/B _08947_/A vssd1 vssd1 vccd1 vccd1 _09332_/B sky130_fd_sc_hd__or2_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05754__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08874_ _08876_/A _09096_/B vssd1 vssd1 vccd1 vccd1 _08875_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07825_ _07826_/A _07740_/A vssd1 vssd1 vccd1 vccd1 _07846_/A sky130_fd_sc_hd__or2b_1
X_07756_ _07822_/B vssd1 vssd1 vccd1 vccd1 _07757_/C sky130_fd_sc_hd__inv_2
X_06707_ _06288_/Y _06707_/B _06707_/C vssd1 vssd1 vccd1 vccd1 _06708_/B sky130_fd_sc_hd__nand3b_1
X_09426_ _09426_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _09431_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ _07690_/B _07692_/B _07690_/C vssd1 vssd1 vccd1 vccd1 _07688_/C sky130_fd_sc_hd__nand3_1
X_06638_ _06638_/A _08656_/A _06638_/C vssd1 vssd1 vccd1 vccd1 _06639_/B sky130_fd_sc_hd__nand3_1
X_09357_ _09357_/A vssd1 vssd1 vccd1 vccd1 _09378_/B sky130_fd_sc_hd__inv_2
X_06569_ _08399_/B _06569_/B _06569_/C vssd1 vssd1 vccd1 vccd1 _08399_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ input17/X vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08308_ _08307_/B _08308_/B _08308_/C vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_34_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08239_ _08239_/A vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__inv_2
XFILLER_0_50_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10201_ _10484_/Q hold75/X vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__or2_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _10138_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__nand2_1
X_10063_ _10063_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _10063_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05855__A _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05940_ _09816_/B _09988_/A vssd1 vssd1 vccd1 vccd1 _06339_/A sky130_fd_sc_hd__nand2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10508__CLK _10509_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05871_ _05871_/A _05871_/B _05871_/C vssd1 vssd1 vccd1 vccd1 _05875_/C sky130_fd_sc_hd__nand3_1
X_08590_ _08589_/B _08590_/B _08590_/C vssd1 vssd1 vccd1 vccd1 _08591_/B sky130_fd_sc_hd__nand3b_1
X_07610_ _07610_/A _07610_/B vssd1 vssd1 vccd1 vccd1 _07611_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06686__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ _07573_/B _07571_/B vssd1 vssd1 vccd1 vccd1 _07542_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07472_ _07534_/B _07534_/C vssd1 vssd1 vccd1 vccd1 _07533_/A sky130_fd_sc_hd__nand2_1
X_09211_ input46/X _09720_/B _10051_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _09212_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06423_ _08422_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _06426_/B sky130_fd_sc_hd__nand2_1
X_09142_ _09144_/A _09144_/B vssd1 vssd1 vccd1 vccd1 _09143_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06354_ _06354_/A vssd1 vssd1 vccd1 vccd1 _06355_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05305_ input4/X vssd1 vssd1 vccd1 vccd1 _09533_/B sky130_fd_sc_hd__buf_6
XFILLER_0_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09073_ _09073_/A vssd1 vssd1 vccd1 vccd1 _09079_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06285_ _06288_/A _06288_/B vssd1 vssd1 vccd1 vccd1 _06707_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08024_ _08024_/A vssd1 vssd1 vccd1 vccd1 _08025_/B sky130_fd_sc_hd__inv_2
X_05236_ _05243_/A _05311_/B vssd1 vssd1 vccd1 vccd1 _05242_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09975_ _09975_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08141__A _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _08930_/B _09277_/A vssd1 vssd1 vccd1 vccd1 _08929_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08857_ _08858_/B _08858_/A vssd1 vssd1 vccd1 vccd1 _08857_/Y sky130_fd_sc_hd__nand2_1
X_07808_ _07808_/A _07808_/B vssd1 vssd1 vccd1 vccd1 _07810_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08788_ input5/X vssd1 vssd1 vccd1 vccd1 _10044_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07739_ _08825_/B input55/X vssd1 vssd1 vccd1 vccd1 _07740_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _09664_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05659__B _09361_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10115_ _10115_/A _10115_/B vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10046_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10047_/B sky130_fd_sc_hd__nand2_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09313__C _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06070_ _09684_/B _08272_/B vssd1 vssd1 vccd1 vccd1 _06484_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05585__A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__A2 _10111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09760_ _09980_/A input18/X vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__nand2_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _09962_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _06977_/A sky130_fd_sc_hd__nand2_1
X_09691_ _10034_/A _09696_/C vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__nand2_1
X_08711_ _08711_/A _08711_/B vssd1 vssd1 vccd1 vccd1 _08717_/A sky130_fd_sc_hd__nand2_1
X_05923_ _05923_/A _05923_/B vssd1 vssd1 vccd1 vccd1 _05925_/A sky130_fd_sc_hd__nand2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08642_ _09166_/A _08642_/B _08642_/C vssd1 vssd1 vccd1 vccd1 _08645_/C sky130_fd_sc_hd__nand3_1
XANTENNA__07156__A1 _07709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05854_ _05959_/A _05960_/A vssd1 vssd1 vccd1 vccd1 _05854_/Y sky130_fd_sc_hd__nand2_1
X_08573_ _08573_/A _08574_/A vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07305__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05785_ _05785_/A _05785_/B _05785_/C vssd1 vssd1 vccd1 vccd1 _05786_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07524_ _07898_/B _07524_/B vssd1 vssd1 vccd1 vccd1 _07530_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07455_ _07520_/B _07463_/B vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__nand2_1
X_06406_ _06406_/A _06406_/B vssd1 vssd1 vccd1 vccd1 _06406_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07386_ _07386_/A _07386_/B vssd1 vssd1 vccd1 vccd1 _07386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ _09414_/B _09125_/B _09126_/B vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_72_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06337_ _06340_/B vssd1 vssd1 vccd1 vccd1 _06342_/A sky130_fd_sc_hd__inv_2
XFILLER_0_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _09056_/A vssd1 vssd1 vccd1 vccd1 _09057_/B sky130_fd_sc_hd__inv_2
X_06268_ _05796_/Y _06268_/B _06268_/C vssd1 vssd1 vccd1 vccd1 _06269_/B sky130_fd_sc_hd__nand3b_1
X_08007_ _09854_/B _09601_/B _09988_/A _09987_/A vssd1 vssd1 vccd1 vccd1 _08102_/A
+ sky130_fd_sc_hd__and4_1
X_05219_ _05219_/A _05219_/B _05219_/C vssd1 vssd1 vccd1 vccd1 _05338_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06199_ _06199_/A _06199_/B _06199_/C vssd1 vssd1 vccd1 vccd1 _06201_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09958_ _09967_/B _09967_/A vssd1 vssd1 vccd1 vccd1 _09958_/Y sky130_fd_sc_hd__nor2_1
X_08909_ _08907_/Y _09262_/B _08909_/C vssd1 vssd1 vccd1 vccd1 _09262_/A sky130_fd_sc_hd__nand3b_1
X_09889_ input54/X _10111_/B vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05942__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05389__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput82 hold63/A vssd1 vssd1 vccd1 vccd1 y_o[24] sky130_fd_sc_hd__buf_12
Xoutput71 _10494_/Q vssd1 vssd1 vccd1 vccd1 y_o[14] sky130_fd_sc_hd__buf_12
Xoutput93 _10485_/Q vssd1 vssd1 vccd1 vccd1 y_o[5] sky130_fd_sc_hd__buf_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09324__B _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _10029_/A _10029_/B vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05570_ _05981_/B _05981_/A vssd1 vssd1 vccd1 vccd1 _05571_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_85_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ _07188_/Y _07239_/Y _07187_/A vssd1 vssd1 vccd1 vccd1 _07475_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07171_ _07171_/A _07170_/A vssd1 vssd1 vccd1 vccd1 _07172_/B sky130_fd_sc_hd__or2b_1
X_06122_ _05605_/C _05605_/B _06121_/Y vssd1 vssd1 vccd1 vccd1 _06129_/B sky130_fd_sc_hd__a21oi_1
X_06053_ _06594_/B _06594_/A vssd1 vssd1 vccd1 vccd1 _06098_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09812_ _09814_/B vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09743_ _09745_/C vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06955_ _07008_/A _07007_/A vssd1 vssd1 vccd1 vccd1 _06955_/Y sky130_fd_sc_hd__nor2_1
X_09674_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__nand2_1
X_06886_ _06886_/A _06886_/B vssd1 vssd1 vccd1 vccd1 _07025_/C sky130_fd_sc_hd__nand2_1
X_05906_ _05906_/A _05906_/B _05906_/C vssd1 vssd1 vccd1 vccd1 _05907_/B sky130_fd_sc_hd__nand3_1
X_08625_ _08625_/A _08893_/A vssd1 vssd1 vccd1 vccd1 _08628_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07035__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05837_ _05948_/B vssd1 vssd1 vccd1 vccd1 _05947_/A sky130_fd_sc_hd__inv_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08556_/A vssd1 vssd1 vccd1 vccd1 _08557_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07507_ _07507_/A _07507_/B vssd1 vssd1 vccd1 vccd1 _07511_/B sky130_fd_sc_hd__nand2_1
X_05768_ _10026_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _05787_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08487_ _08279_/B _08279_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__o21a_1
X_05699_ _09548_/A input12/X vssd1 vssd1 vccd1 vccd1 _05706_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07438_ _10112_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07369_ _07369_/A _07369_/B vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__nand2_1
X_09108_ _09107_/B _09108_/B _09406_/B vssd1 vssd1 vccd1 vccd1 _09406_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ _10480_/Q hold43/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__or2_1
X_09039_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09042_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_60_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09596__A2 _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05847__B _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06740_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06749_/B sky130_fd_sc_hd__inv_2
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06671_ _06781_/A _06782_/A vssd1 vssd1 vccd1 vccd1 _06671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08410_ _08410_/A _08410_/B vssd1 vssd1 vccd1 vccd1 _08652_/A sky130_fd_sc_hd__nand2_1
X_05622_ _05629_/C vssd1 vssd1 vccd1 vccd1 _05626_/B sky130_fd_sc_hd__inv_2
X_09390_ input52/X vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__inv_2
XFILLER_0_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ _08341_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _08342_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05553_ _05562_/A _06043_/A vssd1 vssd1 vccd1 vccd1 _06087_/B sky130_fd_sc_hd__nand2_1
X_08272_ _09496_/B _08272_/B vssd1 vssd1 vccd1 vccd1 _08274_/B sky130_fd_sc_hd__nand2_1
X_05484_ _05478_/Y _05480_/Y _05485_/A vssd1 vssd1 vccd1 vccd1 _05487_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09220__D _09533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07223_ _07223_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07229_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08414__A _08651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ _07154_/A _07154_/B vssd1 vssd1 vccd1 vccd1 _07709_/A sky130_fd_sc_hd__nand2_2
X_06105_ _06402_/B _06105_/B vssd1 vssd1 vccd1 vccd1 _06183_/B sky130_fd_sc_hd__nand2_1
X_07085_ _07345_/A _07347_/A vssd1 vssd1 vccd1 vccd1 _07085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06036_ _06041_/A _06457_/A vssd1 vssd1 vccd1 vccd1 _06505_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07987_ _07989_/A _07989_/B vssd1 vssd1 vccd1 vccd1 _07988_/A sky130_fd_sc_hd__nand2_1
X_09726_ _09718_/Y _09719_/X _09727_/A vssd1 vssd1 vccd1 vccd1 _09730_/A sky130_fd_sc_hd__o21ai_1
X_06938_ _06938_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _07090_/B sky130_fd_sc_hd__nand2_1
X_09657_ _09661_/B _09683_/A vssd1 vssd1 vccd1 vccd1 _09660_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06869_ _07030_/B _07029_/A vssd1 vssd1 vccd1 vccd1 _07033_/C sky130_fd_sc_hd__nand2_1
X_09588_ _09588_/A _09589_/A _09845_/A vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__nand3_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08876_/C vssd1 vssd1 vccd1 vccd1 _08875_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08539_/A vssd1 vssd1 vccd1 vccd1 _08540_/C sky130_fd_sc_hd__inv_2
XFILLER_0_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _10509_/CLK hold8/X fanout100/X vssd1 vssd1 vccd1 vccd1 _10501_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__06109__A _09685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08324__A _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _10432_/A _10434_/A vssd1 vssd1 vccd1 vccd1 _10433_/A sky130_fd_sc_hd__and2_1
X_10363_ hold57/X vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__inv_2
XANTENNA__05667__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10294_ _10298_/A hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__xor2_1
XFILLER_0_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05858__A _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08890_ _08890_/A _08890_/B vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06689__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _08055_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07911_/A sky130_fd_sc_hd__nor2_1
X_07841_ _07841_/A _07841_/B vssd1 vssd1 vccd1 vccd1 _07841_/Y sky130_fd_sc_hd__nand2_1
X_07772_ _08866_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _07849_/B sky130_fd_sc_hd__nand2_1
X_09511_ _09829_/A _09511_/B _09511_/C vssd1 vssd1 vccd1 vccd1 _09515_/C sky130_fd_sc_hd__nand3_1
X_06723_ _09963_/A _09601_/B vssd1 vssd1 vccd1 vccd1 _06725_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09442_ _09443_/B _09443_/A vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__or2_1
XFILLER_0_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06654_ _06654_/A _06654_/B _06654_/C vssd1 vssd1 vccd1 vccd1 _06823_/C sky130_fd_sc_hd__nand3_1
X_09373_ _09076_/Y _09079_/B _09077_/A vssd1 vssd1 vccd1 vccd1 _09375_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09257__A1 _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05605_ _05605_/A _05605_/B _05605_/C vssd1 vssd1 vccd1 vccd1 _05606_/B sky130_fd_sc_hd__nand3_1
X_06585_ _06585_/A _06585_/B vssd1 vssd1 vccd1 vccd1 _06587_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ _08814_/B vssd1 vssd1 vccd1 vccd1 _10084_/D sky130_fd_sc_hd__inv_2
XFILLER_0_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05536_ _05540_/C vssd1 vssd1 vccd1 vccd1 _05537_/C sky130_fd_sc_hd__inv_2
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05467_ _09022_/C _08272_/B vssd1 vssd1 vccd1 vccd1 _05867_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08186_ _08186_/A _08186_/B _08186_/C vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05398_ _05398_/A vssd1 vssd1 vccd1 vccd1 _05399_/C sky130_fd_sc_hd__inv_2
X_07206_ _07206_/A _07206_/B vssd1 vssd1 vccd1 vccd1 _07207_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05768__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ _07137_/A _07137_/B vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__nand2_1
X_07068_ _09560_/B _08247_/B vssd1 vssd1 vccd1 vccd1 _07206_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06019_ _06019_/A _06019_/B _06019_/C vssd1 vssd1 vccd1 vccd1 _06021_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06111__B _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _10043_/A _10052_/A vssd1 vssd1 vccd1 vccd1 _09714_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08319__A _08319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07877__B _09953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ hold68/X vssd1 vssd1 vccd1 vccd1 _10502_/D sky130_fd_sc_hd__clkbuf_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ hold81/A _10277_/B vssd1 vssd1 vccd1 vccd1 _10299_/C sky130_fd_sc_hd__and2b_1
XANTENNA__09723__A2 _10051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__B2 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__A1 _09951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05860__B _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06370_ _06370_/A _06370_/B vssd1 vssd1 vccd1 vccd1 _06747_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06972__A _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05321_ input3/X vssd1 vssd1 vccd1 vccd1 _10043_/B sky130_fd_sc_hd__buf_6
XFILLER_0_71_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08040_ _08040_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _08042_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05252_ _05219_/C _05219_/B _05251_/Y vssd1 vssd1 vccd1 vccd1 _05285_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09991_ _09991_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08942_ _08942_/A _09297_/A vssd1 vssd1 vccd1 vccd1 _08947_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08873_ _08872_/B _08873_/B _09071_/A vssd1 vssd1 vccd1 vccd1 _09096_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07824_ _07741_/Y _07824_/B vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__nand2b_1
X_07755_ _07755_/A _07767_/A vssd1 vssd1 vccd1 vccd1 _07822_/B sky130_fd_sc_hd__nand2_1
X_07686_ _07695_/B _07695_/A vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__nor2_1
X_06706_ _06288_/Y _06705_/Y _06287_/A vssd1 vssd1 vccd1 vccd1 _06708_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09425_ _09427_/C vssd1 vssd1 vccd1 vccd1 _09426_/B sky130_fd_sc_hd__inv_2
XANTENNA__08139__A _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__A _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06637_ _06637_/A _06637_/B vssd1 vssd1 vccd1 vccd1 _06639_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ _09356_/A _09356_/B vssd1 vssd1 vccd1 vccd1 _09378_/A sky130_fd_sc_hd__nor2_1
X_06568_ _06570_/A _06571_/A vssd1 vssd1 vccd1 vccd1 _06569_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06882__A _09022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09287_ _09447_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08307_ _08307_/A _08307_/B vssd1 vssd1 vccd1 vccd1 _08309_/A sky130_fd_sc_hd__nand2_1
X_06499_ _06499_/A _06499_/B _08306_/B vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05519_ _05538_/B _05539_/C _05539_/B vssd1 vssd1 vccd1 vccd1 _06022_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08238_ _08238_/A _08239_/A vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08169_ _08169_/A _08169_/B _08175_/A vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__nand3_2
X_10200_ _10200_/A hold19/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__xor2_1
X_10131_ _10131_/A _10131_/B _10131_/C vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10062_ _10063_/B _10063_/A vssd1 vssd1 vccd1 vccd1 _10062_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10003__A2 _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10329_ _10329_/A hold6/X vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__and2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06032__A _07216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05870_ _05870_/A _05870_/B vssd1 vssd1 vccd1 vccd1 _05875_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06686__B _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _07571_/A _07571_/B _07540_/C vssd1 vssd1 vccd1 vccd1 _07573_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07471_ _07471_/A _07471_/B _07471_/C vssd1 vssd1 vccd1 vccd1 _07534_/C sky130_fd_sc_hd__nand3_1
X_09210_ input46/X _10051_/A _09720_/B _09560_/B vssd1 vssd1 vccd1 vccd1 _09210_/X
+ sky130_fd_sc_hd__and4_1
X_06422_ input16/X vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09141_ _09141_/A _09141_/B _09141_/C vssd1 vssd1 vccd1 vccd1 _09144_/B sky130_fd_sc_hd__nand3_1
X_06353_ _06353_/A vssd1 vssd1 vccd1 vccd1 _06355_/A sky130_fd_sc_hd__inv_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ input51/X _10111_/B vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05304_ _05559_/B _05309_/C vssd1 vssd1 vccd1 vccd1 _05308_/A sky130_fd_sc_hd__nand2_1
X_08023_ _08023_/A vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__inv_2
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06284_ _09963_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _06288_/B sky130_fd_sc_hd__nand2_1
X_05235_ _09816_/B _08689_/A vssd1 vssd1 vccd1 vccd1 _05311_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08422__A _08422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _09977_/B _09977_/C vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08141__B _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _08924_/B _08925_/B _09277_/B vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__nand3b_1
X_08856_ _09140_/A _09141_/A vssd1 vssd1 vccd1 vccd1 _08856_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06877__A _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07807_ _07807_/A _07807_/B vssd1 vssd1 vccd1 vccd1 _07925_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08787_ _08794_/A _08995_/A vssd1 vssd1 vccd1 vccd1 _09014_/B sky130_fd_sc_hd__nand2_1
X_05999_ _05515_/C _05515_/B _05998_/Y vssd1 vssd1 vccd1 vccd1 _06018_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07738_ _07741_/A _07741_/B vssd1 vssd1 vccd1 vccd1 _07824_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07669_ _07654_/Y _07640_/C _07655_/Y vssd1 vssd1 vccd1 vccd1 _07691_/A sky130_fd_sc_hd__a21oi_1
X_09408_ _09407_/B _09408_/B _09408_/C vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _09338_/B _09339_/B _09339_/C vssd1 vssd1 vccd1 vccd1 _09340_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10114_ input52/X _09854_/B input53/X _09601_/B vssd1 vssd1 vccd1 vccd1 _10115_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10045_ _09199_/A _09684_/B _09548_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _10046_/B
+ sky130_fd_sc_hd__a22o_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09313__D _09313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06027__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05585__B _08780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _09960_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _07097_/B sky130_fd_sc_hd__nand2_1
X_09690_ _09690_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09696_/C sky130_fd_sc_hd__nand2_1
X_08710_ _09962_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _08711_/B sky130_fd_sc_hd__nand2_1
X_05922_ _05924_/C vssd1 vssd1 vccd1 vccd1 _05923_/B sky130_fd_sc_hd__inv_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09550__B1 _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ _09166_/B _08641_/B vssd1 vssd1 vccd1 vccd1 _08645_/B sky130_fd_sc_hd__nand2_1
X_05853_ _05924_/B _05924_/C _05852_/Y vssd1 vssd1 vccd1 vccd1 _05960_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__07156__A2 _07709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ _08572_/A _08572_/B vssd1 vssd1 vccd1 vccd1 _08574_/A sky130_fd_sc_hd__nand2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05784_ _05784_/A _05784_/B vssd1 vssd1 vccd1 vccd1 _05786_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07523_ _07524_/B _07523_/B _07523_/C vssd1 vssd1 vccd1 vccd1 _07898_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10490__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ _07454_/A _07454_/B vssd1 vssd1 vccd1 vccd1 _07463_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06405_ _06406_/B _06406_/A vssd1 vssd1 vccd1 vccd1 _06405_/Y sky130_fd_sc_hd__nand2_1
X_07385_ _07386_/B _07386_/A vssd1 vssd1 vccd1 vccd1 _07385_/Y sky130_fd_sc_hd__nand2_1
X_09124_ _09124_/A _09124_/B vssd1 vssd1 vccd1 vccd1 _09126_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06336_ _06739_/B _06739_/C vssd1 vssd1 vccd1 vccd1 _06744_/A sky130_fd_sc_hd__nand2_1
X_09055_ _09055_/A _09055_/B vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__nor2_1
X_06267_ _05796_/Y _06266_/Y _05795_/A vssd1 vssd1 vccd1 vccd1 _06269_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08006_ _08103_/A vssd1 vssd1 vccd1 vccd1 _08006_/Y sky130_fd_sc_hd__inv_2
X_05218_ _05251_/A _05251_/B vssd1 vssd1 vccd1 vccd1 _05219_/C sky130_fd_sc_hd__nand2_1
X_06198_ _06399_/A _06198_/B _06198_/C vssd1 vssd1 vccd1 vccd1 _06199_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07991__A _08337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _09262_/B _08909_/C _08907_/Y vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__a21bo_1
X_09888_ _09631_/B input54/X _10126_/B _09629_/X vssd1 vssd1 vccd1 vccd1 _10109_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08839_/A _08839_/B vssd1 vssd1 vccd1 vccd1 _08839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10507__RESET_B fanout99/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput83 hold49/A vssd1 vssd1 vccd1 vccd1 y_o[25] sky130_fd_sc_hd__buf_12
Xoutput72 _10495_/Q vssd1 vssd1 vccd1 vccd1 y_o[15] sky130_fd_sc_hd__buf_12
Xoutput94 _10486_/Q vssd1 vssd1 vccd1 vccd1 y_o[6] sky130_fd_sc_hd__buf_12
XFILLER_0_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10028_ _09528_/A _09816_/B _09685_/A _09496_/B vssd1 vssd1 vccd1 vccd1 _10029_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09324__C _09816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08099__B1 _10112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07170_ _07170_/A _07171_/A vssd1 vssd1 vccd1 vccd1 _07172_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06121_ _06121_/A _06121_/B vssd1 vssd1 vccd1 vccd1 _06121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06052_ _05571_/C _05571_/B _05981_/Y vssd1 vssd1 vccd1 vccd1 _06594_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09814_/B sky130_fd_sc_hd__nand2_1
X_09742_ _09742_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09745_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06954_ _07011_/C vssd1 vssd1 vccd1 vccd1 _07010_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09673_ _09675_/B _09941_/B vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__nand2_1
X_06885_ _06885_/A _06885_/B _06885_/C vssd1 vssd1 vccd1 vccd1 _06886_/B sky130_fd_sc_hd__nand3_1
X_05905_ _05905_/A _05905_/B vssd1 vssd1 vccd1 vccd1 _05907_/A sky130_fd_sc_hd__nand2_1
X_08624_ _08623_/B _08624_/B _08886_/C vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__07035__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05836_ _05948_/B _05947_/B vssd1 vssd1 vccd1 vccd1 _05918_/C sky130_fd_sc_hd__nand2_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08555_ _08551_/Y _08553_/Y _08556_/A vssd1 vssd1 vccd1 vccd1 _08558_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05767_ _05787_/A _05787_/B vssd1 vssd1 vccd1 vccd1 _05770_/A sky130_fd_sc_hd__nand2_1
X_07506_ _07508_/C vssd1 vssd1 vccd1 vccd1 _07507_/B sky130_fd_sc_hd__inv_2
X_05698_ input43/X vssd1 vssd1 vccd1 vccd1 _09548_/A sky130_fd_sc_hd__buf_4
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08486_ _08490_/B _08737_/A vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07437_ _07437_/A _07437_/B vssd1 vssd1 vccd1 vccd1 _07442_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07368_ _07370_/C vssd1 vssd1 vccd1 vccd1 _07369_/B sky130_fd_sc_hd__inv_2
X_09107_ _09107_/A _09107_/B vssd1 vssd1 vccd1 vccd1 _09115_/B sky130_fd_sc_hd__nand2_1
X_06319_ _06321_/A _06321_/B vssd1 vssd1 vccd1 vccd1 _06320_/A sky130_fd_sc_hd__nand2_1
X_07299_ _07299_/A _07299_/B vssd1 vssd1 vccd1 vccd1 _07321_/A sky130_fd_sc_hd__nor2_1
X_09038_ _09358_/A _09038_/B vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_99_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__A3 _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10470__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06670_ _06774_/C _06774_/B _06669_/Y vssd1 vssd1 vccd1 vccd1 _06782_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05621_ _05621_/A _05621_/B vssd1 vssd1 vccd1 vccd1 _05629_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08340_ _08340_/A vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__inv_2
X_05552_ _06043_/B _05552_/B _05552_/C vssd1 vssd1 vccd1 vccd1 _06043_/A sky130_fd_sc_hd__nand3_2
X_08271_ input6/X _09313_/D vssd1 vssd1 vccd1 vccd1 _08274_/A sky130_fd_sc_hd__nand2_1
X_05483_ _09960_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _05485_/A sky130_fd_sc_hd__nand2_1
X_07222_ _07222_/A _07222_/B _07222_/C vssd1 vssd1 vccd1 vccd1 _07223_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_42_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07153_ _07153_/A _07153_/B vssd1 vssd1 vccd1 vccd1 _07154_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06104_ _05626_/C _05626_/B _05979_/Y vssd1 vssd1 vccd1 vccd1 _06105_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07084_ _07350_/C vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__inv_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06035_ _06034_/B _06457_/B _06035_/C vssd1 vssd1 vccd1 vccd1 _06457_/A sky130_fd_sc_hd__nand3b_2
X_07986_ _07986_/A _07986_/B _07986_/C vssd1 vssd1 vccd1 vccd1 _08087_/B sky130_fd_sc_hd__nand3_2
X_09725_ _09725_/A _09725_/B vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__xor2_1
X_06937_ _06937_/A _06937_/B vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__nand2_1
X_09656_ _09656_/A _09683_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_96_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ input49/X input50/X _08862_/B _08866_/B vssd1 vssd1 vccd1 vccd1 _08876_/C
+ sky130_fd_sc_hd__and4_1
X_06868_ input5/X _08422_/A vssd1 vssd1 vccd1 vccd1 _07029_/A sky130_fd_sc_hd__nand2_1
X_09587_ _09587_/A _09587_/B _09845_/B vssd1 vssd1 vccd1 vccd1 _09845_/A sky130_fd_sc_hd__nand3_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05819_ _08866_/B vssd1 vssd1 vccd1 vccd1 _10126_/B sky130_fd_sc_hd__clkbuf_8
X_06799_ _06842_/A _06841_/A vssd1 vssd1 vccd1 vccd1 _06799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A _08539_/A vssd1 vssd1 vccd1 vccd1 _08547_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08469_ _08469_/A _08470_/A vssd1 vssd1 vccd1 vccd1 _08476_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ _10511_/CLK _10500_/D fanout100/X vssd1 vssd1 vccd1 vccd1 _10500_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__06109__B _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ _10431_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__nand2_1
X_10362_ hold62/X vssd1 vssd1 vccd1 vccd1 _10506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10293_ _10293_/A hold28/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05204__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06689__B _09361_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _07841_/A _07841_/B vssd1 vssd1 vccd1 vccd1 _07842_/A sky130_fd_sc_hd__nor2_1
X_07771_ _07789_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07806_/A sky130_fd_sc_hd__nand2_1
X_09510_ _09510_/A _09510_/B vssd1 vssd1 vccd1 vccd1 _09515_/B sky130_fd_sc_hd__nand2_1
X_06722_ _09962_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _06725_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09081__A _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _09789_/B _09441_/B vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__nand2_1
X_06653_ _06653_/A _06653_/B vssd1 vssd1 vccd1 vccd1 _06823_/B sky130_fd_sc_hd__nand2_1
X_09372_ _09372_/A _09372_/B vssd1 vssd1 vccd1 vccd1 _09375_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05604_ _05604_/A vssd1 vssd1 vccd1 vccd1 _05605_/B sky130_fd_sc_hd__inv_2
X_06584_ _06590_/A _06590_/B vssd1 vssd1 vccd1 vccd1 _06589_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08323_ _10043_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05535_ _05535_/A _05535_/B vssd1 vssd1 vccd1 vccd1 _05540_/C sky130_fd_sc_hd__nand2_1
X_08254_ _08464_/A _08258_/C vssd1 vssd1 vccd1 vccd1 _08504_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05466_ _09022_/D _09313_/D vssd1 vssd1 vccd1 vccd1 _05866_/A sky130_fd_sc_hd__nand2_1
X_08185_ _08153_/A _08153_/B _08184_/Y vssd1 vssd1 vccd1 vccd1 _08186_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_6_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05397_ _05397_/A _05405_/A _05397_/C vssd1 vssd1 vccd1 vccd1 _05399_/B sky130_fd_sc_hd__nand3_1
X_07205_ _07205_/A _07205_/B vssd1 vssd1 vccd1 vccd1 _07207_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05768__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07136_ _07138_/A vssd1 vssd1 vccd1 vccd1 _07137_/B sky130_fd_sc_hd__inv_2
X_07067_ _07088_/B _07088_/A vssd1 vssd1 vccd1 vccd1 _07078_/B sky130_fd_sc_hd__nand2_1
X_06018_ _06018_/A _06018_/B _06018_/C vssd1 vssd1 vccd1 vccd1 _06019_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09256__A _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _09733_/A _09733_/C vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__nand2_1
X_07969_ _09392_/C _09777_/A _07859_/C vssd1 vssd1 vccd1 vccd1 _07970_/B sky130_fd_sc_hd__o21ai_1
X_09639_ _09917_/A _09645_/C vssd1 vssd1 vccd1 vccd1 _09931_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08335__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ _10414_/A _10416_/A vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__and2_1
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ hold67/X _10349_/A vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__and2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _10493_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _10277_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09487__A2 _09485_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05320_ _05320_/A _05320_/B vssd1 vssd1 vccd1 vccd1 _05376_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06972__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05251_ _05251_/A _05251_/B vssd1 vssd1 vccd1 vccd1 _05251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09990_ _09990_/A _09990_/B vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_86_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08941_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _09297_/A sky130_fd_sc_hd__nand2_1
X_08872_ _08872_/A _08872_/B vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09804__A _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ _07823_/A _07823_/B vssd1 vssd1 vccd1 vccd1 _07865_/A sky130_fd_sc_hd__nand2_1
X_07754_ _07767_/B _07754_/B _07754_/C vssd1 vssd1 vccd1 vccd1 _07767_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_79_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07685_ _07692_/B _07692_/C vssd1 vssd1 vccd1 vccd1 _07695_/A sky130_fd_sc_hd__nand2_1
X_06705_ _06707_/C vssd1 vssd1 vccd1 vccd1 _06705_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09424_ _09424_/A _09424_/B vssd1 vssd1 vccd1 vccd1 _09427_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08139__B _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__B _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06636_ _08656_/A _06638_/C vssd1 vssd1 vccd1 vccd1 _06637_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09355_ _09412_/B _09658_/B vssd1 vssd1 vccd1 vccd1 _09410_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06567_ _06572_/C vssd1 vssd1 vccd1 vccd1 _06569_/B sky130_fd_sc_hd__inv_2
XANTENNA__06882__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ _09286_/A _09286_/B vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__nand2_1
X_08306_ _08306_/A _08306_/B vssd1 vssd1 vccd1 vccd1 _08307_/B sky130_fd_sc_hd__nand2_1
X_06498_ _06501_/A _06500_/B _08281_/A vssd1 vssd1 vccd1 vccd1 _08306_/B sky130_fd_sc_hd__nand3_1
X_05518_ _05518_/A _05518_/B _05518_/C vssd1 vssd1 vccd1 vccd1 _05539_/B sky130_fd_sc_hd__nand3_1
X_08237_ _08237_/A _08237_/B vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__xor2_1
X_05449_ _05449_/A _05449_/B vssd1 vssd1 vccd1 vccd1 _05454_/C sky130_fd_sc_hd__nand2_1
X_08168_ _08168_/A _08168_/B vssd1 vssd1 vccd1 vccd1 _08170_/A sky130_fd_sc_hd__nand2_1
X_08099_ _09601_/B _09988_/A _10112_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _08100_/B
+ sky130_fd_sc_hd__a22o_1
X_07119_ _07119_/A _07119_/B vssd1 vssd1 vccd1 vccd1 _07121_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10061_ _10067_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _10066_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10328_ _10500_/Q hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__nand2_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ hold103/X vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__inv_2
XFILLER_0_56_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07470_ _07470_/A _07470_/B vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__nand2_1
X_06421_ _06426_/A vssd1 vssd1 vccd1 vccd1 _06425_/A sky130_fd_sc_hd__inv_2
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09140_ _09140_/A _09140_/B vssd1 vssd1 vccd1 vccd1 _09144_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06352_ _06749_/A _06750_/A vssd1 vssd1 vccd1 vccd1 _06742_/B sky130_fd_sc_hd__nand2_1
X_09071_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09090_/B sky130_fd_sc_hd__and2_1
X_06283_ _09361_/C vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05303_ _05303_/A _05303_/B vssd1 vssd1 vccd1 vccd1 _05309_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08022_ _08031_/B vssd1 vssd1 vccd1 vccd1 _08029_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05234_ input58/X vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__buf_8
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09973_ _09973_/A _09973_/B _09973_/C vssd1 vssd1 vccd1 vccd1 _09977_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08924_ _08924_/A _08924_/B vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07038__B _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _08853_/Y _08593_/B _08854_/Y vssd1 vssd1 vccd1 vccd1 _09141_/A sky130_fd_sc_hd__a21oi_4
X_08786_ _08785_/B _08995_/B _08786_/C vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__nand3b_1
X_07806_ _07806_/A _07806_/B vssd1 vssd1 vccd1 vccd1 _07807_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06877__B _08689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ _08810_/B input33/X vssd1 vssd1 vccd1 vccd1 _07741_/B sky130_fd_sc_hd__nand2_1
X_05998_ _05998_/A _05998_/B vssd1 vssd1 vccd1 vccd1 _05998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07668_ _07668_/A _07668_/B vssd1 vssd1 vccd1 vccd1 _07691_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09407_ _09407_/A _09407_/B vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__nand2_1
X_06619_ _08655_/A _08413_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _06635_/A sky130_fd_sc_hd__nand3_2
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07602_/B sky130_fd_sc_hd__nand2_1
X_09338_ _09338_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _09340_/A sky130_fd_sc_hd__nand2_1
X_09269_ _09981_/B input17/X vssd1 vssd1 vccd1 vccd1 _09270_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09709__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10113_ _10113_/A _10113_/B _10113_/C _10113_/D vssd1 vssd1 vccd1 vccd1 _10115_/A
+ sky130_fd_sc_hd__or4_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
X_10044_ _10044_/A _10044_/B _10044_/C _10044_/D vssd1 vssd1 vccd1 vccd1 _10046_/A
+ sky130_fd_sc_hd__or4_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06027__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ _09528_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _07399_/B sky130_fd_sc_hd__nand2_1
X_05921_ _05924_/A _05924_/B vssd1 vssd1 vccd1 vccd1 _05923_/A sky130_fd_sc_hd__nand2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09550__A1 _09199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__B2 _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ _09166_/A vssd1 vssd1 vccd1 vccd1 _08641_/B sky130_fd_sc_hd__inv_2
X_05852_ _05852_/A _05852_/B vssd1 vssd1 vccd1 vccd1 _05852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08571_ _08571_/A _08870_/A vssd1 vssd1 vccd1 vccd1 _08572_/B sky130_fd_sc_hd__nand2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05783_ _05785_/C vssd1 vssd1 vccd1 vccd1 _05784_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07522_ _07609_/B _07610_/B vssd1 vssd1 vccd1 vccd1 _07523_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07453_ _07453_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07454_/A sky130_fd_sc_hd__nand2_1
X_06404_ _06404_/A _06404_/B vssd1 vssd1 vccd1 vccd1 _06599_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09123_ _08851_/C _08851_/B _08899_/B vssd1 vssd1 vccd1 vccd1 _09124_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07384_ _07643_/A vssd1 vssd1 vccd1 vccd1 _07406_/A sky130_fd_sc_hd__inv_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06335_ _06335_/A _06335_/B _06335_/C vssd1 vssd1 vccd1 vccd1 _06739_/C sky130_fd_sc_hd__nand3_1
X_09054_ _09060_/A _09060_/B vssd1 vssd1 vccd1 vccd1 _09059_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06266_ _06268_/C vssd1 vssd1 vccd1 vccd1 _06266_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08005_ _10112_/B _09986_/A vssd1 vssd1 vccd1 vccd1 _08103_/A sky130_fd_sc_hd__nand2_1
X_05217_ _05217_/A vssd1 vssd1 vccd1 vccd1 _05219_/B sky130_fd_sc_hd__inv_2
XANTENNA__07049__A _09022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06197_ _06399_/B _06197_/B vssd1 vssd1 vccd1 vccd1 _06199_/A sky130_fd_sc_hd__nand2_1
X_09956_ _09956_/A _09956_/B vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__xor2_1
X_09887_ input56/X _10126_/B vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__nand2_1
X_08907_ _09986_/A input18/X vssd1 vssd1 vccd1 vccd1 _08907_/Y sky130_fd_sc_hd__nand2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05792__A _09963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08838_ _08839_/B _08839_/A vssd1 vssd1 vccd1 vccd1 _08838_/Y sky130_fd_sc_hd__nand2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08769_ _08901_/A _08769_/B vssd1 vssd1 vccd1 vccd1 _08770_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput84 hold60/A vssd1 vssd1 vccd1 vccd1 y_o[26] sky130_fd_sc_hd__buf_12
Xoutput73 _10496_/Q vssd1 vssd1 vccd1 vccd1 y_o[16] sky130_fd_sc_hd__buf_12
Xoutput95 _10487_/Q vssd1 vssd1 vccd1 vccd1 y_o[7] sky130_fd_sc_hd__buf_12
X_10027_ _10027_/A _10027_/B _10027_/C _10027_/D vssd1 vssd1 vccd1 vccd1 _10029_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__09324__D _09496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05207__A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__B2 _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__A1 _09601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09599__B2 _09854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09599__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06120_ _06129_/A _06534_/A vssd1 vssd1 vccd1 vccd1 _06128_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06051_ _06100_/B _06100_/C vssd1 vssd1 vccd1 vccd1 _06594_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ _09957_/A _09814_/C vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__nand2_1
X_09741_ _09741_/A vssd1 vssd1 vccd1 vccd1 _09742_/B sky130_fd_sc_hd__inv_2
X_06953_ _06953_/A _06953_/B vssd1 vssd1 vccd1 vccd1 _07011_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05904_ _05906_/A _05906_/B vssd1 vssd1 vccd1 vccd1 _05905_/A sky130_fd_sc_hd__nand2_1
X_09672_ _09672_/A _09672_/B _09682_/A vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__nand3_2
X_06884_ _06884_/A vssd1 vssd1 vccd1 vccd1 _06885_/B sky130_fd_sc_hd__inv_2
X_08623_ _08623_/A _08623_/B vssd1 vssd1 vccd1 vccd1 _08625_/A sky130_fd_sc_hd__nand2_1
X_05835_ input6/X _08689_/A vssd1 vssd1 vccd1 vccd1 _05947_/B sky130_fd_sc_hd__nand2_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08554_ _10043_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__nand2_1
X_05766_ _05765_/B _05766_/B vssd1 vssd1 vccd1 vccd1 _05787_/B sky130_fd_sc_hd__nand2b_1
X_07505_ _07542_/A _07539_/A vssd1 vssd1 vccd1 vccd1 _07505_/Y sky130_fd_sc_hd__nand2_1
X_08485_ _08737_/B _08485_/B _08485_/C vssd1 vssd1 vccd1 vccd1 _08737_/A sky130_fd_sc_hd__nand3_1
X_05697_ _05729_/A _05729_/B vssd1 vssd1 vccd1 vccd1 _05728_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _07440_/B vssd1 vssd1 vccd1 vccd1 _07437_/B sky130_fd_sc_hd__inv_2
X_07367_ _07365_/Y _07312_/B _07366_/Y vssd1 vssd1 vccd1 vccd1 _07370_/C sky130_fd_sc_hd__a21oi_1
X_09106_ input52/X _10126_/B vssd1 vssd1 vccd1 vccd1 _09107_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06318_ _06318_/A _06318_/B vssd1 vssd1 vccd1 vccd1 _06321_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ _09037_/A vssd1 vssd1 vccd1 vccd1 _09038_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07298_ _07298_/A vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__inv_2
XFILLER_0_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06249_ _06695_/A _06696_/B vssd1 vssd1 vccd1 vccd1 _06699_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09211__B1 _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09942_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09722__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10469__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05620_ _05620_/A _05620_/B _05620_/C vssd1 vssd1 vccd1 vccd1 _05621_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_86_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08248__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05551_ _05551_/A vssd1 vssd1 vccd1 vccd1 _05552_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _08313_/A _08314_/B vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__nand2_1
X_05482_ input28/X vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__buf_6
X_07221_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07222_/C sky130_fd_sc_hd__inv_2
XFILLER_0_89_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07152_ _07707_/B _07710_/B _07706_/B vssd1 vssd1 vccd1 vccd1 _10428_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06103_ _06404_/A _06103_/B vssd1 vssd1 vccd1 vccd1 _06402_/B sky130_fd_sc_hd__nand2_1
X_07083_ _07092_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07350_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06034_ _06034_/A _06034_/B vssd1 vssd1 vccd1 vccd1 _06041_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07985_ _08091_/B vssd1 vssd1 vccd1 vccd1 _07986_/B sky130_fd_sc_hd__inv_2
X_09724_ _09724_/A _09723_/X vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__or2b_1
X_06936_ _06936_/A _06936_/B vssd1 vssd1 vccd1 vccd1 _06937_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _09655_/A vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__inv_2
X_06867_ input4/X input44/X vssd1 vssd1 vccd1 vccd1 _07030_/B sky130_fd_sc_hd__nand2_2
X_05818_ _08862_/B vssd1 vssd1 vccd1 vccd1 _10111_/B sky130_fd_sc_hd__buf_4
X_08606_ _08628_/A vssd1 vssd1 vccd1 vccd1 _08627_/A sky130_fd_sc_hd__inv_2
X_09586_ _09586_/A vssd1 vssd1 vccd1 vccd1 _09587_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ _06843_/C vssd1 vssd1 vccd1 vccd1 _06834_/C sky130_fd_sc_hd__inv_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08537_ _08537_/A _08537_/B vssd1 vssd1 vccd1 vccd1 _08539_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05749_ _05749_/A _05749_/B _05749_/C vssd1 vssd1 vccd1 vccd1 _05886_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08468_ _08468_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _08470_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07997__A _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ _07419_/A _07419_/B vssd1 vssd1 vccd1 vccd1 _07610_/B sky130_fd_sc_hd__nand2_1
X_08399_ _08399_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__and2_1
XFILLER_0_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ _10431_/B _10431_/A vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__or2_1
X_10361_ hold61/X _10365_/A vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__and2_1
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ _10290_/Y hold114/A vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09499__B1 _09962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05204__B _08420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07770_ _07770_/A _07770_/B _07770_/C vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__nand3_2
X_06721_ _09960_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _06937_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09440_ _10000_/A _09998_/B _09999_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _09441_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06652_ _06654_/B _06654_/C vssd1 vssd1 vccd1 vccd1 _06653_/A sky130_fd_sc_hd__nand2_1
X_09371_ _09372_/B _09372_/A vssd1 vssd1 vccd1 vccd1 _09375_/A sky130_fd_sc_hd__or2_1
X_05603_ _05603_/A _05604_/A vssd1 vssd1 vccd1 vccd1 _05606_/A sky130_fd_sc_hd__nand2_1
X_06583_ _06583_/A _06583_/B _06583_/C vssd1 vssd1 vccd1 vccd1 _06590_/B sky130_fd_sc_hd__nand3_1
X_08322_ _08322_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08332_/B sky130_fd_sc_hd__and2_1
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05534_ _05534_/A _05534_/B _05534_/C vssd1 vssd1 vccd1 vccd1 _05535_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08706__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08258_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07204_ _07169_/C _07169_/B _07165_/Y vssd1 vssd1 vccd1 vccd1 _07208_/A sky130_fd_sc_hd__a21o_1
X_05465_ _05826_/A _05826_/B vssd1 vssd1 vccd1 vccd1 _05825_/A sky130_fd_sc_hd__nand2_1
X_08184_ _08184_/A _08184_/B vssd1 vssd1 vccd1 vccd1 _08184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06226__A _09684_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05396_ _05405_/B _05396_/B vssd1 vssd1 vccd1 vccd1 _05399_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07135_ _07132_/Y _07666_/B _07134_/Y vssd1 vssd1 vccd1 vccd1 _07684_/B sky130_fd_sc_hd__a21oi_1
X_07066_ _07080_/A _07080_/B vssd1 vssd1 vccd1 vccd1 _07088_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06017_ _06017_/A _06017_/B vssd1 vssd1 vccd1 vccd1 _06019_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09256__B _09987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _08023_/A _08024_/A vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__nand2_1
X_09707_ _09705_/A _09705_/B _09701_/Y vssd1 vssd1 vccd1 vccd1 _09733_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06919_ _07111_/B _07110_/B vssd1 vssd1 vccd1 vccd1 _07109_/C sky130_fd_sc_hd__nand2_1
X_07899_ _07899_/A _07899_/B vssd1 vssd1 vccd1 vccd1 _07903_/C sky130_fd_sc_hd__nand2_1
X_09638_ _09638_/A _09638_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09645_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10460__CLK _10494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _09569_/A _09569_/B vssd1 vssd1 vccd1 vccd1 _09572_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05305__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10413_ _10413_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10416_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10344_ _10344_/A hold66/X vssd1 vssd1 vccd1 vccd1 _10349_/A sky130_fd_sc_hd__nand2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10275_ _10493_/Q hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05250_ _05291_/B _05291_/C _05249_/Y vssd1 vssd1 vccd1 vccd1 _05500_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08940_ _08941_/B _08941_/A vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__or2_1
X_08871_ _08569_/B _08870_/Y _08567_/Y vssd1 vssd1 vccd1 vccd1 _08872_/B sky130_fd_sc_hd__a21oi_1
X_07822_ _07822_/A _07822_/B vssd1 vssd1 vccd1 vccd1 _07823_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10483__CLK _10495_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _07753_/A vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__inv_2
X_07684_ _07684_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07692_/C sky130_fd_sc_hd__nand2_1
X_06704_ _06946_/A _06946_/B vssd1 vssd1 vccd1 vccd1 _06710_/A sky130_fd_sc_hd__nand2_1
X_09423_ _09137_/A _09137_/B _09134_/C vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__a21o_1
X_06635_ _06635_/A _06635_/B _06635_/C vssd1 vssd1 vccd1 vccd1 _06638_/C sky130_fd_sc_hd__nand3_1
X_09354_ _09353_/B _09433_/A _09354_/C vssd1 vssd1 vccd1 vccd1 _09658_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06566_ _06566_/A _06566_/B vssd1 vssd1 vccd1 vccd1 _06572_/C sky130_fd_sc_hd__xor2_1
X_08305_ _08308_/B _08308_/C vssd1 vssd1 vccd1 vccd1 _08307_/A sky130_fd_sc_hd__nand2_1
X_09285_ _09286_/B _09286_/A vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__or2_1
X_06497_ _06501_/C vssd1 vssd1 vccd1 vccd1 _06500_/B sky130_fd_sc_hd__inv_2
X_05517_ _05517_/A _05998_/B vssd1 vssd1 vccd1 vccd1 _05518_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08236_ _08236_/A _08236_/B vssd1 vssd1 vccd1 vccd1 _08237_/B sky130_fd_sc_hd__nand2_1
X_05448_ _05448_/A _05448_/B _05448_/C vssd1 vssd1 vccd1 vccd1 _05449_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07994__B _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ _08169_/A vssd1 vssd1 vccd1 vccd1 _08168_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09267__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05379_ _05380_/A _05380_/B vssd1 vssd1 vccd1 vccd1 _05379_/Y sky130_fd_sc_hd__nand2_1
X_07118_ _07363_/C _07356_/A vssd1 vssd1 vccd1 vccd1 _07119_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08098_ _09601_/B _10112_/B _09988_/A _09987_/A vssd1 vssd1 vccd1 vccd1 _08098_/X
+ sky130_fd_sc_hd__and4_1
X_07049_ _09022_/D _07960_/B vssd1 vssd1 vccd1 vccd1 _07052_/A sky130_fd_sc_hd__nand2_1
X_10060_ _10060_/A _10060_/B _10060_/C vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10327_ _10500_/Q hold5/X vssd1 vssd1 vccd1 vccd1 _10329_/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _10491_/Q hold102/X vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__nand2_1
X_10189_ _10482_/Q hold17/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07425__A _08814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06420_ _08420_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _06426_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06351_ _06759_/C _06759_/B _06350_/Y vssd1 vssd1 vccd1 vccd1 _06750_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09070_ _08832_/C _08832_/B _08819_/A vssd1 vssd1 vccd1 vccd1 _09091_/A sky130_fd_sc_hd__a21o_1
X_05302_ _05302_/A _05302_/B vssd1 vssd1 vccd1 vccd1 _05559_/B sky130_fd_sc_hd__nand2_1
X_06282_ _09962_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _06288_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08021_ _08114_/B _08019_/Y _08020_/Y vssd1 vssd1 vccd1 vccd1 _08031_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05233_ input8/X vssd1 vssd1 vccd1 vccd1 _09816_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09972_ _09790_/A _09971_/Y _09949_/Y vssd1 vssd1 vccd1 vccd1 _09973_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__10026__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ _08923_/A _09291_/A vssd1 vssd1 vccd1 vccd1 _08924_/B sky130_fd_sc_hd__nand2_1
X_08854_ _08854_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _08854_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08785_ _08785_/A _08785_/B vssd1 vssd1 vccd1 vccd1 _08794_/A sky130_fd_sc_hd__nand2_1
X_05997_ _06018_/A _06018_/C vssd1 vssd1 vccd1 vccd1 _06017_/A sky130_fd_sc_hd__nand2_1
X_07805_ _07805_/A _07893_/A _07893_/B vssd1 vssd1 vccd1 vccd1 _08055_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07736_ _08814_/B input44/X vssd1 vssd1 vccd1 vccd1 _07741_/A sky130_fd_sc_hd__nand2_1
X_07667_ _07667_/A _07667_/B _07667_/C vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nand3_1
X_09406_ _09406_/A _09406_/B vssd1 vssd1 vccd1 vccd1 _09407_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06618_ _06618_/A _06618_/B _06618_/C vssd1 vssd1 vccd1 vccd1 _06620_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07598_ _07598_/A _07788_/A vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__nand2_1
X_09337_ _09337_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09338_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06549_ _06549_/A _06549_/B vssd1 vssd1 vccd1 vccd1 _06554_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07070__A _08810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ input18/X vssd1 vssd1 vccd1 vccd1 _09270_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08219_ _08219_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08220_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09709__B _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ _09199_/A _09548_/A _10052_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _09200_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10112_ input54/X _10112_/B vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10043_ _10043_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _10047_/A sky130_fd_sc_hd__nand2_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09953__D_N _09775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ _05920_/A _05920_/B _05920_/C vssd1 vssd1 vccd1 vccd1 _05924_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09550__A2 _10043_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05851_ _06366_/C _05851_/B vssd1 vssd1 vccd1 vccd1 _05924_/C sky130_fd_sc_hd__nand2_1
X_08570_ _08870_/A _08571_/A vssd1 vssd1 vccd1 vccd1 _08572_/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07521_ _07536_/B _07516_/Y _07517_/Y vssd1 vssd1 vccd1 vccd1 _07609_/B sky130_fd_sc_hd__a21oi_1
X_05782_ _06187_/A _05782_/B vssd1 vssd1 vccd1 vccd1 _05785_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_9_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07452_ _07452_/A _07453_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07520_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06403_ _06401_/Y _06182_/B _06402_/Y vssd1 vssd1 vccd1 vccd1 _06616_/B sky130_fd_sc_hd__a21o_1
X_07383_ _07527_/B _07526_/B _07525_/A vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _09122_/A _09352_/A vssd1 vssd1 vccd1 vccd1 _09124_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06334_ _06334_/A _06334_/B _06334_/C vssd1 vssd1 vccd1 vccd1 _06335_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09053_ _09053_/A _09053_/B _09399_/A vssd1 vssd1 vccd1 vccd1 _09060_/B sky130_fd_sc_hd__nand3_1
X_06265_ _06658_/A _06658_/B vssd1 vssd1 vccd1 vccd1 _06271_/A sky130_fd_sc_hd__nand2_1
X_08004_ _09854_/B _09988_/A _09601_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _08004_/X
+ sky130_fd_sc_hd__a22o_1
X_05216_ _05216_/A _05216_/B vssd1 vssd1 vccd1 vccd1 _05219_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06234__A _10052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06196_ _06196_/A _06196_/B _06196_/C vssd1 vssd1 vccd1 vccd1 _06201_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__B _07960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09955_ _09955_/A _09955_/B vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__nand2_1
X_09886_ _09908_/A _09908_/C vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__nand2_1
X_08906_ _09751_/A _09762_/B _08904_/C vssd1 vssd1 vccd1 vccd1 _08909_/C sky130_fd_sc_hd__o21ai_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05792__B _08825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ _09056_/A _08843_/C vssd1 vssd1 vccd1 vccd1 _09111_/B sky130_fd_sc_hd__nand2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08471_/B _08471_/C _08673_/B vssd1 vssd1 vccd1 vccd1 _08770_/A sky130_fd_sc_hd__a21boi_1
X_08699_ _08703_/B _08927_/A vssd1 vssd1 vccd1 vccd1 _08702_/A sky130_fd_sc_hd__nand2_1
X_07719_ _07719_/A _07719_/B vssd1 vssd1 vccd1 vccd1 _07722_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06409__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 hold57/A vssd1 vssd1 vccd1 vccd1 y_o[27] sky130_fd_sc_hd__buf_12
Xoutput74 _10497_/Q vssd1 vssd1 vccd1 vccd1 y_o[17] sky130_fd_sc_hd__buf_12
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput96 _10488_/Q vssd1 vssd1 vccd1 vccd1 y_o[8] sky130_fd_sc_hd__buf_12
XFILLER_0_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10026_ _10026_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _10030_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08099__A2 _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09599__A2 _10083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06050_ _06099_/B _06100_/B _06100_/C vssd1 vssd1 vccd1 vccd1 _06404_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06054__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09740_ _09740_/A _09740_/B vssd1 vssd1 vccd1 vccd1 _09742_/A sky130_fd_sc_hd__nor2_1
X_06952_ _06952_/A _06952_/B vssd1 vssd1 vccd1 vccd1 _06953_/B sky130_fd_sc_hd__nand2_1
.ends

